module top(
  input LIOB33_SING_X0Y100_IOB_X0Y100_IPAD,
  input LIOB33_X0Y101_IOB_X0Y101_IPAD,
  input LIOB33_X0Y101_IOB_X0Y102_IPAD,
  input LIOB33_X0Y103_IOB_X0Y103_IPAD,
  input LIOB33_X0Y103_IOB_X0Y104_IPAD,
  input LIOB33_X0Y105_IOB_X0Y105_IPAD,
  input LIOB33_X0Y105_IOB_X0Y106_IPAD,
  input LIOB33_X0Y107_IOB_X0Y107_IPAD,
  input LIOB33_X0Y107_IOB_X0Y108_IPAD,
  input LIOB33_X0Y109_IOB_X0Y109_IPAD,
  input LIOB33_X0Y109_IOB_X0Y110_IPAD,
  input LIOB33_X0Y111_IOB_X0Y111_IPAD,
  input LIOB33_X0Y111_IOB_X0Y112_IPAD,
  input LIOB33_X0Y113_IOB_X0Y113_IPAD,
  input LIOB33_X0Y113_IOB_X0Y114_IPAD,
  input LIOB33_X0Y115_IOB_X0Y115_IPAD,
  input LIOB33_X0Y115_IOB_X0Y116_IPAD,
  input LIOB33_X0Y117_IOB_X0Y117_IPAD,
  input RIOB33_SING_X105Y100_IOB_X1Y100_IPAD,
  input RIOB33_X105Y101_IOB_X1Y101_IPAD,
  input RIOB33_X105Y101_IOB_X1Y102_IPAD,
  input RIOB33_X105Y103_IOB_X1Y103_IPAD,
  input RIOB33_X105Y103_IOB_X1Y104_IPAD,
  input RIOB33_X105Y105_IOB_X1Y105_IPAD,
  input RIOB33_X105Y105_IOB_X1Y106_IPAD,
  input RIOB33_X105Y107_IOB_X1Y107_IPAD,
  input RIOB33_X105Y107_IOB_X1Y108_IPAD,
  input RIOB33_X105Y109_IOB_X1Y109_IPAD,
  input RIOB33_X105Y109_IOB_X1Y110_IPAD,
  input RIOB33_X105Y111_IOB_X1Y111_IPAD,
  input RIOB33_X105Y111_IOB_X1Y112_IPAD,
  input RIOB33_X105Y113_IOB_X1Y113_IPAD,
  output LIOB33_SING_X0Y149_IOB_X0Y149_OPAD,
  output LIOB33_X0Y117_IOB_X0Y118_OPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD,
  output LIOB33_X0Y125_IOB_X0Y125_OPAD,
  output LIOB33_X0Y125_IOB_X0Y126_OPAD,
  output LIOB33_X0Y127_IOB_X0Y127_OPAD,
  output LIOB33_X0Y127_IOB_X0Y128_OPAD,
  output LIOB33_X0Y129_IOB_X0Y129_OPAD,
  output LIOB33_X0Y129_IOB_X0Y130_OPAD,
  output LIOB33_X0Y131_IOB_X0Y131_OPAD,
  output LIOB33_X0Y131_IOB_X0Y132_OPAD,
  output LIOB33_X0Y133_IOB_X0Y133_OPAD,
  output LIOB33_X0Y133_IOB_X0Y134_OPAD,
  output LIOB33_X0Y135_IOB_X0Y135_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output LIOB33_X0Y141_IOB_X0Y141_OPAD,
  output LIOB33_X0Y141_IOB_X0Y142_OPAD,
  output LIOB33_X0Y143_IOB_X0Y143_OPAD,
  output LIOB33_X0Y145_IOB_X0Y145_OPAD,
  output LIOB33_X0Y145_IOB_X0Y146_OPAD,
  output LIOB33_X0Y147_IOB_X0Y147_OPAD,
  output LIOB33_X0Y147_IOB_X0Y148_OPAD
  );
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_AMUX;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_AO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_AO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_BO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_BO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_CO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_CO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_DO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_DO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_AMUX;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_AO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_AO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_BO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_BO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_CO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_CO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_DO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_DO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_AMUX;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_AO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_BMUX;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_BO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_CO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_DO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_DO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_AMUX;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_AO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_BMUX;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_BO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_CO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_CO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_DMUX;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_DO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_DO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_AMUX;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_AO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_BO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_BO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_CO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_CO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_DO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_DO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_AMUX;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_AO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_BO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_BO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_CO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_CO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_DO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_DO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_AMUX;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_AO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_BMUX;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_BO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_BO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_CO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_DO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_DO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_AMUX;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_AO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_BO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_CO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_CO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_DO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_AMUX;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_BO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_CO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_DO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_DO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_AO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_AO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_BO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_BO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_CO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_CO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_DO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_DO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_AMUX;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_AO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_BMUX;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_BO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_BO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_CMUX;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_CO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_CO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_DO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_DO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_AO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_AO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_BO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_BO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_CO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_CO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_DO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_AMUX;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_AO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_BMUX;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_BO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_CO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_CO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_DO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_DO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_AMUX;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_AO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_BO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_CO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_CO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_DO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_AMUX;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_AO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_AO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_BO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_BO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_CO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_DO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_DO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_AO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_AO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_BO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_BO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_CO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_CO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_DO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_DO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_AO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_AO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_BO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_BO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_CO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_DO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_DO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_AMUX;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_AO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_AO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_BMUX;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_BO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_CO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_CO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_DO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_DO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_AMUX;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_AO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_AO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_BO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_BO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_CO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_DO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_DO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_AO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_AO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_BO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_BO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_CO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_CO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_DO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_DO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_AMUX;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_AO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_BMUX;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_BO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_CO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_DO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_DO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_AO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_AO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_BO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_CO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_DO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_BO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_CO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_DO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_AO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_BO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_CO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_DO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_DO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AMUX;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BMUX;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_DO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AMUX;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_BMUX;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_BO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_DO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AMUX;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_A_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_BO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_BO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_B_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_C_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_DO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X4Y110_D_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_AO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_A_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_BO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_B_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_CO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_C_XOR;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D1;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D2;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D3;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D4;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_DO5;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D_CY;
  wire [0:0] CLBLL_L_X4Y110_SLICE_X5Y110_D_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_BO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_DO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_BO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_CO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_DO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AMUX;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_BO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_DO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_BO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_DO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AMUX;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_DO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_AMUX;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_AO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_A_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_BMUX;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_BO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_B_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CMUX;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_C_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_DO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X4Y114_D_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_AMUX;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_AO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_AO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_A_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_BO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_BO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_B_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CMUX;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_CO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_C_XOR;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D1;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D2;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D3;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D4;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_DO5;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_DO6;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D_CY;
  wire [0:0] CLBLL_L_X4Y114_SLICE_X5Y114_D_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_A_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_BO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_B_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_C_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_DO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X4Y115_D_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AMUX;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_A_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_BO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_B_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_CO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_C_XOR;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D1;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D2;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D3;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D4;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_DO5;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_DO6;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D_CY;
  wire [0:0] CLBLL_L_X4Y115_SLICE_X5Y115_D_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_AMUX;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_AO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_AO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_BMUX;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_BO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_BO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_CMUX;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_CO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_CO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_DO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_DO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_AMUX;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_AO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_AO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_BO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_BO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_CO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_CO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_DO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_DO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_AO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_AO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_BO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_CO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_CO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_DMUX;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_DO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_DO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_AMUX;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_AO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_AO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_BMUX;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_BO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_BO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_CMUX;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_CO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_CO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_DO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_DO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_AO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_AO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_BO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_BO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_CMUX;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_CO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_CO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_DMUX;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_DO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_DO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_AO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_AO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_BO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_BO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_CO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_CO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_DO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_DO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_AO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_AO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_BO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_CO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_CO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_DO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_DO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_AO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_BO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_BO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_CO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_DO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_DO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_AO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_AO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_BO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_CO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_CO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_DO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_DO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_AMUX;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_AO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_BO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_CO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_DO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_AMUX;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_AO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_BO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_CO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_DO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_AMUX;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_AO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_BMUX;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_BO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_CO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_DO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_AMUX;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_AO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_BO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_CO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_DO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_AMUX;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_AO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_AO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_BO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_CO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_DO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_AMUX;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_AO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_AO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_BO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_BO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_CO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_DO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_DO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_AMUX;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_AO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_AO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_BO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_CO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_CO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_DMUX;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_DO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_AO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_AO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_BO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_BO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_CO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_CO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_DO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_AMUX;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_AO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_AO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_BMUX;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_BO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_CO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_DMUX;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_DO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_DO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_AMUX;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_AO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_A_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_BO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_BO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_B_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_CO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_CO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_C_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_DO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X12Y112_D_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_AMUX;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_AO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_AO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_A_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_BO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_B_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_CO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_CO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_C_XOR;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D1;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D2;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D3;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D4;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_DO5;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_DO6;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D_CY;
  wire [0:0] CLBLM_L_X10Y112_SLICE_X13Y112_D_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_AMUX;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_AO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_A_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_BO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_B_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_CO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_C_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_DO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X12Y113_D_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_AO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_AO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_A_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_BO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_B_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_CO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_C_XOR;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D1;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D2;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D3;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D4;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_DO5;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D_CY;
  wire [0:0] CLBLM_L_X10Y113_SLICE_X13Y113_D_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_AO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_AO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_A_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_BO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_BO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_B_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_CO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_CO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_C_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_DO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_DO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X16Y107_D_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_AO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_AO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_A_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_BO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_BO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_B_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_CO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_CO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_C_XOR;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D1;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D2;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D3;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D4;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_DO5;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_DO6;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D_CY;
  wire [0:0] CLBLM_L_X12Y107_SLICE_X17Y107_D_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_AO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_AO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_A_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_BO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_BO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_B_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_CO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_CO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_C_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_DO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_DO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X16Y108_D_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_AO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_AO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_A_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_BO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_BO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_B_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_CO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_CO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_C_XOR;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D1;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D2;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D3;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D4;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_DO5;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_DO6;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D_CY;
  wire [0:0] CLBLM_L_X12Y108_SLICE_X17Y108_D_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_AO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_AO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_A_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_BO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_BO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_B_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_CO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_CO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_C_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_DO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_DO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X16Y109_D_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_AO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_AO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_A_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_BO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_BO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_B_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_CO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_CO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_C_XOR;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D1;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D2;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D3;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D4;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_DO5;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_DO6;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D_CY;
  wire [0:0] CLBLM_L_X12Y109_SLICE_X17Y109_D_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_AO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_AO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_A_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_BO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_BO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_B_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_CO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_CO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_C_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_DO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_DO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X16Y110_D_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_AO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_AO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_A_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_BO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_BO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_B_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_CMUX;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_CO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_CO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_C_XOR;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D1;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D2;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D3;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D4;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_DO5;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_DO6;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D_CY;
  wire [0:0] CLBLM_L_X12Y110_SLICE_X17Y110_D_XOR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A1;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A2;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A3;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A4;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_AMUX;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_AO5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_AO6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A_CY;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A_XOR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B1;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B2;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B3;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B4;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_BO5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_BO6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B_CY;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B_XOR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C1;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C2;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C3;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C4;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_CO5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_CO6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C_CY;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C_XOR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D1;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D2;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D3;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D4;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_DO5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_DO6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D_CY;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D_XOR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A1;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A2;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A3;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A4;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_AMUX;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_AO5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_AO6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A_CY;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A_XOR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B1;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B2;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B3;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B4;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_BO5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_BO6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B_CY;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B_XOR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C1;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C2;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C3;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C4;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_CO5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_CO6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C_CY;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C_XOR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D1;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D2;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D3;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D4;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_DO5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_DO6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D_CY;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_AMUX;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_AO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_AO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_BO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_BO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_CO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_CO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_DO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_DO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_AO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_AO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_BO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_BO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_CO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_CO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_DO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_DO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_AO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_BO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_BO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_CO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_CO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_DO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_DO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_AO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_AO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_BO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_BO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_CO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_CO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_DO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_DO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_AMUX;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_AO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_AO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_BO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_BO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_CO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_CO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_DO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_DO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_AO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_AO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_BO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_BO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_CO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_CO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_DO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_DO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_AO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_AO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_BO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_BO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_CO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_CO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_DO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_DO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_AMUX;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_AO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_BO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_BO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_CO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_CO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_DO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_DO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_AMUX;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_AO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_AO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_BO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_CO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_CO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_DO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_DO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_AMUX;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_AO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_BO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_BO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_CO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_CO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_DO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_DO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_AMUX;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_AO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_BO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_CO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_CO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_DO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_DO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_AO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_BO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_BO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_CO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_CO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_DO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_DO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_AO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_AO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_BO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_CO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_DO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_DO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_AMUX;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_AO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_BO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_BO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_CO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_CO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_DO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_DO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_AMUX;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_AO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_BMUX;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_BO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_CO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_DO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_AMUX;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_AO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_BO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_CO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_DO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_AO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_BO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_CO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_DO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_AMUX;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_AO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_BMUX;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_BO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_CO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_DO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_DO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_AO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_BO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_CO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_DO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_AMUX;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_AO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_BO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_CO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_DO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_DO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AMUX;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_A_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_BMUX;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_BO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_B_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_CO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_C_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_DO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X10Y113_D_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_AO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_A_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_BO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_B_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_CO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_CO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_C_XOR;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D1;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D2;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D3;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D4;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_DO5;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_DO6;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D_CY;
  wire [0:0] CLBLM_L_X8Y113_SLICE_X11Y113_D_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_AMUX;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_AO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_AO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_A_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_BMUX;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_BO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_BO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_B_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_CO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_CO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_C_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_DO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_DO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X10Y114_D_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_AO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_AO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_A_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_BO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_BO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_B_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_CO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_CO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_C_XOR;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D1;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D2;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D3;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D4;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_DO5;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_DO6;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D_CY;
  wire [0:0] CLBLM_L_X8Y114_SLICE_X11Y114_D_XOR;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A1;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A2;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A3;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A4;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_AMUX;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_AO5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_AO6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A_CY;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A_XOR;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B1;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B2;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B3;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B4;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_BO5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_BO6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B_CY;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B_XOR;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C1;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C2;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C3;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C4;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_CO5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_CO6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C_CY;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C_XOR;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D1;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D2;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D3;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D4;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_DO5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_DO6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D_CY;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D_XOR;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A1;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A2;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A3;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A4;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_AO5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_AO6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A_CY;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A_XOR;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B1;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B2;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B3;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B4;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_BO5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_BO6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B_CY;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B_XOR;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C1;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C2;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C3;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C4;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_CO5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_CO6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C_CY;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C_XOR;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D1;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D2;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D3;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D4;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_DO5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_DO6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D_CY;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_AMUX;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_AO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_AO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_BO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_BO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_CO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_CO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_DO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_DO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_AMUX;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_AO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_AO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_BMUX;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_BO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_BO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_CO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_CO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_DO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_DO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_AMUX;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_AO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_BO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_CO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_DO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_DO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_AMUX;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_AO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_AO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_BO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_CO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_CO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_DO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_DO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_AMUX;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_AO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_AO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_BMUX;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_BO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_BO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_CO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_CO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_DO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_DO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_AMUX;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_AO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_AO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_BMUX;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_BO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_BO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_CMUX;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_CO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_CO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_DO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_DO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_AO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_AO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_BMUX;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_BO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_CO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_CO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_DO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_DO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_AMUX;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_AO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_AO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_BO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_BO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_CMUX;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_CO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_DO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_DO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_AO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_AO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_BO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_CO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_CO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_DO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_DO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_AO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_BMUX;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_BO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_BO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_CO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_CO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_DO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_DO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_AMUX;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_AO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_AO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_BO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_BO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_CO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_CO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_DO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_DO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_AMUX;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_AO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_AO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_BO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_BO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_CMUX;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_CO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_CO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_DO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_DO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_AMUX;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_AO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_AO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_A_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_BO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_BO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_B_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_CO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_CO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_C_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_DO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_DO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X14Y111_D_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_AO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_AO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_A_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_BO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_BO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_B_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_CO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_CO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_C_XOR;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D1;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D2;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D3;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D4;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_DO5;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_DO6;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D_CY;
  wire [0:0] CLBLM_R_X11Y111_SLICE_X15Y111_D_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_AO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_AO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_BO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_BO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_CO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_CO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_DO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_DO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_AO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_AO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_BO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_BO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_CO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_CO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_DO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_DO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_AMUX;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_AO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_AO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_BMUX;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_BO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_BO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_CMUX;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_CO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_CO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_DO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_DO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_AMUX;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_AO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_AO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_BMUX;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_BO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_CO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_CO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_DO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_DO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_AMUX;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_AO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_BO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_BO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_CO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_CO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_DO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_DO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_AMUX;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_AO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_AO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_BO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_CO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_DO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_DO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_AO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_AO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_BO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_BO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_CO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_DO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_DO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_AMUX;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_AO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_AO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_BO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_CO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_CO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_DO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_DO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_AO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_BO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_BO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_CO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_DO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_DO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_AMUX;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_AO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_AO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_BMUX;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_BO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_BO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_CO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_DO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_DO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_AMUX;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_AO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_AO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_BO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_BO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_CMUX;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_CO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_CO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_DO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_AO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_BO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_CO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_DO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AMUX;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_BO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_BO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_DO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_DO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AMUX;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_BMUX;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_BO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CMUX;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_DO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AMUX;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_BMUX;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_BO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_CO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_DO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AMUX;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_BO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_CO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_DO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_AMUX;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_BO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_CO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_DO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_DO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AMUX;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_BO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_CO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_DO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_BO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_CO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_DO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AMUX;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BMUX;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_DO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D_XOR;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_A;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_A1;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_A2;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_A3;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_A4;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_A5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_A6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_AMUX;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_AO5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_AO6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_A_CY;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_A_XOR;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_B;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_B1;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_B2;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_B3;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_B4;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_B5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_B6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_BO5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_BO6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_B_CY;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_B_XOR;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_C;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_C1;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_C2;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_C3;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_C4;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_C5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_C6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_CO5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_CO6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_C_CY;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_C_XOR;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_D;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_D1;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_D2;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_D3;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_D4;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_D5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_D6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_DO5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_DO6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_D_CY;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_D_XOR;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_A;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_A1;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_A2;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_A3;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_A4;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_A5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_A6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_AMUX;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_AO5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_AO6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_A_CY;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_A_XOR;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_B;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_B1;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_B2;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_B3;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_B4;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_B5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_B6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_BO5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_BO6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_B_CY;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_B_XOR;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_C;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_C1;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_C2;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_C3;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_C4;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_C5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_C6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_CO5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_CO6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_C_CY;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_C_XOR;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_D;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_D1;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_D2;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_D3;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_D4;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_D5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_D6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_DO5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_DO6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_D_CY;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_D_XOR;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_A;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_A1;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_A2;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_A3;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_A4;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_A5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_A6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_AMUX;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_AO5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_AO6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_A_CY;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_A_XOR;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_B;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_B1;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_B2;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_B3;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_B4;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_B5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_B6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_BO5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_BO6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_B_CY;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_B_XOR;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_C;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_C1;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_C2;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_C3;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_C4;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_C5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_C6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_CO5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_CO6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_C_CY;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_C_XOR;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_D;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_D1;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_D2;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_D3;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_D4;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_D5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_D6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_DO5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_DO6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_D_CY;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_D_XOR;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_A;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_A1;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_A2;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_A3;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_A4;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_A5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_A6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_AMUX;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_AO5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_AO6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_A_CY;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_A_XOR;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_B;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_B1;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_B2;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_B3;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_B4;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_B5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_B6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_BO5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_BO6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_B_CY;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_B_XOR;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_C;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_C1;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_C2;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_C3;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_C4;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_C5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_C6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_CO5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_CO6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_C_CY;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_C_XOR;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_D;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_D1;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_D2;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_D3;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_D4;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_D5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_D6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_DO5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_DO6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_D_CY;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_D_XOR;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A1;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A2;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A3;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A4;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_AMUX;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_AO5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_AO6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A_CY;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A_XOR;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B1;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B2;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B3;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B4;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_BO5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_BO6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B_CY;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B_XOR;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C1;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C2;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C3;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C4;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_CO5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_CO6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C_CY;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C_XOR;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D1;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D2;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D3;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D4;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_DO5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_DO6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D_CY;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D_XOR;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A1;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A2;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A3;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A4;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_AO5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_AO6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A_CY;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A_XOR;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B1;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B2;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B3;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B4;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_BO5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_BO6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B_CY;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B_XOR;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C1;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C2;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C3;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C4;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_CO5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_CO6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C_CY;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C_XOR;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D1;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D2;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D3;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D4;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_DO5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_DO6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D_CY;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_AO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_AO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_BO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_BO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_CO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_CO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_DO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_DO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_AO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_AO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_BO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_BO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_CO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_CO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_DO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_DO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_AMUX;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_AO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_BO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_BO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_CO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_CO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_DMUX;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_DO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_DO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_AO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_AO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_BO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_BO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_CO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_DO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_DO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_AMUX;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_AO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_BO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_CO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_DO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_AO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_AO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_BO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_CO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_CO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_DO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_DO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_AMUX;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_AO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_BO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_CO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_CO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_DO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_AO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_AO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_BO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_CO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_CO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_DO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_DO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_AO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_BO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_CO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_DO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_AO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_AO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_BO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_CO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_DO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_DO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_AO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_BO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_CO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_DO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AMUX;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_BO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_CO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_DO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_DO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_AO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_BO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_CO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_DO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_AO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_BO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_CO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_DO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_AMUX;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_AO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_BO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_CO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_DO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_AO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_BO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_CO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_DO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AMUX;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_BO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_CO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_DO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_BO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_BO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_CO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_CO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_DO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_AMUX;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_AO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_A_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_BO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_B_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_CO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_C_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_DO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X6Y113_D_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_AMUX;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_AO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_A_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_BMUX;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_BO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_B_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_CO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_CO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_C_XOR;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D1;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D2;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D3;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D4;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_DO5;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_DO6;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D_CY;
  wire [0:0] CLBLM_R_X5Y113_SLICE_X7Y113_D_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_AMUX;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_AO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_AO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_A_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_BO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_B_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_CO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_C_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_DO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_DO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X6Y114_D_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_AMUX;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_AO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_AO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_A_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_BO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_BO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_B_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_CO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_CO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_C_XOR;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D1;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D2;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D3;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D4;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_DO5;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_DO6;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D_CY;
  wire [0:0] CLBLM_R_X5Y114_SLICE_X7Y114_D_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_AMUX;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_AO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_A_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_BO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_B_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_CO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_C_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_DO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X6Y115_D_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_AMUX;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_AO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_A_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_BO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_BO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_B_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_CO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_C_XOR;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D1;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D2;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D3;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D4;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_DO5;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D_CY;
  wire [0:0] CLBLM_R_X5Y115_SLICE_X7Y115_D_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AMUX;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_BO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_DO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_BO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_BO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_DO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D_XOR;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A1;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A2;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A3;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A4;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_AMUX;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_AO5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_AO6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A_CY;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A_XOR;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B1;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B2;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B3;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B4;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_BMUX;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_BO5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_BO6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B_CY;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B_XOR;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C1;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C2;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C3;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C4;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_CMUX;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_CO5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_CO6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C_CY;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C_XOR;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D1;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D2;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D3;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D4;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_DO5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_DO6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D_CY;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D_XOR;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A1;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A2;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A3;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A4;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_AMUX;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_AO5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_AO6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A_CY;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A_XOR;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B1;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B2;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B3;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B4;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_BO5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_BO6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B_CY;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B_XOR;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C1;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C2;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C3;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C4;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_CMUX;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_CO5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_CO6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C_CY;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C_XOR;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D1;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D2;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D3;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D4;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_DO5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_DO6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D_CY;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_AO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_AO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_BO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_BO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_CO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_CO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_DO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_DO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_AO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_AO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_BO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_BO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_CO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_CO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_DO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_DO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_AMUX;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_AO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_AO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_BMUX;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_BO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_BO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_CO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_CO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_DO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_DO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_AO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_AO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_BO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_BO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_CO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_CO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_DO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_DO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_AMUX;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_AO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_AO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_BO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_BO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_CO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_CO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_DO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_DO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_AO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_AO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_BO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_BO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_CO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_CO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_DO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_DO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_AMUX;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_AO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_BO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_BO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_CO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_DO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_DO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_AO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_AO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_BO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_BO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_CO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_CO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_DO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_DO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_AMUX;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_AO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_BO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_BO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_CO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_CO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_DO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_DO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_AMUX;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_AO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_AO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_BMUX;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_BO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_CO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_CO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_DO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_DO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_AO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_BO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_CO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_CO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_DO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_DO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_AMUX;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_AO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_BO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_CO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_DO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_DO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_AMUX;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_AO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_BMUX;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_BO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_CO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_DO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_AO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_BO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_BO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_CO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_DO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_AMUX;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_AO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_AO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_BO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_CO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_DO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_AMUX;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_BO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_CO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_DO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_AMUX;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_AO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_BO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_CO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_DO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_AMUX;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_AO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_BO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_CO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_DO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_DO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_AO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_BO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_CO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_DO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_BO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_CO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_DO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AMUX;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_A_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_BO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_B_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_CO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_C_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_DO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X8Y113_D_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AMUX;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_A_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_BMUX;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_BO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_B_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_CO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_C_XOR;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D1;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D2;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D3;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D4;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_DO5;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D_CY;
  wire [0:0] CLBLM_R_X7Y113_SLICE_X9Y113_D_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_AO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_A_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_BO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_B_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_CO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_C_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_DO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X8Y114_D_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_AMUX;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_AO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_A_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_BO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_B_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_CMUX;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_CO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_CO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_C_XOR;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D1;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D2;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D3;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D4;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_DO5;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D_CY;
  wire [0:0] CLBLM_R_X7Y114_SLICE_X9Y114_D_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_AMUX;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_AO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_BMUX;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_BO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_BO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_CMUX;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_CO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_CO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_DO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_DO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_AO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_AO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_BO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_BO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_CO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_CO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_DO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D_XOR;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_I;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_O;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_O;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_D;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_O;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_O;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_O;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_TQ;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_I;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_D;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_O;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y105_SLICE_X0Y105_DO5),
.O6(CLBLL_L_X2Y105_SLICE_X0Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y105_SLICE_X0Y105_CO5),
.O6(CLBLL_L_X2Y105_SLICE_X0Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f13137f13137f7f)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLM_R_X3Y107_SLICE_X2Y107_BO6),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(CLBLL_L_X2Y105_SLICE_X0Y105_AO6),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLL_L_X2Y105_SLICE_X0Y105_BO5),
.O6(CLBLL_L_X2Y105_SLICE_X0Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3935c6c9f5f60a0)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLM_R_X3Y104_SLICE_X2Y104_BO6),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(CLBLM_R_X3Y104_SLICE_X3Y104_BO6),
.I5(CLBLL_L_X2Y106_SLICE_X0Y106_AO5),
.O5(CLBLL_L_X2Y105_SLICE_X0Y105_AO5),
.O6(CLBLL_L_X2Y105_SLICE_X0Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he080fef8fef8e080)
  ) CLBLL_L_X2Y105_SLICE_X1Y105_DLUT (
.I0(CLBLM_R_X3Y104_SLICE_X2Y104_BO6),
.I1(CLBLL_L_X2Y106_SLICE_X0Y106_AO5),
.I2(CLBLM_R_X3Y104_SLICE_X2Y104_AO6),
.I3(CLBLM_R_X3Y109_SLICE_X3Y109_AO5),
.I4(CLBLM_R_X3Y104_SLICE_X3Y104_BO6),
.I5(CLBLL_L_X4Y104_SLICE_X4Y104_AO6),
.O5(CLBLL_L_X2Y105_SLICE_X1Y105_DO5),
.O6(CLBLL_L_X2Y105_SLICE_X1Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a69a59669a5965a)
  ) CLBLL_L_X2Y105_SLICE_X1Y105_CLUT (
.I0(CLBLL_L_X4Y104_SLICE_X4Y104_AO6),
.I1(CLBLL_L_X2Y106_SLICE_X0Y106_AO5),
.I2(CLBLM_R_X3Y104_SLICE_X2Y104_AO6),
.I3(CLBLM_R_X3Y109_SLICE_X3Y109_AO5),
.I4(CLBLM_R_X3Y104_SLICE_X3Y104_BO6),
.I5(CLBLM_R_X3Y104_SLICE_X2Y104_BO6),
.O5(CLBLL_L_X2Y105_SLICE_X1Y105_CO5),
.O6(CLBLL_L_X2Y105_SLICE_X1Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he9c94fefb9391f1f)
  ) CLBLL_L_X2Y105_SLICE_X1Y105_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLL_L_X2Y105_SLICE_X1Y105_BO5),
.O6(CLBLL_L_X2Y105_SLICE_X1Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3fc03fc0eaea8080)
  ) CLBLL_L_X2Y105_SLICE_X1Y105_ALUT (
.I0(CLBLL_L_X2Y106_SLICE_X0Y106_AO5),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(CLBLL_L_X2Y105_SLICE_X1Y105_BO6),
.I4(CLBLM_R_X3Y104_SLICE_X2Y104_BO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y105_SLICE_X1Y105_AO5),
.O6(CLBLL_L_X2Y105_SLICE_X1Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_DO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8778778878878877)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(CLBLL_L_X2Y105_SLICE_X0Y105_AO6),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(CLBLM_R_X3Y107_SLICE_X2Y107_BO6),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_CO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc95593ff36aa6c00)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_BLUT (
.I0(CLBLL_L_X2Y107_SLICE_X0Y107_AO5),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(CLBLL_L_X2Y105_SLICE_X1Y105_AO6),
.I5(CLBLL_L_X2Y105_SLICE_X0Y105_AO6),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_BO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7bc00cc040c0ccc0)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_ALUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_AO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd00d4004fddff44f)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_DLUT (
.I0(CLBLL_L_X2Y106_SLICE_X1Y106_AO6),
.I1(CLBLL_L_X2Y106_SLICE_X0Y106_CO6),
.I2(CLBLM_R_X3Y105_SLICE_X2Y105_AO6),
.I3(CLBLL_L_X2Y106_SLICE_X1Y106_AO5),
.I4(CLBLM_R_X3Y108_SLICE_X2Y108_DO6),
.I5(CLBLL_L_X2Y106_SLICE_X1Y106_BO6),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_DO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4800de5ac000fcf0)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(CLBLL_L_X2Y106_SLICE_X0Y106_BO6),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(CLBLM_R_X3Y108_SLICE_X2Y108_DO6),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_CO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000ff000000)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(1'b1),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_BO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ff000000)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(1'b1),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_AO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfec4c804c804c80)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_DLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLL_L_X2Y108_SLICE_X0Y108_CO6),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(CLBLL_L_X2Y107_SLICE_X0Y107_CO6),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_DO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h63ffc6aa9c003955)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_CLUT (
.I0(CLBLL_L_X2Y107_SLICE_X0Y107_AO6),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(CLBLL_L_X2Y108_SLICE_X0Y108_BO5),
.I5(CLBLM_R_X3Y107_SLICE_X2Y107_AO6),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_CO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3bbcf770c443088f)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(CLBLL_L_X2Y107_SLICE_X1Y107_AO6),
.I3(CLBLL_L_X2Y108_SLICE_X0Y108_AO5),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLM_R_X3Y107_SLICE_X3Y107_CO6),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_BO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc3300ff4d4d0505)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_ALUT (
.I0(CLBLL_L_X2Y106_SLICE_X0Y106_AO6),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(CLBLL_L_X2Y107_SLICE_X1Y107_AO5),
.I3(CLBLM_R_X3Y107_SLICE_X3Y107_CO6),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_AO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h956aa95656565656)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_DLUT (
.I0(CLBLM_R_X3Y105_SLICE_X2Y105_AO6),
.I1(CLBLL_L_X2Y106_SLICE_X0Y106_CO6),
.I2(CLBLM_R_X3Y108_SLICE_X2Y108_DO6),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_DO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h96693cc36969c3c3)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLL_L_X2Y106_SLICE_X0Y106_BO6),
.I2(CLBLM_R_X3Y108_SLICE_X2Y108_DO6),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_CO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha59a556a9a5a6aaa)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_BLUT (
.I0(CLBLL_L_X2Y107_SLICE_X1Y107_DO6),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLL_L_X2Y107_SLICE_X0Y107_DO6),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(CLBLL_L_X2Y107_SLICE_X1Y107_CO6),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_BO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h59aacc00c455ffff)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_ALUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_AO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf773fddc3110c440)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_DLUT (
.I0(CLBLL_L_X2Y108_SLICE_X0Y108_AO6),
.I1(CLBLL_L_X2Y109_SLICE_X0Y109_CO6),
.I2(CLBLL_L_X2Y110_SLICE_X0Y110_AO6),
.I3(CLBLL_L_X2Y111_SLICE_X0Y111_AO6),
.I4(CLBLM_R_X3Y108_SLICE_X2Y108_AO6),
.I5(CLBLL_L_X2Y108_SLICE_X1Y108_AO6),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_DO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8fff0888f8888000)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(CLBLL_L_X2Y108_SLICE_X0Y108_DO6),
.I5(CLBLL_L_X2Y107_SLICE_X0Y107_BO6),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_CO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aaff00d4d4fcfc)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_BLUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(CLBLL_L_X2Y108_SLICE_X0Y108_AO5),
.I2(CLBLL_L_X2Y107_SLICE_X1Y107_AO6),
.I3(CLBLL_L_X2Y109_SLICE_X0Y109_CO6),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_BO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6e44a288b333ff77)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_ALUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_AO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3b2b230fce8e8c0)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_DLUT (
.I0(CLBLM_R_X3Y108_SLICE_X2Y108_BO6),
.I1(CLBLM_R_X3Y107_SLICE_X2Y107_CO6),
.I2(CLBLM_R_X3Y109_SLICE_X2Y109_AO6),
.I3(CLBLL_L_X2Y108_SLICE_X1Y108_AO5),
.I4(CLBLL_L_X2Y108_SLICE_X0Y108_CO6),
.I5(CLBLL_L_X2Y106_SLICE_X1Y106_AO6),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_DO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hebc38200af0f0a00)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(CLBLL_L_X2Y107_SLICE_X1Y107_DO6),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(CLBLL_L_X2Y108_SLICE_X1Y108_DO6),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_CO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c939393936c6c6c)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_BLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(CLBLM_R_X3Y106_SLICE_X2Y106_AO6),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLL_L_X2Y108_SLICE_X1Y108_CO6),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_BO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00a0a0a0a0)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_ALUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(1'b1),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_AO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c39933963c66cc)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(CLBLL_L_X2Y108_SLICE_X0Y108_CO6),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(CLBLL_L_X2Y107_SLICE_X0Y107_CO6),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_DO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hee917f3ba2dd3377)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_CO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h43c48f08bc3b70f7)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_BLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(CLBLL_L_X2Y108_SLICE_X0Y108_AO6),
.I3(CLBLL_L_X2Y110_SLICE_X0Y110_AO6),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(CLBLL_L_X2Y109_SLICE_X0Y109_CO6),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_BO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h93939393aa5500ff)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_ALUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(CLBLL_L_X2Y107_SLICE_X1Y107_BO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(CLBLL_L_X2Y109_SLICE_X0Y109_BO6),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_AO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_DO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_CO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_BO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fa0609f609fa05f)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(CLBLM_R_X3Y107_SLICE_X2Y107_CO6),
.I4(CLBLM_R_X3Y108_SLICE_X2Y108_BO6),
.I5(CLBLL_L_X2Y108_SLICE_X0Y108_CO6),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_AO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h566af000a9950fff)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(CLBLL_L_X2Y108_SLICE_X0Y108_BO6),
.I3(CLBLL_L_X2Y110_SLICE_X0Y110_CO6),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLL_L_X2Y107_SLICE_X0Y107_BO6),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_DO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha000faaac333c333)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_CLUT (
.I0(CLBLL_L_X2Y110_SLICE_X0Y110_AO6),
.I1(CLBLL_L_X2Y110_SLICE_X1Y110_AO6),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(CLBLL_L_X2Y108_SLICE_X0Y108_AO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_CO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h99995555c03fc03f)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_BLUT (
.I0(CLBLL_L_X2Y110_SLICE_X0Y110_DO6),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLL_L_X2Y109_SLICE_X1Y109_AO6),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_BO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h70f03000b30f43ff)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_ALUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_AO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_DO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_CO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_BO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h083078cc4cfc3c00)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_ALUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_AO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_DO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_CO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888c03f3fc0)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_BLUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(CLBLM_R_X3Y106_SLICE_X3Y106_AO6),
.I4(CLBLM_R_X3Y108_SLICE_X3Y108_AO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_BO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c077777777)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_ALUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_AO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_DO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_CO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h936c6c936c6c9393)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_BLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(CLBLM_R_X3Y108_SLICE_X3Y108_CO6),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(CLBLM_R_X3Y108_SLICE_X3Y108_BO6),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_BO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3c33333a555a555)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_ALUT (
.I0(CLBLM_R_X3Y111_SLICE_X2Y111_CO6),
.I1(CLBLM_R_X3Y109_SLICE_X2Y109_BO6),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_AO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h96693cc35aa5f00f)
  ) CLBLL_L_X4Y104_SLICE_X4Y104_DLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(CLBLM_R_X5Y101_SLICE_X6Y101_BO6),
.I3(CLBLL_L_X4Y104_SLICE_X4Y104_CO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLL_L_X4Y104_SLICE_X4Y104_DO5),
.O6(CLBLL_L_X4Y104_SLICE_X4Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbe3c28be3c2800)
  ) CLBLL_L_X4Y104_SLICE_X4Y104_CLUT (
.I0(CLBLL_L_X4Y104_SLICE_X4Y104_AO6),
.I1(CLBLM_R_X3Y103_SLICE_X3Y103_AO6),
.I2(CLBLM_R_X5Y101_SLICE_X6Y101_AO5),
.I3(CLBLM_R_X3Y104_SLICE_X2Y104_BO5),
.I4(CLBLM_R_X3Y104_SLICE_X2Y104_AO5),
.I5(CLBLM_R_X5Y102_SLICE_X6Y102_AO6),
.O5(CLBLL_L_X4Y104_SLICE_X4Y104_CO5),
.O6(CLBLL_L_X4Y104_SLICE_X4Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9696966996696969)
  ) CLBLL_L_X4Y104_SLICE_X4Y104_BLUT (
.I0(CLBLM_R_X5Y101_SLICE_X6Y101_AO5),
.I1(CLBLM_R_X3Y104_SLICE_X2Y104_AO5),
.I2(CLBLM_R_X3Y103_SLICE_X3Y103_AO6),
.I3(CLBLM_R_X5Y102_SLICE_X6Y102_AO6),
.I4(CLBLL_L_X4Y104_SLICE_X4Y104_AO6),
.I5(CLBLM_R_X3Y104_SLICE_X2Y104_BO5),
.O5(CLBLL_L_X4Y104_SLICE_X4Y104_BO5),
.O6(CLBLL_L_X4Y104_SLICE_X4Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000cccc0000)
  ) CLBLL_L_X4Y104_SLICE_X4Y104_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(1'b1),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y104_SLICE_X4Y104_AO5),
.O6(CLBLL_L_X4Y104_SLICE_X4Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff7b5a127b5a1200)
  ) CLBLL_L_X4Y104_SLICE_X5Y104_DLUT (
.I0(CLBLM_R_X5Y103_SLICE_X6Y103_BO6),
.I1(CLBLM_R_X5Y103_SLICE_X6Y103_CO6),
.I2(CLBLM_R_X5Y105_SLICE_X6Y105_AO6),
.I3(CLBLL_L_X4Y105_SLICE_X5Y105_AO5),
.I4(CLBLL_L_X4Y105_SLICE_X5Y105_BO5),
.I5(CLBLL_L_X4Y104_SLICE_X5Y104_BO6),
.O5(CLBLL_L_X4Y104_SLICE_X5Y104_DO5),
.O6(CLBLL_L_X4Y104_SLICE_X5Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a6696669655a555)
  ) CLBLL_L_X4Y104_SLICE_X5Y104_CLUT (
.I0(CLBLM_R_X5Y103_SLICE_X6Y103_BO6),
.I1(CLBLM_R_X5Y103_SLICE_X6Y103_CO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLL_L_X4Y104_SLICE_X5Y104_BO6),
.O5(CLBLL_L_X4Y104_SLICE_X5Y104_CO5),
.O6(CLBLL_L_X4Y104_SLICE_X5Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8f08ff88f8808800)
  ) CLBLL_L_X4Y104_SLICE_X5Y104_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(CLBLL_L_X4Y104_SLICE_X4Y104_CO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_R_X5Y101_SLICE_X6Y101_BO6),
.O5(CLBLL_L_X4Y104_SLICE_X5Y104_BO5),
.O6(CLBLL_L_X4Y104_SLICE_X5Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5695a96695a96a5)
  ) CLBLL_L_X4Y104_SLICE_X5Y104_ALUT (
.I0(CLBLL_L_X4Y105_SLICE_X5Y105_BO5),
.I1(CLBLM_R_X5Y103_SLICE_X6Y103_CO6),
.I2(CLBLM_R_X5Y105_SLICE_X6Y105_AO6),
.I3(CLBLL_L_X4Y104_SLICE_X5Y104_BO6),
.I4(CLBLM_R_X5Y103_SLICE_X6Y103_BO6),
.I5(CLBLL_L_X4Y105_SLICE_X5Y105_AO5),
.O5(CLBLL_L_X4Y104_SLICE_X5Y104_AO5),
.O6(CLBLL_L_X4Y104_SLICE_X5Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf990f55090905050)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_DLUT (
.I0(CLBLM_R_X3Y104_SLICE_X3Y104_DO6),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(CLBLM_R_X3Y105_SLICE_X3Y105_CO6),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLL_L_X4Y105_SLICE_X4Y105_DO5),
.O6(CLBLL_L_X4Y105_SLICE_X4Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf9f990f990f99090)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_CLUT (
.I0(CLBLM_R_X5Y105_SLICE_X6Y105_BO6),
.I1(CLBLL_L_X4Y105_SLICE_X5Y105_AO5),
.I2(CLBLL_L_X4Y105_SLICE_X5Y105_BO6),
.I3(CLBLL_L_X4Y104_SLICE_X4Y104_DO6),
.I4(CLBLM_R_X3Y105_SLICE_X3Y105_CO6),
.I5(CLBLL_L_X4Y105_SLICE_X5Y105_AO6),
.O5(CLBLL_L_X4Y105_SLICE_X4Y105_CO5),
.O6(CLBLL_L_X4Y105_SLICE_X4Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93936c36c9c936)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_BLUT (
.I0(CLBLM_R_X3Y105_SLICE_X3Y105_CO6),
.I1(CLBLL_L_X4Y105_SLICE_X5Y105_BO6),
.I2(CLBLL_L_X4Y105_SLICE_X5Y105_AO6),
.I3(CLBLL_L_X4Y105_SLICE_X5Y105_AO5),
.I4(CLBLM_R_X5Y105_SLICE_X6Y105_BO6),
.I5(CLBLL_L_X4Y104_SLICE_X4Y104_DO6),
.O5(CLBLL_L_X4Y105_SLICE_X4Y105_BO5),
.O6(CLBLL_L_X4Y105_SLICE_X4Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h963cccccc3966666)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_ALUT (
.I0(CLBLM_R_X3Y105_SLICE_X3Y105_CO6),
.I1(CLBLM_R_X5Y105_SLICE_X6Y105_BO6),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(CLBLL_L_X4Y104_SLICE_X4Y104_DO6),
.O5(CLBLL_L_X4Y105_SLICE_X4Y105_AO5),
.O6(CLBLL_L_X4Y105_SLICE_X4Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h96665aaa6999a555)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_DLUT (
.I0(CLBLM_R_X5Y101_SLICE_X6Y101_CO6),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(CLBLL_L_X4Y104_SLICE_X5Y104_BO6),
.O5(CLBLL_L_X4Y105_SLICE_X5Y105_DO5),
.O6(CLBLL_L_X4Y105_SLICE_X5Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he7184db2659acf30)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLL_L_X4Y105_SLICE_X5Y105_DO6),
.I2(CLBLL_L_X4Y105_SLICE_X4Y105_DO6),
.I3(CLBLL_L_X4Y104_SLICE_X5Y104_CO6),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLL_L_X4Y105_SLICE_X5Y105_CO5),
.O6(CLBLL_L_X4Y105_SLICE_X5Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000ff000000)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(1'b1),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y105_SLICE_X5Y105_BO5),
.O6(CLBLL_L_X4Y105_SLICE_X5Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f000f000)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y105_SLICE_X5Y105_AO5),
.O6(CLBLL_L_X4Y105_SLICE_X5Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_DO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969966996699696)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_CLUT (
.I0(CLBLL_L_X4Y104_SLICE_X5Y104_AO6),
.I1(CLBLL_L_X4Y105_SLICE_X4Y105_CO6),
.I2(CLBLL_L_X4Y106_SLICE_X4Y106_AO6),
.I3(CLBLL_L_X4Y106_SLICE_X4Y106_AO5),
.I4(CLBLM_R_X3Y106_SLICE_X2Y106_DO6),
.I5(CLBLL_L_X4Y105_SLICE_X4Y105_BO6),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_CO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a56fcfc95a90303)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(CLBLM_R_X3Y106_SLICE_X3Y106_CO6),
.I2(CLBLM_R_X3Y107_SLICE_X3Y107_DO6),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(CLBLL_L_X4Y106_SLICE_X4Y106_CO6),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_BO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00aa00aa00)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(1'b1),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_AO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_DO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_CO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_BO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996669999666996)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_ALUT (
.I0(CLBLL_L_X4Y104_SLICE_X5Y104_DO6),
.I1(CLBLM_R_X5Y106_SLICE_X6Y106_AO6),
.I2(CLBLL_L_X4Y106_SLICE_X4Y106_AO6),
.I3(CLBLM_R_X5Y104_SLICE_X6Y104_AO6),
.I4(CLBLL_L_X4Y104_SLICE_X5Y104_AO6),
.I5(CLBLL_L_X4Y105_SLICE_X4Y105_CO6),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_AO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc639639c39c69c63)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_DLUT (
.I0(CLBLL_L_X4Y107_SLICE_X4Y107_AO6),
.I1(CLBLL_L_X4Y106_SLICE_X4Y106_CO6),
.I2(CLBLM_R_X3Y106_SLICE_X3Y106_CO6),
.I3(CLBLL_L_X4Y107_SLICE_X4Y107_AO5),
.I4(CLBLM_R_X3Y107_SLICE_X3Y107_DO6),
.I5(CLBLL_L_X4Y107_SLICE_X4Y107_BO6),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_DO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h60f6f6f6a0fafafa)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_CLUT (
.I0(CLBLL_L_X4Y105_SLICE_X4Y105_AO6),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(CLBLM_R_X3Y106_SLICE_X2Y106_DO6),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_CO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000cc00cc00)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_BO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f000f000)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_AO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_DO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a5c30f965a3cf0)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(CLBLM_R_X5Y105_SLICE_X6Y105_CO6),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLL_L_X4Y107_SLICE_X5Y107_BO6),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_CO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hebc3bb3382002200)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(CLBLL_L_X4Y104_SLICE_X5Y104_CO6),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLL_L_X4Y105_SLICE_X4Y105_CO6),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_BO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93a05f936c5fa0)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(CLBLL_L_X4Y104_SLICE_X5Y104_CO6),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLL_L_X4Y105_SLICE_X4Y105_CO6),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_AO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h405480a8d5fdeafe)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_DLUT (
.I0(CLBLL_L_X4Y106_SLICE_X5Y106_AO6),
.I1(CLBLL_L_X4Y107_SLICE_X5Y107_AO6),
.I2(CLBLL_L_X4Y107_SLICE_X4Y107_CO6),
.I3(CLBLL_L_X4Y107_SLICE_X4Y107_AO5),
.I4(CLBLM_R_X5Y107_SLICE_X6Y107_AO6),
.I5(CLBLL_L_X4Y107_SLICE_X4Y107_BO5),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_DO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h95a96a566a5695a9)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_CLUT (
.I0(CLBLL_L_X4Y106_SLICE_X5Y106_AO6),
.I1(CLBLL_L_X4Y107_SLICE_X5Y107_AO6),
.I2(CLBLL_L_X4Y107_SLICE_X4Y107_CO6),
.I3(CLBLL_L_X4Y107_SLICE_X4Y107_AO5),
.I4(CLBLM_R_X5Y107_SLICE_X6Y107_AO6),
.I5(CLBLL_L_X4Y107_SLICE_X4Y107_BO5),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_CO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h90c06f3f3595ca6a)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_BLUT (
.I0(CLBLL_L_X4Y107_SLICE_X5Y107_AO6),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(CLBLL_L_X4Y106_SLICE_X5Y106_AO6),
.I5(CLBLL_L_X4Y107_SLICE_X4Y107_CO6),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_BO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h96663ccc6999c333)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(CLBLL_L_X4Y105_SLICE_X5Y105_CO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(CLBLL_L_X4Y107_SLICE_X4Y107_CO6),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_AO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_DO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfff3b3f3fbf222a)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_CLUT (
.I0(CLBLL_L_X4Y107_SLICE_X5Y107_CO6),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(CLBLM_R_X5Y107_SLICE_X6Y107_DO6),
.I5(CLBLL_L_X4Y108_SLICE_X5Y108_BO6),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_CO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffdf5f135f4c00)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(CLBLL_L_X4Y105_SLICE_X5Y105_CO6),
.I5(CLBLL_L_X4Y107_SLICE_X4Y107_CO6),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_BO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8a1975e620b3df4c)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_ALUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(CLBLL_L_X4Y107_SLICE_X5Y107_CO6),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(CLBLL_L_X4Y108_SLICE_X5Y108_BO6),
.I4(CLBLM_R_X5Y107_SLICE_X6Y107_BO6),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_AO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a5695a995a96a56)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_DLUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.I1(CLBLL_L_X4Y108_SLICE_X5Y108_CO6),
.I2(CLBLL_L_X4Y109_SLICE_X5Y109_BO5),
.I3(CLBLL_L_X4Y109_SLICE_X4Y109_AO5),
.I4(CLBLM_R_X5Y109_SLICE_X6Y109_DO6),
.I5(CLBLM_R_X3Y109_SLICE_X3Y109_BO5),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_DO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h936cc936c936936c)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_CLUT (
.I0(CLBLL_L_X4Y109_SLICE_X4Y109_AO6),
.I1(CLBLL_L_X4Y109_SLICE_X5Y109_CO6),
.I2(CLBLM_R_X3Y108_SLICE_X3Y108_DO6),
.I3(CLBLL_L_X4Y109_SLICE_X4Y109_AO5),
.I4(CLBLL_L_X4Y108_SLICE_X5Y108_AO6),
.I5(CLBLL_L_X4Y109_SLICE_X5Y109_AO6),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_CO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3c3c33f030303)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y109_SLICE_X5Y109_BO5),
.I2(CLBLL_L_X4Y108_SLICE_X5Y108_CO6),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_BO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0cc00cc00)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_AO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb42d4bd24bd2b42d)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_DLUT (
.I0(CLBLL_L_X4Y109_SLICE_X5Y109_BO5),
.I1(CLBLL_L_X4Y109_SLICE_X4Y109_AO5),
.I2(CLBLM_R_X5Y108_SLICE_X6Y108_BO6),
.I3(CLBLL_L_X4Y108_SLICE_X5Y108_CO6),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.I5(CLBLL_L_X4Y109_SLICE_X5Y109_BO6),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_DO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2bd4d42bd42b2bd4)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_CLUT (
.I0(CLBLL_L_X4Y109_SLICE_X5Y109_AO6),
.I1(CLBLM_R_X5Y107_SLICE_X6Y107_DO6),
.I2(CLBLL_L_X4Y108_SLICE_X4Y108_DO6),
.I3(CLBLM_R_X7Y108_SLICE_X8Y108_AO6),
.I4(CLBLM_L_X8Y111_SLICE_X11Y111_AO6),
.I5(CLBLM_R_X5Y107_SLICE_X6Y107_CO6),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_CO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf0c0c0cc33c3c3c)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y107_SLICE_X6Y107_CO6),
.I2(CLBLM_R_X7Y108_SLICE_X8Y108_AO6),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_BO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00cc0033ff)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(1'b1),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(CLBLL_L_X4Y108_SLICE_X5Y108_AO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_AO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5fad4e8d4e850a0)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_DLUT (
.I0(CLBLL_L_X4Y110_SLICE_X4Y110_AO6),
.I1(CLBLM_R_X3Y109_SLICE_X3Y109_BO5),
.I2(CLBLM_R_X5Y112_SLICE_X6Y112_AO6),
.I3(CLBLM_R_X5Y109_SLICE_X6Y109_BO6),
.I4(CLBLL_L_X4Y109_SLICE_X4Y109_BO5),
.I5(CLBLM_R_X5Y109_SLICE_X6Y109_CO6),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_DO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4004d00df44ffddf)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_CLUT (
.I0(CLBLL_L_X4Y110_SLICE_X4Y110_AO6),
.I1(CLBLM_R_X5Y110_SLICE_X7Y110_AO6),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_AO5),
.I3(CLBLM_R_X7Y109_SLICE_X8Y109_CO6),
.I4(CLBLM_R_X5Y109_SLICE_X6Y109_AO6),
.I5(CLBLM_R_X3Y110_SLICE_X3Y110_AO6),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_CO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5965a69965a69a5)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_BLUT (
.I0(CLBLM_R_X5Y112_SLICE_X6Y112_AO6),
.I1(CLBLL_L_X4Y109_SLICE_X4Y109_BO5),
.I2(CLBLM_R_X5Y109_SLICE_X6Y109_BO6),
.I3(CLBLM_R_X5Y109_SLICE_X6Y109_CO6),
.I4(CLBLL_L_X4Y110_SLICE_X4Y110_AO6),
.I5(CLBLM_R_X3Y109_SLICE_X3Y109_BO5),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_BO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0c0ff00c0)
  ) CLBLL_L_X4Y110_SLICE_X4Y110_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLM_R_X5Y110_SLICE_X7Y110_AO6),
.I4(CLBLM_R_X5Y109_SLICE_X6Y109_AO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X4Y110_AO5),
.O6(CLBLL_L_X4Y110_SLICE_X4Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_DO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_CO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_BO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h399993336369c9c3)
  ) CLBLL_L_X4Y110_SLICE_X5Y110_ALUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(CLBLM_R_X7Y109_SLICE_X8Y109_CO6),
.I2(CLBLM_R_X5Y109_SLICE_X6Y109_AO6),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLM_R_X5Y110_SLICE_X7Y110_AO6),
.O5(CLBLL_L_X4Y110_SLICE_X5Y110_AO5),
.O6(CLBLL_L_X4Y110_SLICE_X5Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_DO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_CO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h96695aa56969a5a5)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_BLUT (
.I0(CLBLL_L_X4Y110_SLICE_X4Y110_DO6),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(CLBLL_L_X4Y110_SLICE_X5Y110_AO6),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_BO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h157f40d57f7fd5d5)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_ALUT (
.I0(CLBLL_L_X4Y110_SLICE_X4Y110_DO6),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(CLBLL_L_X4Y110_SLICE_X5Y110_AO6),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_AO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_DO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_CO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_BO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_AO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999966696669666)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_DLUT (
.I0(CLBLL_L_X4Y110_SLICE_X4Y110_CO6),
.I1(CLBLL_L_X4Y112_SLICE_X5Y112_AO6),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_DO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd777411141114111)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_CLUT (
.I0(CLBLL_L_X4Y110_SLICE_X4Y110_CO6),
.I1(CLBLL_L_X4Y112_SLICE_X5Y112_AO6),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_CO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2d87787887872d87)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(CLBLL_L_X4Y112_SLICE_X5Y112_AO6),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_AO6),
.I5(CLBLL_L_X4Y110_SLICE_X4Y110_AO5),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_BO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3fc0c03fc0c0c0c0)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(CLBLM_R_X5Y111_SLICE_X6Y111_CO6),
.I4(CLBLM_R_X5Y110_SLICE_X7Y110_BO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_AO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_DO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_CO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_BO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h693cccccc3699999)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_ALUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_CO6),
.I1(CLBLM_R_X7Y111_SLICE_X8Y111_CO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(CLBLM_R_X5Y110_SLICE_X7Y110_BO6),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_AO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7e8156a9d42bfc03)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_DLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLM_R_X5Y110_SLICE_X7Y110_BO6),
.I2(CLBLM_R_X5Y111_SLICE_X6Y111_CO6),
.I3(CLBLM_R_X7Y109_SLICE_X9Y109_BO6),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(LIOB33_X0Y113_IOB_X0Y113_I),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_DO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9c6339c6639cc639)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_CLUT (
.I0(CLBLL_L_X4Y110_SLICE_X4Y110_CO6),
.I1(CLBLM_R_X7Y113_SLICE_X8Y113_DO6),
.I2(CLBLM_R_X3Y112_SLICE_X3Y112_AO5),
.I3(CLBLL_L_X4Y113_SLICE_X4Y113_AO5),
.I4(CLBLL_L_X4Y113_SLICE_X4Y113_DO6),
.I5(CLBLL_L_X4Y113_SLICE_X4Y113_BO6),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_CO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2b000000ff2b0303)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_BLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(CLBLM_R_X5Y111_SLICE_X6Y111_CO6),
.I2(CLBLM_R_X5Y110_SLICE_X7Y110_BO6),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLM_R_X7Y109_SLICE_X9Y109_BO6),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_BO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000f000f000)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_AO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_DO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_CO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_BO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_AO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heb82af0ac3000f00)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_DLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_R_X5Y111_SLICE_X6Y111_DO6),
.I3(CLBLL_L_X4Y113_SLICE_X4Y113_BO6),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_DO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887877887788778)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(CLBLM_R_X5Y111_SLICE_X6Y111_DO6),
.I3(CLBLL_L_X4Y113_SLICE_X4Y113_BO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(LIOB33_X0Y113_IOB_X0Y113_I),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_CO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h96c33c968ecf0c8e)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_BLUT (
.I0(CLBLM_R_X3Y111_SLICE_X3Y111_DO6),
.I1(CLBLL_L_X4Y114_SLICE_X5Y114_BO6),
.I2(CLBLL_L_X4Y114_SLICE_X4Y114_DO6),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_CO6),
.I4(CLBLL_L_X4Y114_SLICE_X4Y114_CO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_BO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h9999666633330000)
  ) CLBLL_L_X4Y114_SLICE_X4Y114_ALUT (
.I0(CLBLM_R_X3Y111_SLICE_X3Y111_DO6),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_CO6),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X4Y114_SLICE_X4Y114_CO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X4Y114_AO5),
.O6(CLBLL_L_X4Y114_SLICE_X4Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaff8aef0aaf08ae)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_DLUT (
.I0(CLBLM_R_X5Y114_SLICE_X6Y114_AO6),
.I1(CLBLL_L_X4Y114_SLICE_X4Y114_AO5),
.I2(CLBLL_L_X4Y114_SLICE_X4Y114_DO6),
.I3(CLBLL_L_X4Y114_SLICE_X5Y114_CO6),
.I4(CLBLM_R_X3Y112_SLICE_X3Y112_DO6),
.I5(CLBLL_L_X4Y114_SLICE_X5Y114_BO6),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_DO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he8c088008e0ceecc)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_R_X5Y112_SLICE_X6Y112_BO6),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(CLBLM_R_X7Y113_SLICE_X8Y113_AO6),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_CO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887887787787788)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(LIOB33_X0Y113_IOB_X0Y113_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(CLBLM_R_X7Y113_SLICE_X8Y113_AO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_R_X5Y112_SLICE_X6Y112_BO6),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_BO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h965aa596cc3333cc)
  ) CLBLL_L_X4Y114_SLICE_X5Y114_ALUT (
.I0(CLBLM_R_X5Y114_SLICE_X6Y114_AO5),
.I1(CLBLM_R_X5Y114_SLICE_X6Y114_AO6),
.I2(CLBLM_R_X7Y114_SLICE_X8Y114_AO6),
.I3(CLBLL_L_X4Y114_SLICE_X4Y114_BO5),
.I4(CLBLL_L_X4Y114_SLICE_X5Y114_CO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y114_SLICE_X5Y114_AO5),
.O6(CLBLL_L_X4Y114_SLICE_X5Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_DO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_CO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_BO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y115_SLICE_X4Y115_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X4Y115_AO5),
.O6(CLBLL_L_X4Y115_SLICE_X4Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_DO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_CO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000bb22bb22ffff)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_BLUT (
.I0(CLBLL_L_X4Y114_SLICE_X5Y114_DO6),
.I1(CLBLM_R_X5Y114_SLICE_X6Y114_AO5),
.I2(1'b1),
.I3(CLBLM_R_X7Y114_SLICE_X8Y114_AO6),
.I4(CLBLM_R_X7Y114_SLICE_X8Y114_BO6),
.I5(CLBLM_R_X5Y115_SLICE_X6Y115_BO6),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_BO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h669966992db42db4)
  ) CLBLL_L_X4Y115_SLICE_X5Y115_ALUT (
.I0(CLBLM_R_X5Y116_SLICE_X6Y116_CO6),
.I1(CLBLM_R_X5Y115_SLICE_X6Y115_AO5),
.I2(CLBLM_R_X5Y114_SLICE_X7Y114_AO6),
.I3(CLBLM_R_X7Y114_SLICE_X8Y114_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y115_SLICE_X5Y115_AO5),
.O6(CLBLL_L_X4Y115_SLICE_X5Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y102_SLICE_X10Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y102_SLICE_X10Y102_DO5),
.O6(CLBLM_L_X8Y102_SLICE_X10Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y102_SLICE_X10Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y102_SLICE_X10Y102_CO5),
.O6(CLBLM_L_X8Y102_SLICE_X10Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y102_SLICE_X10Y102_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y102_SLICE_X10Y102_BO5),
.O6(CLBLM_L_X8Y102_SLICE_X10Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd505ffff6a5af000)
  ) CLBLM_L_X8Y102_SLICE_X10Y102_ALUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y102_SLICE_X10Y102_AO5),
.O6(CLBLM_L_X8Y102_SLICE_X10Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y102_SLICE_X11Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y102_SLICE_X11Y102_DO5),
.O6(CLBLM_L_X8Y102_SLICE_X11Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2abfbf2a02abab02)
  ) CLBLM_L_X8Y102_SLICE_X11Y102_CLUT (
.I0(CLBLM_L_X8Y102_SLICE_X11Y102_AO6),
.I1(CLBLM_L_X8Y102_SLICE_X10Y102_AO6),
.I2(CLBLM_L_X10Y103_SLICE_X12Y103_CO6),
.I3(CLBLM_L_X10Y103_SLICE_X12Y103_AO6),
.I4(CLBLM_L_X10Y103_SLICE_X13Y103_BO6),
.I5(CLBLM_R_X7Y102_SLICE_X9Y102_AO5),
.O5(CLBLM_L_X8Y102_SLICE_X11Y102_CO5),
.O6(CLBLM_L_X8Y102_SLICE_X11Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h599aa665a665599a)
  ) CLBLM_L_X8Y102_SLICE_X11Y102_BLUT (
.I0(CLBLM_L_X10Y103_SLICE_X12Y103_AO6),
.I1(CLBLM_R_X7Y102_SLICE_X9Y102_AO5),
.I2(CLBLM_L_X8Y102_SLICE_X10Y102_AO6),
.I3(CLBLM_L_X10Y103_SLICE_X12Y103_CO6),
.I4(CLBLM_L_X8Y102_SLICE_X11Y102_AO6),
.I5(CLBLM_L_X10Y103_SLICE_X13Y103_BO6),
.O5(CLBLM_L_X8Y102_SLICE_X11Y102_BO5),
.O6(CLBLM_L_X8Y102_SLICE_X11Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a088888888)
  ) CLBLM_L_X8Y102_SLICE_X11Y102_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y102_SLICE_X11Y102_AO5),
.O6(CLBLM_L_X8Y102_SLICE_X11Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf770f88077008800)
  ) CLBLM_L_X8Y103_SLICE_X10Y103_DLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(CLBLM_L_X8Y102_SLICE_X11Y102_CO6),
.I4(CLBLM_L_X10Y104_SLICE_X12Y104_CO6),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_L_X8Y103_SLICE_X10Y103_DO5),
.O6(CLBLM_L_X8Y103_SLICE_X10Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd1b72e48953f6ac0)
  ) CLBLM_L_X8Y103_SLICE_X10Y103_CLUT (
.I0(CLBLM_L_X8Y103_SLICE_X10Y103_AO6),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(CLBLM_L_X10Y103_SLICE_X13Y103_AO6),
.I4(CLBLM_L_X10Y104_SLICE_X12Y104_CO6),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_L_X8Y103_SLICE_X10Y103_CO5),
.O6(CLBLM_L_X8Y103_SLICE_X10Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9666999669996669)
  ) CLBLM_L_X8Y103_SLICE_X10Y103_BLUT (
.I0(CLBLM_L_X10Y103_SLICE_X12Y103_DO6),
.I1(CLBLM_L_X10Y103_SLICE_X12Y103_BO6),
.I2(CLBLM_R_X7Y104_SLICE_X8Y104_AO6),
.I3(CLBLM_R_X7Y102_SLICE_X9Y102_CO6),
.I4(CLBLM_L_X8Y102_SLICE_X11Y102_BO6),
.I5(CLBLM_L_X8Y102_SLICE_X11Y102_CO6),
.O5(CLBLM_L_X8Y103_SLICE_X10Y103_BO5),
.O6(CLBLM_L_X8Y103_SLICE_X10Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h08088f8f88778877)
  ) CLBLM_L_X8Y103_SLICE_X10Y103_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(CLBLM_L_X8Y102_SLICE_X10Y102_AO6),
.I3(CLBLM_R_X7Y103_SLICE_X9Y103_AO6),
.I4(CLBLM_L_X10Y103_SLICE_X12Y103_CO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y103_SLICE_X10Y103_AO5),
.O6(CLBLM_L_X8Y103_SLICE_X10Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y103_SLICE_X11Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y103_SLICE_X11Y103_DO5),
.O6(CLBLM_L_X8Y103_SLICE_X11Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y103_SLICE_X11Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y103_SLICE_X11Y103_CO5),
.O6(CLBLM_L_X8Y103_SLICE_X11Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y103_SLICE_X11Y103_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y103_SLICE_X11Y103_BO5),
.O6(CLBLM_L_X8Y103_SLICE_X11Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h66cc96cc96cc9933)
  ) CLBLM_L_X8Y103_SLICE_X11Y103_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(CLBLM_L_X10Y103_SLICE_X13Y103_BO6),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(CLBLM_L_X8Y102_SLICE_X10Y102_AO6),
.I5(CLBLM_L_X10Y103_SLICE_X12Y103_CO6),
.O5(CLBLM_L_X8Y103_SLICE_X11Y103_AO5),
.O6(CLBLM_L_X8Y103_SLICE_X11Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff6c6c6c6c000000)
  ) CLBLM_L_X8Y104_SLICE_X10Y104_DLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(CLBLM_L_X8Y103_SLICE_X10Y103_CO6),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(CLBLM_R_X7Y104_SLICE_X9Y104_AO6),
.O5(CLBLM_L_X8Y104_SLICE_X10Y104_DO5),
.O6(CLBLM_L_X8Y104_SLICE_X10Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h96663ccc6999c333)
  ) CLBLM_L_X8Y104_SLICE_X10Y104_CLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(CLBLM_L_X8Y103_SLICE_X10Y103_CO6),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(CLBLM_R_X7Y104_SLICE_X9Y104_AO6),
.O5(CLBLM_L_X8Y104_SLICE_X10Y104_CO5),
.O6(CLBLM_L_X8Y104_SLICE_X10Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff6f6f6666060600)
  ) CLBLM_L_X8Y104_SLICE_X10Y104_BLUT (
.I0(CLBLM_L_X8Y105_SLICE_X10Y105_AO5),
.I1(CLBLM_L_X10Y104_SLICE_X12Y104_AO6),
.I2(CLBLM_L_X8Y104_SLICE_X11Y104_AO6),
.I3(CLBLM_R_X7Y104_SLICE_X9Y104_AO6),
.I4(CLBLM_L_X8Y105_SLICE_X10Y105_AO6),
.I5(CLBLM_R_X7Y105_SLICE_X8Y105_AO5),
.O5(CLBLM_L_X8Y104_SLICE_X10Y104_BO5),
.O6(CLBLM_L_X8Y104_SLICE_X10Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h9969696666969699)
  ) CLBLM_L_X8Y104_SLICE_X10Y104_ALUT (
.I0(CLBLM_L_X8Y105_SLICE_X10Y105_AO5),
.I1(CLBLM_L_X10Y104_SLICE_X12Y104_AO6),
.I2(CLBLM_L_X8Y104_SLICE_X11Y104_AO6),
.I3(CLBLM_R_X7Y104_SLICE_X9Y104_AO6),
.I4(CLBLM_L_X8Y105_SLICE_X10Y105_AO6),
.I5(CLBLM_R_X7Y105_SLICE_X8Y105_AO5),
.O5(CLBLM_L_X8Y104_SLICE_X10Y104_AO5),
.O6(CLBLM_L_X8Y104_SLICE_X10Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y104_SLICE_X11Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y104_SLICE_X11Y104_DO5),
.O6(CLBLM_L_X8Y104_SLICE_X11Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y104_SLICE_X11Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y104_SLICE_X11Y104_CO5),
.O6(CLBLM_L_X8Y104_SLICE_X11Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y104_SLICE_X11Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y104_SLICE_X11Y104_BO5),
.O6(CLBLM_L_X8Y104_SLICE_X11Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h966669995aaaa555)
  ) CLBLM_L_X8Y104_SLICE_X11Y104_ALUT (
.I0(CLBLM_L_X10Y104_SLICE_X12Y104_CO6),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLM_L_X8Y102_SLICE_X11Y102_CO6),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_L_X8Y104_SLICE_X11Y104_AO5),
.O6(CLBLM_L_X8Y104_SLICE_X11Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y105_SLICE_X10Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y105_SLICE_X10Y105_DO5),
.O6(CLBLM_L_X8Y105_SLICE_X10Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h963c69c369c369c3)
  ) CLBLM_L_X8Y105_SLICE_X10Y105_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(CLBLM_L_X10Y105_SLICE_X13Y105_CO6),
.I2(CLBLM_L_X8Y103_SLICE_X10Y103_DO6),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_L_X8Y105_SLICE_X10Y105_CO5),
.O6(CLBLM_L_X8Y105_SLICE_X10Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4cb3807f26d9ea15)
  ) CLBLM_L_X8Y105_SLICE_X10Y105_BLUT (
.I0(CLBLM_L_X8Y104_SLICE_X10Y104_DO6),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_L_X10Y105_SLICE_X12Y105_BO6),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(CLBLM_L_X8Y105_SLICE_X10Y105_CO6),
.O5(CLBLM_L_X8Y105_SLICE_X10Y105_BO5),
.O6(CLBLM_L_X8Y105_SLICE_X10Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f000f000)
  ) CLBLM_L_X8Y105_SLICE_X10Y105_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y105_SLICE_X10Y105_AO5),
.O6(CLBLM_L_X8Y105_SLICE_X10Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y105_SLICE_X11Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y105_SLICE_X11Y105_DO5),
.O6(CLBLM_L_X8Y105_SLICE_X11Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y105_SLICE_X11Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y105_SLICE_X11Y105_CO5),
.O6(CLBLM_L_X8Y105_SLICE_X11Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y105_SLICE_X11Y105_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y105_SLICE_X11Y105_BO5),
.O6(CLBLM_L_X8Y105_SLICE_X11Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbf2a2a2aea808080)
  ) CLBLM_L_X8Y105_SLICE_X11Y105_ALUT (
.I0(CLBLM_L_X8Y103_SLICE_X10Y103_DO6),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(CLBLM_L_X10Y105_SLICE_X13Y105_CO6),
.O5(CLBLM_L_X8Y105_SLICE_X11Y105_AO5),
.O6(CLBLM_L_X8Y105_SLICE_X11Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y106_SLICE_X10Y106_DO5),
.O6(CLBLM_L_X8Y106_SLICE_X10Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y106_SLICE_X10Y106_CO5),
.O6(CLBLM_L_X8Y106_SLICE_X10Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y106_SLICE_X10Y106_BO5),
.O6(CLBLM_L_X8Y106_SLICE_X10Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y106_SLICE_X10Y106_AO5),
.O6(CLBLM_L_X8Y106_SLICE_X10Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y106_SLICE_X11Y106_DO5),
.O6(CLBLM_L_X8Y106_SLICE_X11Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y106_SLICE_X11Y106_CO5),
.O6(CLBLM_L_X8Y106_SLICE_X11Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hadd5077f522af880)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(CLBLM_L_X8Y105_SLICE_X11Y105_AO6),
.I3(CLBLM_L_X10Y106_SLICE_X12Y106_AO6),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(CLBLM_L_X10Y106_SLICE_X12Y106_CO6),
.O5(CLBLM_L_X8Y106_SLICE_X11Y106_BO5),
.O6(CLBLM_L_X8Y106_SLICE_X11Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f000f000)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y106_SLICE_X11Y106_AO5),
.O6(CLBLM_L_X8Y106_SLICE_X11Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heb828282bb222222)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_DLUT (
.I0(CLBLM_R_X7Y106_SLICE_X9Y106_AO6),
.I1(CLBLM_L_X8Y105_SLICE_X10Y105_BO6),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_L_X8Y107_SLICE_X10Y107_DO5),
.O6(CLBLM_L_X8Y107_SLICE_X10Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33c3cc36996)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_CLUT (
.I0(CLBLM_L_X8Y106_SLICE_X11Y106_AO6),
.I1(CLBLM_L_X10Y105_SLICE_X13Y105_BO6),
.I2(CLBLM_L_X8Y107_SLICE_X11Y107_AO6),
.I3(CLBLM_L_X8Y104_SLICE_X10Y104_BO6),
.I4(CLBLM_R_X7Y105_SLICE_X8Y105_CO6),
.I5(CLBLM_L_X8Y104_SLICE_X10Y104_AO6),
.O5(CLBLM_L_X8Y107_SLICE_X10Y107_CO5),
.O6(CLBLM_L_X8Y107_SLICE_X10Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33ca55a0ff0)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(CLBLM_R_X7Y106_SLICE_X9Y106_AO6),
.I3(CLBLM_L_X8Y105_SLICE_X10Y105_BO6),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_L_X8Y107_SLICE_X10Y107_BO5),
.O6(CLBLM_L_X8Y107_SLICE_X10Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h965a3cf069a5c30f)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(CLBLM_L_X8Y104_SLICE_X10Y104_BO6),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLM_L_X10Y105_SLICE_X12Y105_BO6),
.O5(CLBLM_L_X8Y107_SLICE_X10Y107_AO5),
.O6(CLBLM_L_X8Y107_SLICE_X10Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9696966996696969)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_DLUT (
.I0(CLBLM_L_X10Y106_SLICE_X13Y106_CO6),
.I1(CLBLM_L_X8Y106_SLICE_X11Y106_AO5),
.I2(CLBLM_L_X10Y108_SLICE_X13Y108_CO6),
.I3(CLBLM_L_X8Y107_SLICE_X11Y107_AO5),
.I4(CLBLM_L_X10Y105_SLICE_X13Y105_DO6),
.I5(CLBLM_L_X10Y106_SLICE_X13Y106_BO6),
.O5(CLBLM_L_X8Y107_SLICE_X11Y107_DO5),
.O6(CLBLM_L_X8Y107_SLICE_X11Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8e71718e718e8e71)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_CLUT (
.I0(CLBLM_L_X8Y107_SLICE_X11Y107_AO6),
.I1(CLBLM_L_X8Y104_SLICE_X10Y104_BO6),
.I2(CLBLM_L_X10Y105_SLICE_X13Y105_BO6),
.I3(CLBLM_L_X8Y107_SLICE_X11Y107_AO5),
.I4(CLBLM_L_X10Y105_SLICE_X13Y105_DO6),
.I5(CLBLM_L_X10Y106_SLICE_X13Y106_BO6),
.O5(CLBLM_L_X8Y107_SLICE_X11Y107_CO5),
.O6(CLBLM_L_X8Y107_SLICE_X11Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7707070f8808080)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(CLBLM_L_X8Y104_SLICE_X10Y104_BO6),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_L_X10Y105_SLICE_X12Y105_BO6),
.O5(CLBLM_L_X8Y107_SLICE_X11Y107_BO5),
.O6(CLBLM_L_X8Y107_SLICE_X11Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00aa00aa00)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(1'b1),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y107_SLICE_X11Y107_AO5),
.O6(CLBLM_L_X8Y107_SLICE_X11Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he88ec00cfccfe88e)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_DLUT (
.I0(CLBLM_L_X8Y108_SLICE_X10Y108_AO6),
.I1(CLBLM_L_X8Y109_SLICE_X11Y109_AO5),
.I2(CLBLM_L_X8Y107_SLICE_X11Y107_CO6),
.I3(CLBLM_L_X8Y108_SLICE_X10Y108_AO5),
.I4(CLBLM_R_X7Y106_SLICE_X9Y106_AO6),
.I5(CLBLM_L_X8Y107_SLICE_X10Y107_AO6),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_DO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33c3cc36996)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_CLUT (
.I0(CLBLM_L_X8Y108_SLICE_X10Y108_AO6),
.I1(CLBLM_L_X8Y109_SLICE_X11Y109_AO5),
.I2(CLBLM_L_X8Y107_SLICE_X11Y107_CO6),
.I3(CLBLM_L_X8Y108_SLICE_X10Y108_AO5),
.I4(CLBLM_R_X7Y106_SLICE_X9Y106_AO6),
.I5(CLBLM_L_X8Y107_SLICE_X10Y107_AO6),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_CO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h695aa56996a55a96)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_BLUT (
.I0(CLBLM_L_X8Y107_SLICE_X11Y107_BO6),
.I1(CLBLM_R_X7Y106_SLICE_X9Y106_AO6),
.I2(CLBLM_L_X8Y108_SLICE_X11Y108_AO6),
.I3(CLBLM_L_X8Y107_SLICE_X10Y107_AO6),
.I4(CLBLM_L_X8Y108_SLICE_X10Y108_AO6),
.I5(CLBLM_L_X8Y108_SLICE_X10Y108_AO5),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_BO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0f0f00000)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(1'b1),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_AO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd444e888fcccc000)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_DLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(CLBLM_L_X10Y105_SLICE_X13Y105_DO6),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(CLBLM_L_X10Y106_SLICE_X12Y106_CO6),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_DO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h965a66aa69a59955)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_CLUT (
.I0(CLBLM_L_X8Y106_SLICE_X11Y106_BO6),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(CLBLM_L_X8Y107_SLICE_X11Y107_BO6),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_CO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7f8708070807080)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(CLBLM_L_X8Y107_SLICE_X11Y107_BO6),
.I3(CLBLM_L_X8Y106_SLICE_X11Y106_BO6),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(RIOB33_X105Y101_IOB_X1Y102_I),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_BO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h9669696966999999)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_ALUT (
.I0(CLBLM_L_X10Y106_SLICE_X12Y106_CO6),
.I1(CLBLM_L_X10Y105_SLICE_X13Y105_DO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_AO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd24b2db42db4d24b)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_DLUT (
.I0(CLBLM_L_X8Y108_SLICE_X11Y108_AO6),
.I1(CLBLM_L_X8Y108_SLICE_X10Y108_AO5),
.I2(CLBLM_L_X8Y107_SLICE_X11Y107_DO6),
.I3(CLBLM_L_X8Y107_SLICE_X11Y107_BO6),
.I4(CLBLM_R_X7Y109_SLICE_X8Y109_AO5),
.I5(CLBLM_L_X8Y109_SLICE_X11Y109_AO6),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_DO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996669999666996)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_CLUT (
.I0(CLBLM_L_X8Y109_SLICE_X10Y109_AO6),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_AO5),
.I2(CLBLM_L_X8Y108_SLICE_X10Y108_DO6),
.I3(CLBLM_L_X10Y109_SLICE_X12Y109_BO6),
.I4(CLBLM_L_X8Y109_SLICE_X10Y109_DO6),
.I5(CLBLM_R_X5Y109_SLICE_X7Y109_AO5),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_CO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h639cc6399c6339c6)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_BLUT (
.I0(CLBLM_L_X8Y107_SLICE_X10Y107_DO6),
.I1(CLBLM_L_X8Y109_SLICE_X11Y109_BO6),
.I2(CLBLM_L_X8Y108_SLICE_X11Y108_CO6),
.I3(CLBLM_L_X8Y108_SLICE_X11Y108_BO6),
.I4(CLBLM_L_X8Y109_SLICE_X11Y109_AO5),
.I5(CLBLM_L_X8Y109_SLICE_X11Y109_AO6),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_BO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf45ef8a5d04ae08)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_ALUT (
.I0(CLBLM_R_X7Y109_SLICE_X8Y109_AO5),
.I1(CLBLM_L_X8Y107_SLICE_X11Y107_BO6),
.I2(CLBLM_L_X8Y108_SLICE_X11Y108_AO6),
.I3(CLBLM_L_X8Y109_SLICE_X11Y109_AO6),
.I4(CLBLM_L_X8Y107_SLICE_X11Y107_DO6),
.I5(CLBLM_L_X8Y108_SLICE_X10Y108_AO5),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_AO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_DO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd444fccce888c000)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLM_L_X8Y108_SLICE_X11Y108_DO6),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(CLBLM_R_X11Y109_SLICE_X14Y109_AO6),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_CO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h966966993cc3cc33)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(CLBLM_L_X8Y108_SLICE_X11Y108_DO6),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(CLBLM_R_X11Y109_SLICE_X14Y109_AO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_BO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000aa00aa00)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_AO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_DO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_CO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9669699666999966)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_BLUT (
.I0(CLBLM_L_X8Y108_SLICE_X11Y108_BO6),
.I1(CLBLM_L_X8Y109_SLICE_X11Y109_BO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(CLBLM_L_X8Y108_SLICE_X10Y108_DO6),
.I4(CLBLM_L_X8Y109_SLICE_X11Y109_AO6),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_BO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000ff000000)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(1'b1),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_AO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfae0800080800000)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_DLUT (
.I0(CLBLM_L_X12Y110_SLICE_X17Y110_AO6),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(RIOB33_X105Y111_IOB_X1Y111_I),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_DO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff7fffffffffff)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_CLUT (
.I0(CLBLM_R_X7Y107_SLICE_X8Y107_BO6),
.I1(CLBLM_L_X10Y110_SLICE_X13Y110_BO6),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(CLBLM_L_X10Y111_SLICE_X13Y111_AO6),
.I5(CLBLM_R_X11Y110_SLICE_X15Y110_DO6),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_CO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff7fffffff)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X11Y109_SLICE_X14Y109_AO6),
.I3(CLBLM_L_X10Y108_SLICE_X13Y108_DO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_BO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc000066aa66aa)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_ALUT (
.I0(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(1'b1),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_AO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a95956a956a6a95)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_DLUT (
.I0(CLBLM_L_X8Y109_SLICE_X10Y109_AO6),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_L_X10Y110_SLICE_X13Y110_CO6),
.I4(CLBLM_L_X10Y112_SLICE_X12Y112_AO6),
.I5(CLBLM_L_X8Y109_SLICE_X11Y109_CO6),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_DO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff69690069006900)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_CLUT (
.I0(CLBLM_L_X8Y109_SLICE_X11Y109_BO6),
.I1(CLBLM_L_X8Y109_SLICE_X11Y109_AO6),
.I2(CLBLM_L_X8Y108_SLICE_X11Y108_BO6),
.I3(CLBLM_L_X8Y108_SLICE_X10Y108_DO6),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_CO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h956aa9566a9556a9)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_BLUT (
.I0(CLBLM_L_X10Y112_SLICE_X12Y112_AO6),
.I1(CLBLM_L_X8Y108_SLICE_X11Y108_BO6),
.I2(CLBLM_L_X8Y109_SLICE_X11Y109_AO6),
.I3(CLBLM_L_X10Y110_SLICE_X13Y110_CO6),
.I4(CLBLM_L_X8Y109_SLICE_X11Y109_BO6),
.I5(CLBLM_L_X8Y109_SLICE_X11Y109_CO6),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_BO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he8d4a050d4e850a0)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_ALUT (
.I0(CLBLM_L_X10Y112_SLICE_X12Y112_AO6),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(CLBLM_L_X8Y109_SLICE_X10Y109_AO6),
.I3(CLBLM_L_X10Y110_SLICE_X13Y110_CO6),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLM_L_X8Y109_SLICE_X11Y109_CO6),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_AO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbba2b300aa202000)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_DLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(CLBLM_R_X11Y111_SLICE_X14Y111_CO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(CLBLM_L_X8Y111_SLICE_X11Y111_AO5),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(CLBLM_R_X11Y111_SLICE_X14Y111_AO5),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_DO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8f70e31c7f8013ec)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_CLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(CLBLM_R_X11Y111_SLICE_X14Y111_AO5),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(CLBLM_R_X11Y111_SLICE_X14Y111_AO6),
.I4(CLBLM_R_X11Y111_SLICE_X14Y111_CO6),
.I5(RIOB33_X105Y107_IOB_X1Y108_I),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_CO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00000096965a5a)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_BLUT (
.I0(CLBLM_L_X10Y111_SLICE_X13Y111_CO6),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(CLBLM_R_X11Y111_SLICE_X14Y111_DO6),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_BO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00003cf03cf0)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(CLBLM_R_X11Y111_SLICE_X14Y111_AO6),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_AO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hde5a4800eeaa8800)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_DLUT (
.I0(CLBLM_L_X10Y111_SLICE_X12Y111_AO6),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(CLBLM_L_X10Y112_SLICE_X12Y112_DO6),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_DO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb2e82288e8e88888)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_CLUT (
.I0(CLBLM_L_X8Y111_SLICE_X10Y111_AO6),
.I1(CLBLM_L_X8Y112_SLICE_X11Y112_AO6),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_CO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4d17dd7744114d17)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_BLUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_AO5),
.I1(CLBLM_L_X10Y110_SLICE_X12Y110_BO6),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_AO6),
.I3(CLBLM_R_X5Y111_SLICE_X6Y111_AO5),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_AO6),
.I5(CLBLM_L_X10Y112_SLICE_X12Y112_BO6),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_BO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6966996996996696)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_ALUT (
.I0(CLBLM_R_X5Y112_SLICE_X6Y112_AO5),
.I1(CLBLM_L_X8Y113_SLICE_X11Y113_BO6),
.I2(CLBLM_L_X8Y113_SLICE_X11Y113_AO6),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_BO6),
.I4(CLBLM_R_X7Y113_SLICE_X9Y113_AO6),
.I5(CLBLM_R_X7Y113_SLICE_X9Y113_CO6),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_AO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_DO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_CO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_BO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969699669969696)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_ALUT (
.I0(CLBLM_L_X10Y112_SLICE_X12Y112_AO5),
.I1(CLBLM_L_X10Y110_SLICE_X13Y110_BO6),
.I2(CLBLM_L_X10Y111_SLICE_X13Y111_AO6),
.I3(CLBLM_L_X10Y112_SLICE_X12Y112_AO6),
.I4(CLBLM_L_X10Y110_SLICE_X13Y110_CO6),
.I5(CLBLM_L_X8Y109_SLICE_X11Y109_CO6),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_AO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h966969695aa5a5a5)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_DLUT (
.I0(CLBLM_L_X10Y111_SLICE_X12Y111_AO6),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(CLBLM_L_X10Y112_SLICE_X12Y112_DO6),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_DO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h099900099fff999f)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_CLUT (
.I0(CLBLM_L_X8Y114_SLICE_X10Y114_AO6),
.I1(CLBLM_L_X8Y113_SLICE_X11Y113_CO6),
.I2(CLBLM_L_X8Y112_SLICE_X10Y112_CO6),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_AO5),
.I4(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.I5(CLBLM_R_X7Y113_SLICE_X9Y113_AO6),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_CO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h18e79c63d42b50af)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_BLUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(CLBLM_L_X8Y112_SLICE_X10Y112_CO6),
.I3(CLBLM_L_X8Y113_SLICE_X11Y113_CO6),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_BO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha55a5a5aff000000)
  ) CLBLM_L_X8Y113_SLICE_X10Y113_ALUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_DO6),
.I1(1'b1),
.I2(CLBLM_L_X8Y112_SLICE_X10Y112_CO6),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y113_SLICE_X10Y113_AO5),
.O6(CLBLM_L_X8Y113_SLICE_X10Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h63c6cc999c39cc99)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_DLUT (
.I0(CLBLM_L_X10Y112_SLICE_X13Y112_DO6),
.I1(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y113_SLICE_X12Y113_AO5),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(RIOB33_X105Y107_IOB_X1Y107_I),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_DO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc369966996c33c)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_CLUT (
.I0(CLBLM_L_X10Y112_SLICE_X13Y112_BO6),
.I1(CLBLM_L_X10Y112_SLICE_X12Y112_CO6),
.I2(CLBLM_L_X10Y112_SLICE_X13Y112_CO6),
.I3(CLBLM_R_X7Y114_SLICE_X9Y114_AO6),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_AO5),
.I5(CLBLM_L_X10Y112_SLICE_X12Y112_DO6),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_CO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h044ccddf0113377f)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_BLUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_AO5),
.I1(CLBLM_L_X10Y113_SLICE_X12Y113_BO6),
.I2(CLBLM_L_X10Y112_SLICE_X12Y112_DO6),
.I3(CLBLM_L_X10Y112_SLICE_X13Y112_BO6),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_AO6),
.I5(CLBLM_R_X7Y114_SLICE_X9Y114_AO6),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_BO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h366cc993c993366c)
  ) CLBLM_L_X8Y113_SLICE_X11Y113_ALUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_AO5),
.I1(CLBLM_L_X10Y113_SLICE_X12Y113_BO6),
.I2(CLBLM_L_X10Y112_SLICE_X12Y112_DO6),
.I3(CLBLM_L_X10Y112_SLICE_X13Y112_BO6),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_AO6),
.I5(CLBLM_R_X7Y114_SLICE_X9Y114_AO6),
.O5(CLBLM_L_X8Y113_SLICE_X11Y113_AO5),
.O6(CLBLM_L_X8Y113_SLICE_X11Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_DO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdcc4d44454405000)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_CLUT (
.I0(CLBLM_R_X7Y113_SLICE_X9Y113_BO6),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(CLBLM_L_X10Y112_SLICE_X12Y112_CO6),
.I3(CLBLM_L_X10Y112_SLICE_X13Y112_CO6),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_CO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc33c33cc0ff0ff00)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y114_SLICE_X10Y114_CO6),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(CLBLM_L_X8Y113_SLICE_X11Y113_DO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_BO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c088888888)
  ) CLBLM_L_X8Y114_SLICE_X10Y114_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y114_SLICE_X10Y114_AO5),
.O6(CLBLM_L_X8Y114_SLICE_X10Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_DO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_CO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_BO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y114_SLICE_X11Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y114_SLICE_X11Y114_AO5),
.O6(CLBLM_L_X8Y114_SLICE_X11Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2bd4d42bd42b2bd4)
  ) CLBLM_L_X10Y103_SLICE_X12Y103_DLUT (
.I0(CLBLM_L_X10Y103_SLICE_X12Y103_CO5),
.I1(CLBLM_R_X11Y104_SLICE_X14Y104_AO5),
.I2(CLBLM_L_X10Y103_SLICE_X12Y103_AO6),
.I3(CLBLM_L_X10Y103_SLICE_X12Y103_AO5),
.I4(CLBLM_L_X8Y102_SLICE_X11Y102_AO5),
.I5(CLBLM_L_X10Y104_SLICE_X12Y104_DO6),
.O5(CLBLM_L_X10Y103_SLICE_X12Y103_DO5),
.O6(CLBLM_L_X10Y103_SLICE_X12Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h64a8e428b3f733f7)
  ) CLBLM_L_X10Y103_SLICE_X12Y103_CLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y103_SLICE_X12Y103_CO5),
.O6(CLBLM_L_X10Y103_SLICE_X12Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aa00aa00)
  ) CLBLM_L_X10Y103_SLICE_X12Y103_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(1'b1),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y103_SLICE_X12Y103_BO5),
.O6(CLBLM_L_X10Y103_SLICE_X12Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc0088888888)
  ) CLBLM_L_X10Y103_SLICE_X12Y103_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(1'b1),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y103_SLICE_X12Y103_AO5),
.O6(CLBLM_L_X10Y103_SLICE_X12Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y103_SLICE_X13Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y103_SLICE_X13Y103_DO5),
.O6(CLBLM_L_X10Y103_SLICE_X13Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y103_SLICE_X13Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y103_SLICE_X13Y103_CO5),
.O6(CLBLM_L_X10Y103_SLICE_X13Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcaaaf3f3c5653f3f)
  ) CLBLM_L_X10Y103_SLICE_X13Y103_BLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_L_X10Y103_SLICE_X13Y103_BO5),
.O6(CLBLM_L_X10Y103_SLICE_X13Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ccff007171f5f5)
  ) CLBLM_L_X10Y103_SLICE_X13Y103_ALUT (
.I0(CLBLM_R_X11Y104_SLICE_X14Y104_AO5),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(CLBLM_L_X10Y103_SLICE_X12Y103_CO5),
.I3(CLBLM_L_X10Y103_SLICE_X13Y103_BO6),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y103_SLICE_X13Y103_AO5),
.O6(CLBLM_L_X10Y103_SLICE_X13Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hacccff55a63355ff)
  ) CLBLM_L_X10Y104_SLICE_X12Y104_DLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y107_IOB_X1Y108_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y104_SLICE_X12Y104_DO5),
.O6(CLBLM_L_X10Y104_SLICE_X12Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he62a19d573bf8c40)
  ) CLBLM_L_X10Y104_SLICE_X12Y104_CLUT (
.I0(CLBLM_L_X10Y103_SLICE_X12Y103_CO5),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y104_SLICE_X12Y104_DO6),
.I5(CLBLM_R_X11Y104_SLICE_X14Y104_AO5),
.O5(CLBLM_L_X10Y104_SLICE_X12Y104_CO5),
.O6(CLBLM_L_X10Y104_SLICE_X12Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h099900099fff999f)
  ) CLBLM_L_X10Y104_SLICE_X12Y104_BLUT (
.I0(CLBLM_L_X10Y104_SLICE_X12Y104_DO6),
.I1(CLBLM_L_X10Y103_SLICE_X12Y103_AO5),
.I2(CLBLM_L_X10Y103_SLICE_X12Y103_AO6),
.I3(CLBLM_R_X11Y104_SLICE_X14Y104_AO5),
.I4(CLBLM_L_X10Y103_SLICE_X12Y103_CO5),
.I5(CLBLM_L_X8Y102_SLICE_X11Y102_AO5),
.O5(CLBLM_L_X10Y104_SLICE_X12Y104_BO5),
.O6(CLBLM_L_X10Y104_SLICE_X12Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he11e87781ee17887)
  ) CLBLM_L_X10Y104_SLICE_X12Y104_ALUT (
.I0(CLBLM_L_X10Y103_SLICE_X12Y103_DO6),
.I1(CLBLM_L_X8Y102_SLICE_X11Y102_CO6),
.I2(CLBLM_L_X10Y104_SLICE_X13Y104_CO6),
.I3(CLBLM_L_X10Y104_SLICE_X12Y104_BO6),
.I4(CLBLM_L_X10Y103_SLICE_X12Y103_BO6),
.I5(CLBLM_L_X10Y103_SLICE_X12Y103_BO5),
.O5(CLBLM_L_X10Y104_SLICE_X12Y104_AO5),
.O6(CLBLM_L_X10Y104_SLICE_X12Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h44d41171d4dd7177)
  ) CLBLM_L_X10Y104_SLICE_X13Y104_DLUT (
.I0(CLBLM_L_X10Y104_SLICE_X13Y104_AO6),
.I1(CLBLM_L_X10Y106_SLICE_X13Y106_AO6),
.I2(CLBLM_R_X11Y104_SLICE_X14Y104_AO6),
.I3(CLBLM_R_X11Y105_SLICE_X15Y105_AO5),
.I4(CLBLM_R_X7Y111_SLICE_X9Y111_AO6),
.I5(CLBLM_L_X10Y103_SLICE_X12Y103_AO5),
.O5(CLBLM_L_X10Y104_SLICE_X13Y104_DO5),
.O6(CLBLM_L_X10Y104_SLICE_X13Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93936c36c9c936)
  ) CLBLM_L_X10Y104_SLICE_X13Y104_CLUT (
.I0(CLBLM_L_X10Y103_SLICE_X12Y103_AO5),
.I1(CLBLM_L_X10Y106_SLICE_X13Y106_AO6),
.I2(CLBLM_R_X11Y105_SLICE_X15Y105_AO5),
.I3(CLBLM_R_X7Y111_SLICE_X9Y111_AO6),
.I4(CLBLM_L_X10Y104_SLICE_X13Y104_AO6),
.I5(CLBLM_R_X11Y104_SLICE_X14Y104_AO6),
.O5(CLBLM_L_X10Y104_SLICE_X13Y104_CO5),
.O6(CLBLM_L_X10Y104_SLICE_X13Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3ccc3ccc5fff0555)
  ) CLBLM_L_X10Y104_SLICE_X13Y104_BLUT (
.I0(CLBLM_R_X11Y105_SLICE_X15Y105_AO5),
.I1(CLBLM_L_X10Y104_SLICE_X12Y104_DO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(CLBLM_R_X11Y104_SLICE_X14Y104_AO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y104_SLICE_X13Y104_BO5),
.O6(CLBLM_L_X10Y104_SLICE_X13Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000aa00aa00)
  ) CLBLM_L_X10Y104_SLICE_X13Y104_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(1'b1),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y104_SLICE_X13Y104_AO5),
.O6(CLBLM_L_X10Y104_SLICE_X13Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2db4d24bd24b2db4)
  ) CLBLM_L_X10Y105_SLICE_X12Y105_DLUT (
.I0(CLBLM_L_X10Y104_SLICE_X12Y104_BO6),
.I1(CLBLM_L_X10Y103_SLICE_X12Y103_BO5),
.I2(CLBLM_L_X10Y104_SLICE_X13Y104_AO5),
.I3(CLBLM_L_X10Y104_SLICE_X13Y104_CO6),
.I4(CLBLM_R_X11Y105_SLICE_X14Y105_DO6),
.I5(CLBLM_L_X10Y104_SLICE_X13Y104_DO6),
.O5(CLBLM_L_X10Y105_SLICE_X12Y105_DO5),
.O6(CLBLM_L_X10Y105_SLICE_X12Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9669696966999999)
  ) CLBLM_L_X10Y105_SLICE_X12Y105_CLUT (
.I0(CLBLM_L_X10Y104_SLICE_X12Y104_BO6),
.I1(CLBLM_L_X10Y105_SLICE_X13Y105_AO6),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_L_X10Y105_SLICE_X12Y105_CO5),
.O6(CLBLM_L_X10Y105_SLICE_X12Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he51a8f7015ea7f80)
  ) CLBLM_L_X10Y105_SLICE_X12Y105_BLUT (
.I0(CLBLM_L_X8Y103_SLICE_X10Y103_DO6),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(CLBLM_L_X10Y105_SLICE_X12Y105_DO6),
.I4(CLBLM_L_X10Y105_SLICE_X12Y105_CO6),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_L_X10Y105_SLICE_X12Y105_BO5),
.O6(CLBLM_L_X10Y105_SLICE_X12Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb73f2103ffffa50f)
  ) CLBLM_L_X10Y105_SLICE_X12Y105_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(CLBLM_L_X10Y105_SLICE_X13Y105_AO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y104_SLICE_X12Y104_BO6),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_L_X10Y105_SLICE_X12Y105_AO5),
.O6(CLBLM_L_X10Y105_SLICE_X12Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haf8e8e0afae8e8a0)
  ) CLBLM_L_X10Y105_SLICE_X13Y105_DLUT (
.I0(CLBLM_R_X11Y105_SLICE_X15Y105_BO5),
.I1(CLBLM_L_X10Y105_SLICE_X12Y105_CO6),
.I2(CLBLM_L_X10Y105_SLICE_X12Y105_DO6),
.I3(CLBLM_L_X8Y105_SLICE_X10Y105_AO5),
.I4(CLBLM_L_X8Y103_SLICE_X10Y103_DO6),
.I5(CLBLM_L_X10Y109_SLICE_X12Y109_AO5),
.O5(CLBLM_L_X10Y105_SLICE_X13Y105_DO5),
.O6(CLBLM_L_X10Y105_SLICE_X13Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha96959996a5a9aaa)
  ) CLBLM_L_X10Y105_SLICE_X13Y105_CLUT (
.I0(CLBLM_L_X10Y105_SLICE_X13Y105_AO6),
.I1(CLBLM_L_X10Y103_SLICE_X13Y103_AO5),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X10Y104_SLICE_X13Y104_BO6),
.O5(CLBLM_L_X10Y105_SLICE_X13Y105_CO5),
.O6(CLBLM_L_X10Y105_SLICE_X13Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc93636c9936c6c93)
  ) CLBLM_L_X10Y105_SLICE_X13Y105_BLUT (
.I0(CLBLM_L_X8Y103_SLICE_X10Y103_DO6),
.I1(CLBLM_L_X10Y105_SLICE_X12Y105_DO6),
.I2(CLBLM_L_X10Y105_SLICE_X12Y105_CO6),
.I3(CLBLM_L_X10Y109_SLICE_X12Y109_AO5),
.I4(CLBLM_R_X11Y105_SLICE_X15Y105_BO5),
.I5(CLBLM_L_X8Y105_SLICE_X10Y105_AO5),
.O5(CLBLM_L_X10Y105_SLICE_X13Y105_BO5),
.O6(CLBLM_L_X10Y105_SLICE_X13Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8ef5710a71f58e0a)
  ) CLBLM_L_X10Y105_SLICE_X13Y105_ALUT (
.I0(CLBLM_R_X11Y105_SLICE_X15Y105_AO5),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X11Y104_SLICE_X14Y104_AO6),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(CLBLM_L_X10Y106_SLICE_X13Y106_AO6),
.I5(RIOB33_X105Y107_IOB_X1Y107_I),
.O5(CLBLM_L_X10Y105_SLICE_X13Y105_AO5),
.O6(CLBLM_L_X10Y105_SLICE_X13Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h96695aa53cc3f00f)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(CLBLM_L_X10Y104_SLICE_X13Y104_DO6),
.I3(CLBLM_R_X11Y105_SLICE_X15Y105_CO6),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_L_X10Y106_SLICE_X12Y106_DO5),
.O6(CLBLM_L_X10Y106_SLICE_X12Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2dd2b44bd22d4bb4)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_CLUT (
.I0(CLBLM_L_X10Y105_SLICE_X12Y105_AO6),
.I1(CLBLM_L_X10Y109_SLICE_X12Y109_AO5),
.I2(CLBLM_L_X10Y108_SLICE_X13Y108_AO5),
.I3(CLBLM_R_X11Y106_SLICE_X14Y106_BO6),
.I4(CLBLM_L_X10Y106_SLICE_X12Y106_DO6),
.I5(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.O5(CLBLM_L_X10Y106_SLICE_X12Y106_CO5),
.O6(CLBLM_L_X10Y106_SLICE_X12Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h80eaeaea2abfbfbf)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_BLUT (
.I0(CLBLM_L_X10Y104_SLICE_X13Y104_DO6),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X11Y105_SLICE_X15Y105_CO6),
.O5(CLBLM_L_X10Y106_SLICE_X12Y106_BO5),
.O6(CLBLM_L_X10Y106_SLICE_X12Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h965a69a569a569a5)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_ALUT (
.I0(CLBLM_R_X11Y105_SLICE_X14Y105_CO6),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(CLBLM_L_X10Y105_SLICE_X12Y105_AO6),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_L_X10Y106_SLICE_X12Y106_AO5),
.O6(CLBLM_L_X10Y106_SLICE_X12Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5695a96695a96a5)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_DLUT (
.I0(CLBLM_R_X11Y105_SLICE_X14Y105_BO6),
.I1(CLBLM_L_X10Y104_SLICE_X13Y104_AO5),
.I2(CLBLM_R_X11Y107_SLICE_X14Y107_DO6),
.I3(CLBLM_L_X10Y104_SLICE_X13Y104_DO6),
.I4(CLBLM_L_X8Y110_SLICE_X11Y110_AO6),
.I5(CLBLM_R_X11Y105_SLICE_X14Y105_DO6),
.O5(CLBLM_L_X10Y106_SLICE_X13Y106_DO5),
.O6(CLBLM_L_X10Y106_SLICE_X13Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3b02023bbf2323bf)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_CLUT (
.I0(CLBLM_L_X10Y105_SLICE_X12Y105_AO6),
.I1(CLBLM_L_X10Y107_SLICE_X13Y107_AO5),
.I2(CLBLM_L_X10Y109_SLICE_X12Y109_AO5),
.I3(CLBLM_L_X10Y108_SLICE_X13Y108_AO5),
.I4(CLBLM_L_X10Y106_SLICE_X13Y106_DO6),
.I5(CLBLM_L_X10Y106_SLICE_X12Y106_DO6),
.O5(CLBLM_L_X10Y106_SLICE_X13Y106_CO5),
.O6(CLBLM_L_X10Y106_SLICE_X13Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a55a69965aa596)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_BLUT (
.I0(CLBLM_L_X10Y106_SLICE_X13Y106_DO6),
.I1(CLBLM_L_X10Y109_SLICE_X12Y109_AO5),
.I2(CLBLM_L_X10Y108_SLICE_X13Y108_AO5),
.I3(CLBLM_L_X10Y106_SLICE_X12Y106_DO6),
.I4(CLBLM_L_X10Y105_SLICE_X12Y105_AO6),
.I5(CLBLM_L_X10Y107_SLICE_X13Y107_AO5),
.O5(CLBLM_L_X10Y106_SLICE_X13Y106_BO5),
.O6(CLBLM_L_X10Y106_SLICE_X13Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he2d2aa55ff0f0fff)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_ALUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(RIOB33_X105Y113_IOB_X1Y113_I),
.O5(CLBLM_L_X10Y106_SLICE_X13Y106_AO5),
.O6(CLBLM_L_X10Y106_SLICE_X13Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y107_SLICE_X12Y107_DO5),
.O6(CLBLM_L_X10Y107_SLICE_X12Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf03c3cf08c40cc00)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_CLUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O5(CLBLM_L_X10Y107_SLICE_X12Y107_CO5),
.O6(CLBLM_L_X10Y107_SLICE_X12Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hecece8a0c8800000)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_BLUT (
.I0(CLBLM_L_X10Y110_SLICE_X13Y110_AO5),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(CLBLM_R_X11Y107_SLICE_X14Y107_BO5),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLM_L_X10Y107_SLICE_X12Y107_CO6),
.O5(CLBLM_L_X10Y107_SLICE_X12Y107_BO5),
.O6(CLBLM_L_X10Y107_SLICE_X12Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdb93175f246ce8a0)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_ALUT (
.I0(CLBLM_L_X10Y110_SLICE_X13Y110_AO5),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(CLBLM_R_X11Y107_SLICE_X14Y107_BO5),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLM_L_X10Y107_SLICE_X12Y107_CO6),
.O5(CLBLM_L_X10Y107_SLICE_X12Y107_AO5),
.O6(CLBLM_L_X10Y107_SLICE_X12Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfec88888ec800000)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_DLUT (
.I0(CLBLM_R_X11Y108_SLICE_X15Y108_AO6),
.I1(CLBLM_R_X11Y109_SLICE_X15Y109_AO6),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(CLBLM_R_X11Y107_SLICE_X14Y107_AO6),
.O5(CLBLM_L_X10Y107_SLICE_X13Y107_DO5),
.O6(CLBLM_L_X10Y107_SLICE_X13Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h36c999996c933333)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_CLUT (
.I0(CLBLM_R_X11Y108_SLICE_X15Y108_AO6),
.I1(CLBLM_R_X11Y109_SLICE_X15Y109_AO6),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(CLBLM_R_X11Y107_SLICE_X14Y107_AO6),
.O5(CLBLM_L_X10Y107_SLICE_X13Y107_CO5),
.O6(CLBLM_L_X10Y107_SLICE_X13Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699699669969966)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_BLUT (
.I0(CLBLM_L_X10Y107_SLICE_X12Y107_AO6),
.I1(CLBLM_L_X8Y111_SLICE_X11Y111_BO6),
.I2(CLBLM_R_X11Y105_SLICE_X14Y105_BO6),
.I3(CLBLM_R_X11Y107_SLICE_X14Y107_CO6),
.I4(CLBLM_L_X8Y110_SLICE_X11Y110_AO6),
.I5(CLBLM_R_X11Y107_SLICE_X14Y107_DO6),
.O5(CLBLM_L_X10Y107_SLICE_X13Y107_BO5),
.O6(CLBLM_L_X10Y107_SLICE_X13Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000cc00cc00)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(1'b1),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y107_SLICE_X13Y107_AO5),
.O6(CLBLM_L_X10Y107_SLICE_X13Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000000000)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(RIOB33_X105Y109_IOB_X1Y109_I),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_DO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2dd2b44bd22d4bb4)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_CLUT (
.I0(CLBLM_L_X10Y106_SLICE_X13Y106_CO6),
.I1(CLBLM_L_X8Y106_SLICE_X11Y106_AO5),
.I2(CLBLM_L_X10Y108_SLICE_X13Y108_BO6),
.I3(CLBLM_L_X10Y108_SLICE_X12Y108_AO5),
.I4(CLBLM_L_X10Y108_SLICE_X13Y108_CO6),
.I5(CLBLM_R_X11Y108_SLICE_X14Y108_DO6),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_CO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h956a6a95a95656a9)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_BLUT (
.I0(CLBLM_R_X11Y109_SLICE_X15Y109_AO6),
.I1(CLBLM_L_X10Y108_SLICE_X13Y108_BO6),
.I2(CLBLM_R_X11Y108_SLICE_X14Y108_DO6),
.I3(CLBLM_R_X11Y108_SLICE_X14Y108_CO6),
.I4(CLBLM_L_X10Y108_SLICE_X12Y108_AO6),
.I5(CLBLM_L_X10Y108_SLICE_X12Y108_AO5),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_BO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00f000f000)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_AO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h781ee1e187e1e1e1)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_DLUT (
.I0(CLBLM_L_X10Y109_SLICE_X13Y109_AO6),
.I1(CLBLM_R_X11Y107_SLICE_X14Y107_AO5),
.I2(CLBLM_R_X11Y108_SLICE_X14Y108_AO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(RIOB33_X105Y107_IOB_X1Y107_I),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_DO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h96a5695a5a96a569)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_CLUT (
.I0(CLBLM_L_X10Y107_SLICE_X13Y107_AO6),
.I1(CLBLM_R_X11Y106_SLICE_X14Y106_BO6),
.I2(CLBLM_L_X10Y107_SLICE_X13Y107_BO6),
.I3(CLBLM_L_X10Y108_SLICE_X13Y108_AO5),
.I4(CLBLM_L_X10Y108_SLICE_X13Y108_AO6),
.I5(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_CO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8f08088fef0e0eef)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_BLUT (
.I0(CLBLM_R_X11Y106_SLICE_X14Y106_BO6),
.I1(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I2(CLBLM_L_X10Y107_SLICE_X13Y107_AO6),
.I3(CLBLM_L_X10Y107_SLICE_X13Y107_BO6),
.I4(CLBLM_L_X10Y108_SLICE_X13Y108_AO6),
.I5(CLBLM_L_X10Y108_SLICE_X13Y108_AO5),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_BO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000ff000000)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_AO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_DO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfed5ea54a84080)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_CLUT (
.I0(CLBLM_L_X10Y109_SLICE_X12Y109_AO6),
.I1(CLBLM_L_X8Y108_SLICE_X11Y108_DO6),
.I2(CLBLM_R_X11Y109_SLICE_X14Y109_DO6),
.I3(CLBLM_L_X10Y108_SLICE_X12Y108_CO6),
.I4(CLBLM_R_X7Y109_SLICE_X8Y109_AO5),
.I5(CLBLM_L_X10Y112_SLICE_X12Y112_AO6),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_CO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he81717e817e8e817)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_BLUT (
.I0(CLBLM_R_X7Y109_SLICE_X8Y109_AO5),
.I1(CLBLM_R_X11Y109_SLICE_X14Y109_DO6),
.I2(CLBLM_L_X8Y108_SLICE_X11Y108_DO6),
.I3(CLBLM_L_X10Y112_SLICE_X12Y112_AO6),
.I4(CLBLM_L_X10Y109_SLICE_X12Y109_AO6),
.I5(CLBLM_L_X10Y108_SLICE_X12Y108_CO6),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_BO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f0f00000)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_AO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h963c69c366cc9933)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_L_X10Y108_SLICE_X13Y108_BO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(CLBLM_R_X11Y108_SLICE_X14Y108_AO6),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_DO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8e0c4dcfeeccddff)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_L_X10Y108_SLICE_X13Y108_BO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(CLBLM_R_X11Y108_SLICE_X14Y108_AO6),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_CO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2fbcd043df4c20b3)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(CLBLM_R_X11Y106_SLICE_X14Y106_BO6),
.I4(CLBLM_L_X10Y107_SLICE_X13Y107_BO6),
.I5(RIOB33_X105Y107_IOB_X1Y107_I),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_BO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf4cdf4c936c936c)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(CLBLM_R_X11Y106_SLICE_X14Y106_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_AO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h366cc993c993366c)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_DLUT (
.I0(CLBLM_L_X10Y109_SLICE_X12Y109_AO6),
.I1(CLBLM_L_X10Y112_SLICE_X12Y112_AO5),
.I2(CLBLM_R_X11Y109_SLICE_X14Y109_BO6),
.I3(CLBLM_L_X10Y109_SLICE_X13Y109_DO6),
.I4(CLBLM_L_X10Y112_SLICE_X13Y112_AO5),
.I5(CLBLM_L_X10Y108_SLICE_X12Y108_BO6),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_DO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h04cd01374cdf137f)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_CLUT (
.I0(CLBLM_L_X10Y109_SLICE_X12Y109_AO6),
.I1(CLBLM_L_X10Y108_SLICE_X12Y108_BO6),
.I2(CLBLM_R_X11Y109_SLICE_X14Y109_BO6),
.I3(CLBLM_L_X10Y112_SLICE_X12Y112_AO5),
.I4(CLBLM_L_X10Y112_SLICE_X13Y112_AO5),
.I5(CLBLM_L_X10Y109_SLICE_X13Y109_DO6),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_CO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc93636c9936c6c93)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_BLUT (
.I0(CLBLM_L_X10Y110_SLICE_X12Y110_DO6),
.I1(CLBLM_L_X10Y110_SLICE_X12Y110_CO6),
.I2(CLBLM_L_X10Y109_SLICE_X12Y109_CO6),
.I3(CLBLM_L_X10Y111_SLICE_X12Y111_BO6),
.I4(CLBLM_L_X10Y110_SLICE_X12Y110_AO6),
.I5(CLBLM_L_X10Y110_SLICE_X12Y110_AO5),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_BO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00ff000000)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_AO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff6c6c006c006c00)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_DLUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(CLBLM_R_X11Y110_SLICE_X14Y110_DO6),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(CLBLM_L_X10Y111_SLICE_X13Y111_DO6),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_DO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996a55a96965a5a)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_CLUT (
.I0(CLBLM_R_X11Y109_SLICE_X14Y109_BO6),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(CLBLM_L_X10Y108_SLICE_X13Y108_DO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_CO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdeee48885aaa0000)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_BLUT (
.I0(CLBLM_L_X10Y108_SLICE_X13Y108_DO6),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(CLBLM_R_X11Y109_SLICE_X14Y109_BO6),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_BO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h22aa00004ec6a0a0)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_ALUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(RIOB33_X105Y111_IOB_X1Y111_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_AO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb230f3b22b033f2b)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_DLUT (
.I0(CLBLM_L_X10Y107_SLICE_X13Y107_CO6),
.I1(CLBLM_R_X7Y108_SLICE_X9Y108_AO5),
.I2(CLBLM_L_X10Y111_SLICE_X13Y111_BO5),
.I3(CLBLM_L_X10Y109_SLICE_X13Y109_CO6),
.I4(CLBLM_L_X10Y112_SLICE_X13Y112_AO5),
.I5(CLBLM_R_X11Y109_SLICE_X14Y109_CO6),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_DO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h73e6bf2a8c1940d5)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_CLUT (
.I0(CLBLM_L_X10Y107_SLICE_X13Y107_CO6),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y109_SLICE_X13Y109_CO6),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(CLBLM_R_X11Y109_SLICE_X14Y109_CO6),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_CO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc639639c39c69c63)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_BLUT (
.I0(CLBLM_L_X10Y112_SLICE_X13Y112_AO5),
.I1(CLBLM_L_X10Y111_SLICE_X13Y111_BO5),
.I2(CLBLM_L_X10Y109_SLICE_X13Y109_CO6),
.I3(CLBLM_R_X11Y109_SLICE_X14Y109_CO6),
.I4(CLBLM_L_X10Y107_SLICE_X13Y107_CO6),
.I5(CLBLM_R_X7Y108_SLICE_X9Y108_AO5),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_BO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha93f953f56c06ac0)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y110_SLICE_X13Y110_BO6),
.I2(CLBLM_L_X10Y111_SLICE_X13Y111_AO6),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(CLBLM_L_X10Y111_SLICE_X12Y111_CO6),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_AO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8ee8ee880aa0aa00)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_DLUT (
.I0(CLBLM_L_X12Y110_SLICE_X16Y110_CO6),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLM_R_X11Y110_SLICE_X15Y110_DO6),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_DO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999c33396663ccc)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_CLUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(CLBLM_R_X11Y110_SLICE_X14Y110_DO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(CLBLM_L_X10Y111_SLICE_X13Y111_DO6),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_CO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969a5a5cccc0000)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_BLUT (
.I0(CLBLM_L_X10Y107_SLICE_X13Y107_DO6),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(CLBLM_R_X11Y110_SLICE_X14Y110_AO6),
.I3(1'b1),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_BO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h93936c6cdfdf4c4c)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y109_SLICE_X13Y109_CO6),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(1'b1),
.I4(CLBLM_L_X10Y107_SLICE_X13Y107_CO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_AO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf9f6906090609060)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_DLUT (
.I0(CLBLM_L_X10Y110_SLICE_X13Y110_BO6),
.I1(CLBLM_L_X10Y111_SLICE_X13Y111_AO6),
.I2(CLBLM_L_X10Y109_SLICE_X12Y109_CO6),
.I3(CLBLM_L_X10Y112_SLICE_X12Y112_AO5),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_DO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaf0ea80e0800000)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_CLUT (
.I0(CLBLM_L_X10Y111_SLICE_X13Y111_AO6),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(CLBLM_L_X10Y110_SLICE_X13Y110_BO6),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLM_L_X10Y111_SLICE_X12Y111_BO6),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_CO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3963c963c69c3)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(CLBLM_L_X10Y109_SLICE_X12Y109_CO6),
.I2(CLBLM_L_X10Y111_SLICE_X13Y111_AO6),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(CLBLM_L_X10Y110_SLICE_X13Y110_BO6),
.I5(CLBLM_L_X10Y112_SLICE_X12Y112_AO5),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_BO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000aaaa0000)
  ) CLBLM_L_X10Y112_SLICE_X12Y112_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y112_SLICE_X12Y112_AO5),
.O6(CLBLM_L_X10Y112_SLICE_X12Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8f0eaf8eefaeffee)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_DLUT (
.I0(CLBLM_R_X11Y111_SLICE_X14Y111_BO6),
.I1(CLBLM_L_X10Y111_SLICE_X13Y111_BO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y111_SLICE_X13Y111_AO5),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_DO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9556a59665a65566)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_CLUT (
.I0(CLBLM_R_X11Y111_SLICE_X14Y111_BO6),
.I1(CLBLM_L_X10Y111_SLICE_X13Y111_BO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y111_SLICE_X13Y111_AO5),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_CO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8d72d72887787788)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(CLBLM_L_X10Y110_SLICE_X13Y110_BO6),
.I3(CLBLM_L_X10Y111_SLICE_X12Y111_BO6),
.I4(CLBLM_L_X10Y111_SLICE_X13Y111_AO6),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_BO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00cccc0000)
  ) CLBLM_L_X10Y112_SLICE_X13Y112_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y112_SLICE_X13Y112_AO5),
.O6(CLBLM_L_X10Y112_SLICE_X13Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_DO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h693cc36996c33c96)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_CLUT (
.I0(CLBLM_R_X11Y111_SLICE_X14Y111_BO6),
.I1(CLBLM_L_X10Y113_SLICE_X12Y113_AO6),
.I2(CLBLM_R_X11Y111_SLICE_X14Y111_AO5),
.I3(CLBLM_L_X10Y112_SLICE_X13Y112_AO6),
.I4(CLBLM_L_X10Y111_SLICE_X12Y111_DO6),
.I5(CLBLM_R_X11Y111_SLICE_X14Y111_CO6),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_CO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a5965a5a69a596)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_BLUT (
.I0(CLBLM_L_X10Y111_SLICE_X12Y111_DO6),
.I1(CLBLM_L_X10Y110_SLICE_X12Y110_AO6),
.I2(CLBLM_L_X10Y112_SLICE_X13Y112_AO6),
.I3(CLBLM_L_X10Y111_SLICE_X12Y111_BO6),
.I4(CLBLM_R_X11Y111_SLICE_X14Y111_BO6),
.I5(CLBLM_L_X10Y110_SLICE_X12Y110_CO6),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_BO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f00096669666)
  ) CLBLM_L_X10Y113_SLICE_X12Y113_ALUT (
.I0(CLBLM_R_X11Y111_SLICE_X14Y111_AO5),
.I1(CLBLM_R_X11Y111_SLICE_X14Y111_CO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y113_SLICE_X12Y113_AO5),
.O6(CLBLM_L_X10Y113_SLICE_X12Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_DO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_CO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_BO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y113_SLICE_X13Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y113_SLICE_X13Y113_AO5),
.O6(CLBLM_L_X10Y113_SLICE_X13Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y107_SLICE_X16Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y107_SLICE_X16Y107_DO5),
.O6(CLBLM_L_X12Y107_SLICE_X16Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y107_SLICE_X16Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y107_SLICE_X16Y107_CO5),
.O6(CLBLM_L_X12Y107_SLICE_X16Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y107_SLICE_X16Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y107_SLICE_X16Y107_BO5),
.O6(CLBLM_L_X12Y107_SLICE_X16Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h138a1b0a64a8e428)
  ) CLBLM_L_X12Y107_SLICE_X16Y107_ALUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(RIOB33_X105Y109_IOB_X1Y109_I),
.O5(CLBLM_L_X12Y107_SLICE_X16Y107_AO5),
.O6(CLBLM_L_X12Y107_SLICE_X16Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y107_SLICE_X17Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y107_SLICE_X17Y107_DO5),
.O6(CLBLM_L_X12Y107_SLICE_X17Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y107_SLICE_X17Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y107_SLICE_X17Y107_CO5),
.O6(CLBLM_L_X12Y107_SLICE_X17Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y107_SLICE_X17Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y107_SLICE_X17Y107_BO5),
.O6(CLBLM_L_X12Y107_SLICE_X17Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y107_SLICE_X17Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y107_SLICE_X17Y107_AO5),
.O6(CLBLM_L_X12Y107_SLICE_X17Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y108_SLICE_X16Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y108_SLICE_X16Y108_DO5),
.O6(CLBLM_L_X12Y108_SLICE_X16Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y108_SLICE_X16Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y108_SLICE_X16Y108_CO5),
.O6(CLBLM_L_X12Y108_SLICE_X16Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb61cda700aa0aa00)
  ) CLBLM_L_X12Y108_SLICE_X16Y108_BLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLM_L_X12Y108_SLICE_X16Y108_AO6),
.I5(RIOB33_X105Y111_IOB_X1Y111_I),
.O5(CLBLM_L_X12Y108_SLICE_X16Y108_BO5),
.O6(CLBLM_L_X12Y108_SLICE_X16Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha2a0a000a0000000)
  ) CLBLM_L_X12Y108_SLICE_X16Y108_ALUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(RIOB33_X105Y111_IOB_X1Y111_I),
.O5(CLBLM_L_X12Y108_SLICE_X16Y108_AO5),
.O6(CLBLM_L_X12Y108_SLICE_X16Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y108_SLICE_X17Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y108_SLICE_X17Y108_DO5),
.O6(CLBLM_L_X12Y108_SLICE_X17Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y108_SLICE_X17Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y108_SLICE_X17Y108_CO5),
.O6(CLBLM_L_X12Y108_SLICE_X17Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y108_SLICE_X17Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y108_SLICE_X17Y108_BO5),
.O6(CLBLM_L_X12Y108_SLICE_X17Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y108_SLICE_X17Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y108_SLICE_X17Y108_AO5),
.O6(CLBLM_L_X12Y108_SLICE_X17Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y109_SLICE_X16Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y109_SLICE_X16Y109_DO5),
.O6(CLBLM_L_X12Y109_SLICE_X16Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y109_SLICE_X16Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y109_SLICE_X16Y109_CO5),
.O6(CLBLM_L_X12Y109_SLICE_X16Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y109_SLICE_X16Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y109_SLICE_X16Y109_BO5),
.O6(CLBLM_L_X12Y109_SLICE_X16Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8e8c00080000000)
  ) CLBLM_L_X12Y109_SLICE_X16Y109_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLM_L_X12Y108_SLICE_X16Y108_AO6),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_L_X12Y109_SLICE_X16Y109_AO5),
.O6(CLBLM_L_X12Y109_SLICE_X16Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y109_SLICE_X17Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y109_SLICE_X17Y109_DO5),
.O6(CLBLM_L_X12Y109_SLICE_X17Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y109_SLICE_X17Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y109_SLICE_X17Y109_CO5),
.O6(CLBLM_L_X12Y109_SLICE_X17Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y109_SLICE_X17Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y109_SLICE_X17Y109_BO5),
.O6(CLBLM_L_X12Y109_SLICE_X17Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y109_SLICE_X17Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y109_SLICE_X17Y109_AO5),
.O6(CLBLM_L_X12Y109_SLICE_X17Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1780c8003f808000)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_DLUT (
.I0(CLBLM_L_X12Y108_SLICE_X16Y108_AO6),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(LIOB33_X0Y101_IOB_X0Y101_I),
.O5(CLBLM_L_X12Y110_SLICE_X16Y110_DO5),
.O6(CLBLM_L_X12Y110_SLICE_X16Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf4c4c4cec808080)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLM_L_X12Y110_SLICE_X17Y110_CO6),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(CLBLM_L_X12Y110_SLICE_X16Y110_BO6),
.O5(CLBLM_L_X12Y110_SLICE_X16Y110_CO5),
.O6(CLBLM_L_X12Y110_SLICE_X16Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h46806a006a802a00)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(CLBLM_L_X12Y109_SLICE_X16Y109_AO6),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_L_X12Y110_SLICE_X16Y110_BO5),
.O6(CLBLM_L_X12Y110_SLICE_X16Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996a55ac33c0ff0)
  ) CLBLM_L_X12Y110_SLICE_X16Y110_ALUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(CLBLM_L_X12Y110_SLICE_X17Y110_CO6),
.I3(CLBLM_L_X12Y110_SLICE_X16Y110_BO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLM_L_X12Y110_SLICE_X16Y110_AO5),
.O6(CLBLM_L_X12Y110_SLICE_X16Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd7289f604848c0c0)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_DLUT (
.I0(CLBLM_L_X12Y109_SLICE_X16Y109_AO6),
.I1(RIOB33_X105Y111_IOB_X1Y111_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(RIOB33_X105Y109_IOB_X1Y110_I),
.O5(CLBLM_L_X12Y110_SLICE_X17Y110_DO5),
.O6(CLBLM_L_X12Y110_SLICE_X17Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeecc880aa000000)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_CLUT (
.I0(CLBLM_R_X11Y110_SLICE_X15Y110_AO5),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_R_X11Y108_SLICE_X15Y108_BO6),
.I4(CLBLM_L_X12Y110_SLICE_X17Y110_DO6),
.I5(RIOB33_X105Y109_IOB_X1Y109_I),
.O5(CLBLM_L_X12Y110_SLICE_X17Y110_CO5),
.O6(CLBLM_L_X12Y110_SLICE_X17Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h995a96aa965a66aa)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_BLUT (
.I0(CLBLM_L_X12Y110_SLICE_X17Y110_DO6),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(CLBLM_R_X11Y108_SLICE_X15Y108_BO6),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(CLBLM_R_X11Y110_SLICE_X15Y110_AO5),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_L_X12Y110_SLICE_X17Y110_BO5),
.O6(CLBLM_L_X12Y110_SLICE_X17Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe80c000a0000000)
  ) CLBLM_L_X12Y110_SLICE_X17Y110_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(CLBLM_L_X12Y109_SLICE_X16Y109_AO6),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(RIOB33_X105Y111_IOB_X1Y111_I),
.O5(CLBLM_L_X12Y110_SLICE_X17Y110_AO5),
.O6(CLBLM_L_X12Y110_SLICE_X17Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y103_SLICE_X2Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y103_SLICE_X2Y103_DO5),
.O6(CLBLM_R_X3Y103_SLICE_X2Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y103_SLICE_X2Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y103_SLICE_X2Y103_CO5),
.O6(CLBLM_R_X3Y103_SLICE_X2Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y103_SLICE_X2Y103_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y103_SLICE_X2Y103_BO5),
.O6(CLBLM_R_X3Y103_SLICE_X2Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y103_SLICE_X2Y103_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y103_SLICE_X2Y103_AO5),
.O6(CLBLM_R_X3Y103_SLICE_X2Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y103_SLICE_X3Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y103_SLICE_X3Y103_DO5),
.O6(CLBLM_R_X3Y103_SLICE_X3Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y103_SLICE_X3Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y103_SLICE_X3Y103_CO5),
.O6(CLBLM_R_X3Y103_SLICE_X3Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y103_SLICE_X3Y103_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y103_SLICE_X3Y103_BO5),
.O6(CLBLM_R_X3Y103_SLICE_X3Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hacffa655cc5533ff)
  ) CLBLM_R_X3Y103_SLICE_X3Y103_ALUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_R_X3Y103_SLICE_X3Y103_AO5),
.O6(CLBLM_R_X3Y103_SLICE_X3Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y104_SLICE_X2Y104_DO5),
.O6(CLBLM_R_X3Y104_SLICE_X2Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5af05af0eecc8800)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLM_R_X5Y102_SLICE_X6Y102_AO6),
.I2(CLBLM_R_X3Y104_SLICE_X3Y104_BO6),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(CLBLM_R_X3Y104_SLICE_X2Y104_BO5),
.I5(1'b1),
.O5(CLBLM_R_X3Y104_SLICE_X2Y104_CO5),
.O6(CLBLM_R_X3Y104_SLICE_X2Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3635f5f30b0a0a0)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_BLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y104_SLICE_X2Y104_BO5),
.O6(CLBLM_R_X3Y104_SLICE_X2Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00f000f000)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y104_SLICE_X2Y104_AO5),
.O6(CLBLM_R_X3Y104_SLICE_X2Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h396c936c93399393)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_DLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(CLBLM_R_X5Y101_SLICE_X6Y101_BO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_R_X3Y104_SLICE_X3Y104_AO5),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLM_R_X3Y104_SLICE_X2Y104_CO5),
.O5(CLBLM_R_X3Y104_SLICE_X3Y104_DO5),
.O6(CLBLM_R_X3Y104_SLICE_X3Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h66696999a5a55555)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_CLUT (
.I0(CLBLM_R_X3Y103_SLICE_X3Y103_AO6),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_R_X3Y104_SLICE_X2Y104_BO5),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(CLBLM_R_X5Y102_SLICE_X6Y102_AO6),
.I5(LIOB33_X0Y101_IOB_X0Y101_I),
.O5(CLBLM_R_X3Y104_SLICE_X3Y104_CO5),
.O6(CLBLM_R_X3Y104_SLICE_X3Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbf8f95a5f5050fff)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_BLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X3Y104_SLICE_X3Y104_BO5),
.O6(CLBLM_R_X3Y104_SLICE_X3Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00a5a50f0f)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(1'b1),
.I2(CLBLM_R_X3Y103_SLICE_X3Y103_AO6),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y104_SLICE_X3Y104_AO5),
.O6(CLBLM_R_X3Y104_SLICE_X3Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4cdf80ecdfdfecec)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_DLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLL_L_X2Y105_SLICE_X0Y105_BO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(CLBLM_R_X3Y105_SLICE_X2Y105_BO6),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_R_X3Y105_SLICE_X2Y105_DO5),
.O6(CLBLM_R_X3Y105_SLICE_X2Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93936c936c936c)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLM_R_X3Y104_SLICE_X3Y104_CO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLL_L_X2Y105_SLICE_X1Y105_DO6),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X3Y105_SLICE_X2Y105_CO5),
.O6(CLBLM_R_X3Y105_SLICE_X2Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd21e965ab4783cf0)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_BLUT (
.I0(CLBLL_L_X2Y105_SLICE_X1Y105_AO5),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(CLBLM_R_X3Y104_SLICE_X3Y104_CO6),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLM_R_X3Y104_SLICE_X2Y104_CO6),
.O5(CLBLM_R_X3Y105_SLICE_X2Y105_BO5),
.O6(CLBLM_R_X3Y105_SLICE_X2Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc396963c3c6969c3)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_ALUT (
.I0(CLBLM_R_X3Y107_SLICE_X3Y107_BO5),
.I1(CLBLL_L_X4Y104_SLICE_X4Y104_BO6),
.I2(CLBLM_R_X3Y105_SLICE_X3Y105_AO6),
.I3(CLBLM_R_X3Y107_SLICE_X2Y107_BO6),
.I4(CLBLL_L_X2Y105_SLICE_X1Y105_CO6),
.I5(CLBLL_L_X2Y105_SLICE_X1Y105_DO6),
.O5(CLBLM_R_X3Y105_SLICE_X2Y105_AO5),
.O6(CLBLM_R_X3Y105_SLICE_X2Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996a55ac33c0ff0)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(CLBLM_R_X3Y104_SLICE_X3Y104_DO6),
.I3(CLBLM_R_X3Y105_SLICE_X3Y105_CO6),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLM_R_X3Y105_SLICE_X3Y105_DO5),
.O6(CLBLM_R_X3Y105_SLICE_X3Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff87870087008700)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_CLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(CLBLM_R_X3Y104_SLICE_X3Y104_CO6),
.I3(CLBLL_L_X2Y105_SLICE_X1Y105_DO6),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLM_R_X3Y105_SLICE_X3Y105_CO5),
.O6(CLBLM_R_X3Y105_SLICE_X3Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h693cc36996c33c96)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_BLUT (
.I0(CLBLL_L_X2Y105_SLICE_X1Y105_DO6),
.I1(CLBLL_L_X4Y104_SLICE_X4Y104_CO6),
.I2(CLBLM_R_X5Y102_SLICE_X6Y102_BO6),
.I3(CLBLL_L_X4Y104_SLICE_X4Y104_BO6),
.I4(CLBLM_R_X3Y105_SLICE_X3Y105_AO6),
.I5(CLBLM_R_X3Y105_SLICE_X3Y105_AO5),
.O5(CLBLM_R_X3Y105_SLICE_X3Y105_BO5),
.O6(CLBLM_R_X3Y105_SLICE_X3Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000cccc0000)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(1'b1),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y105_SLICE_X3Y105_AO5),
.O6(CLBLM_R_X3Y105_SLICE_X3Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4504df5d8a08efae)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_DLUT (
.I0(CLBLL_L_X4Y105_SLICE_X5Y105_AO6),
.I1(CLBLM_R_X3Y105_SLICE_X2Y105_CO6),
.I2(CLBLL_L_X2Y106_SLICE_X1Y106_AO5),
.I3(CLBLL_L_X2Y105_SLICE_X0Y105_BO6),
.I4(CLBLL_L_X2Y106_SLICE_X1Y106_BO5),
.I5(CLBLM_R_X3Y105_SLICE_X3Y105_BO6),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_DO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd42b03fc2bd403fc)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(CLBLM_R_X3Y105_SLICE_X2Y105_CO6),
.I2(CLBLL_L_X2Y105_SLICE_X0Y105_BO6),
.I3(CLBLM_R_X3Y105_SLICE_X3Y105_BO6),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_CO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h963c69c366cc9933)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(CLBLL_L_X2Y105_SLICE_X0Y105_BO6),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(CLBLM_R_X3Y105_SLICE_X2Y105_BO6),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_BO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd5b97f132a4680ec)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLL_L_X2Y106_SLICE_X1Y106_CO6),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(CLBLM_R_X3Y106_SLICE_X2Y106_BO6),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLM_R_X3Y106_SLICE_X2Y106_CO6),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_AO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf4c5f007f13ff5f)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLM_R_X3Y106_SLICE_X3Y106_CO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_R_X3Y106_SLICE_X3Y106_BO6),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_DO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf4c7f137f137f13)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(CLBLM_R_X3Y106_SLICE_X2Y106_CO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(CLBLL_L_X2Y106_SLICE_X1Y106_DO6),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_CO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h87781e1ee11e1e1e)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_BLUT (
.I0(CLBLM_R_X3Y105_SLICE_X2Y105_DO6),
.I1(CLBLM_R_X3Y105_SLICE_X3Y105_DO6),
.I2(CLBLL_L_X4Y105_SLICE_X4Y105_AO6),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_BO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h936c5fa06c93a05f)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(CLBLM_R_X3Y106_SLICE_X3Y106_BO6),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(CLBLM_R_X3Y106_SLICE_X3Y106_CO6),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_AO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996669999666996)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_DLUT (
.I0(CLBLL_L_X2Y105_SLICE_X1Y105_BO6),
.I1(CLBLM_R_X3Y107_SLICE_X3Y107_AO5),
.I2(CLBLL_L_X2Y107_SLICE_X1Y107_AO5),
.I3(CLBLM_R_X3Y109_SLICE_X3Y109_AO5),
.I4(CLBLM_R_X3Y108_SLICE_X2Y108_AO5),
.I5(CLBLL_L_X2Y106_SLICE_X0Y106_AO6),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_DO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h96c33c96693cc369)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_CLUT (
.I0(CLBLM_R_X3Y108_SLICE_X2Y108_CO6),
.I1(CLBLL_L_X2Y105_SLICE_X1Y105_CO6),
.I2(CLBLM_R_X3Y107_SLICE_X3Y107_BO5),
.I3(CLBLM_R_X3Y107_SLICE_X3Y107_BO6),
.I4(CLBLM_R_X3Y107_SLICE_X2Y107_DO6),
.I5(CLBLM_R_X3Y107_SLICE_X2Y107_BO6),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_CO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2bafb2fa0a2ba0b2)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_BLUT (
.I0(CLBLM_R_X3Y107_SLICE_X3Y107_AO5),
.I1(CLBLL_L_X2Y107_SLICE_X1Y107_AO5),
.I2(CLBLM_R_X3Y109_SLICE_X3Y109_AO5),
.I3(CLBLL_L_X2Y106_SLICE_X0Y106_AO6),
.I4(CLBLL_L_X2Y105_SLICE_X1Y105_BO6),
.I5(CLBLM_R_X3Y108_SLICE_X2Y108_AO5),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_BO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h693cccccc3699999)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_ALUT (
.I0(CLBLL_L_X2Y107_SLICE_X1Y107_AO5),
.I1(CLBLL_L_X2Y105_SLICE_X1Y105_BO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(CLBLL_L_X2Y106_SLICE_X0Y106_AO6),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_AO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h966969695aa5a5a5)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_DLUT (
.I0(CLBLL_L_X4Y105_SLICE_X4Y105_AO6),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(CLBLM_R_X3Y106_SLICE_X2Y106_DO6),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_DO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he94fb91fc9ef391f)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_CO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000cccc0000)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(1'b1),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_BO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000cc00cc00)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_AO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbf2a7f157f157f15)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_DLUT (
.I0(CLBLM_R_X3Y107_SLICE_X2Y107_AO6),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLM_R_X3Y108_SLICE_X2Y108_CO6),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_DO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc431fdf74010dc73)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_CLUT (
.I0(CLBLM_R_X3Y108_SLICE_X2Y108_AO6),
.I1(CLBLM_R_X3Y107_SLICE_X3Y107_CO6),
.I2(CLBLL_L_X2Y108_SLICE_X0Y108_AO5),
.I3(CLBLM_R_X3Y108_SLICE_X2Y108_AO5),
.I4(CLBLM_R_X3Y107_SLICE_X3Y107_AO6),
.I5(CLBLL_L_X2Y107_SLICE_X1Y107_AO6),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_CO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h953f6ac06ac0953f)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(CLBLM_R_X3Y107_SLICE_X2Y107_AO6),
.I5(CLBLM_R_X3Y108_SLICE_X2Y108_CO6),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_BO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000cccc0000)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_AO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h40c0c4dd0040c0d5)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_DLUT (
.I0(CLBLL_L_X4Y108_SLICE_X4Y108_AO6),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(CLBLM_R_X3Y106_SLICE_X3Y106_DO6),
.I4(CLBLL_L_X4Y108_SLICE_X4Y108_CO6),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_DO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c36c9c993c9c9c9)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_CLUT (
.I0(CLBLL_L_X4Y108_SLICE_X4Y108_AO6),
.I1(CLBLL_L_X4Y108_SLICE_X4Y108_BO6),
.I2(CLBLM_R_X3Y106_SLICE_X3Y106_DO6),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_CO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h050f577f577f5fff)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_BLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(CLBLL_L_X4Y107_SLICE_X4Y107_DO6),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(CLBLM_R_X3Y108_SLICE_X3Y108_AO6),
.I5(CLBLM_R_X3Y106_SLICE_X3Y106_AO6),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_BO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8f08f880f880f880)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_ALUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(CLBLM_R_X3Y106_SLICE_X2Y106_AO6),
.I3(CLBLL_L_X2Y108_SLICE_X1Y108_CO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_AO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_DO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_CO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66cc693369339933)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(CLBLL_L_X4Y106_SLICE_X4Y106_BO6),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(CLBLM_R_X3Y108_SLICE_X3Y108_AO6),
.I5(CLBLM_R_X3Y106_SLICE_X3Y106_AO6),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_BO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00aa00aa00)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_ALUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(1'b1),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_AO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h21b71177b7b77777)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_DLUT (
.I0(CLBLL_L_X4Y108_SLICE_X5Y108_AO6),
.I1(CLBLM_R_X3Y108_SLICE_X3Y108_DO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_DO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9669696966999999)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_CLUT (
.I0(CLBLL_L_X4Y108_SLICE_X5Y108_AO6),
.I1(CLBLM_R_X3Y108_SLICE_X3Y108_DO6),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_CO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he888e888f000f000)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_BLUT (
.I0(CLBLL_L_X4Y109_SLICE_X4Y109_BO5),
.I1(CLBLM_R_X5Y109_SLICE_X6Y109_CO6),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_BO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h99339933f000f000)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_ALUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(CLBLM_R_X5Y109_SLICE_X6Y109_BO6),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_AO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9f603fc0c53a956a)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_DLUT (
.I0(CLBLM_R_X3Y110_SLICE_X2Y110_AO6),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(CLBLM_R_X3Y110_SLICE_X2Y110_CO6),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(CLBLM_R_X3Y111_SLICE_X2Y111_AO6),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_DO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a5aa9699aaa5999)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_CLUT (
.I0(CLBLL_L_X4Y109_SLICE_X5Y109_DO6),
.I1(CLBLL_L_X4Y109_SLICE_X4Y109_BO6),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(CLBLM_R_X3Y109_SLICE_X3Y109_DO6),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_CO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c088888888)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_BO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha55a5a5aff000000)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_ALUT (
.I0(CLBLM_R_X3Y109_SLICE_X3Y109_DO6),
.I1(1'b1),
.I2(CLBLL_L_X4Y109_SLICE_X4Y109_BO6),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_AO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb332fb32ffb2fffa)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_DLUT (
.I0(CLBLL_L_X4Y109_SLICE_X4Y109_BO6),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(CLBLM_R_X3Y109_SLICE_X3Y109_DO6),
.I3(CLBLL_L_X4Y109_SLICE_X4Y109_DO6),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(LIOB33_X0Y113_IOB_X0Y113_I),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_DO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3595ca6a90c06f3f)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_CLUT (
.I0(CLBLM_R_X3Y109_SLICE_X3Y109_AO6),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(CLBLL_L_X4Y110_SLICE_X5Y110_AO6),
.I5(CLBLM_R_X3Y109_SLICE_X3Y109_BO6),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_CO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4fbfda2ab04025d5)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_BLUT (
.I0(CLBLM_R_X3Y109_SLICE_X3Y109_DO6),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(CLBLL_L_X4Y109_SLICE_X4Y109_BO6),
.I5(CLBLL_L_X4Y109_SLICE_X4Y109_DO6),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_BO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00003c3cf0f0)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(CLBLL_L_X4Y110_SLICE_X5Y110_AO6),
.I3(1'b1),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_AO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0082c3eb82c3ebff)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_DLUT (
.I0(CLBLM_R_X3Y109_SLICE_X3Y109_CO6),
.I1(CLBLM_R_X3Y110_SLICE_X2Y110_AO5),
.I2(CLBLL_L_X4Y109_SLICE_X4Y109_CO6),
.I3(CLBLM_R_X3Y109_SLICE_X2Y109_AO5),
.I4(CLBLM_R_X3Y110_SLICE_X2Y110_BO5),
.I5(CLBLM_R_X3Y111_SLICE_X2Y111_BO6),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_DO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h693c0ff0c3690f0f)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_CLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(CLBLL_L_X4Y109_SLICE_X4Y109_CO6),
.I3(CLBLM_R_X3Y109_SLICE_X3Y109_CO6),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(CLBLM_R_X3Y111_SLICE_X2Y111_BO6),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_CO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6cff006c006c006c)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_BLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(CLBLM_R_X3Y108_SLICE_X3Y108_CO6),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(CLBLM_R_X3Y108_SLICE_X3Y108_BO6),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_BO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fff005f5fa0a05f)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_ALUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(1'b1),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(CLBLM_R_X3Y111_SLICE_X2Y111_BO6),
.I4(CLBLM_R_X3Y109_SLICE_X3Y109_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_AO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2f0bbf2f0b022f0b)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_DLUT (
.I0(CLBLM_R_X3Y110_SLICE_X3Y110_AO5),
.I1(CLBLM_R_X3Y112_SLICE_X3Y112_BO6),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_DO6),
.I3(CLBLM_R_X3Y111_SLICE_X3Y111_CO6),
.I4(CLBLL_L_X4Y110_SLICE_X4Y110_DO6),
.I5(CLBLM_R_X3Y111_SLICE_X3Y111_BO6),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_DO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999666996669996)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_CLUT (
.I0(CLBLM_R_X3Y111_SLICE_X3Y111_AO6),
.I1(CLBLM_R_X3Y110_SLICE_X3Y110_DO6),
.I2(CLBLM_R_X3Y111_SLICE_X2Y111_DO6),
.I3(CLBLM_R_X3Y110_SLICE_X3Y110_BO6),
.I4(CLBLM_R_X3Y110_SLICE_X2Y110_BO6),
.I5(CLBLL_L_X4Y110_SLICE_X4Y110_BO6),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_CO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc60af5c6c905fac9)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_BLUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_AO6),
.I1(CLBLM_R_X3Y110_SLICE_X3Y110_DO6),
.I2(CLBLM_R_X5Y110_SLICE_X6Y110_CO6),
.I3(CLBLL_L_X4Y110_SLICE_X4Y110_BO6),
.I4(CLBLM_R_X3Y111_SLICE_X3Y111_AO6),
.I5(CLBLM_R_X3Y111_SLICE_X3Y111_AO5),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_BO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000aa00aa00)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_AO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_DO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_CO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_BO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_AO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00b3002000fb0032)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_DLUT (
.I0(CLBLM_R_X3Y111_SLICE_X3Y111_CO6),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_DO6),
.I2(CLBLM_R_X3Y111_SLICE_X3Y111_BO6),
.I3(CLBLL_L_X4Y113_SLICE_X4Y113_CO6),
.I4(CLBLL_L_X4Y111_SLICE_X4Y111_AO6),
.I5(CLBLL_L_X4Y111_SLICE_X4Y111_BO6),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_DO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h565a59556aaa9a5a)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_CLUT (
.I0(CLBLM_R_X3Y112_SLICE_X3Y112_AO6),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(CLBLM_R_X3Y111_SLICE_X3Y111_BO6),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(CLBLM_R_X3Y110_SLICE_X3Y110_CO6),
.I5(CLBLM_R_X3Y111_SLICE_X3Y111_CO6),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_CO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc0069a5965a)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_BLUT (
.I0(CLBLM_R_X3Y110_SLICE_X3Y110_CO6),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(CLBLM_R_X3Y111_SLICE_X3Y111_BO6),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(CLBLM_R_X3Y111_SLICE_X3Y111_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_BO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc33c0ff0cccc0000)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(CLBLL_L_X4Y111_SLICE_X4Y111_AO6),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_BO6),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_AO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y101_SLICE_X6Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y101_SLICE_X6Y101_DO5),
.O6(CLBLM_R_X5Y101_SLICE_X6Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h18e8e71778888777)
  ) CLBLM_R_X5Y101_SLICE_X6Y101_CLUT (
.I0(CLBLM_R_X5Y101_SLICE_X6Y101_AO6),
.I1(CLBLM_R_X5Y101_SLICE_X7Y101_AO6),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLM_R_X5Y102_SLICE_X7Y102_CO6),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X5Y101_SLICE_X6Y101_CO5),
.O6(CLBLM_R_X5Y101_SLICE_X6Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4db2fafab24d0505)
  ) CLBLM_R_X5Y101_SLICE_X6Y101_BLUT (
.I0(CLBLM_R_X5Y102_SLICE_X6Y102_AO5),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_R_X5Y102_SLICE_X7Y102_AO6),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(CLBLM_R_X5Y102_SLICE_X6Y102_CO6),
.O5(CLBLM_R_X5Y101_SLICE_X6Y101_BO5),
.O6(CLBLM_R_X5Y101_SLICE_X6Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4d054d05cc00cc00)
  ) CLBLM_R_X5Y101_SLICE_X6Y101_ALUT (
.I0(CLBLM_R_X5Y102_SLICE_X6Y102_AO5),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_R_X5Y102_SLICE_X7Y102_AO6),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y101_SLICE_X6Y101_AO5),
.O6(CLBLM_R_X5Y101_SLICE_X6Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y101_SLICE_X7Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y101_SLICE_X7Y101_DO5),
.O6(CLBLM_R_X5Y101_SLICE_X7Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y101_SLICE_X7Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y101_SLICE_X7Y101_CO5),
.O6(CLBLM_R_X5Y101_SLICE_X7Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y101_SLICE_X7Y101_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y101_SLICE_X7Y101_BO5),
.O6(CLBLM_R_X5Y101_SLICE_X7Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6666aaaafcc0f000)
  ) CLBLM_R_X5Y101_SLICE_X7Y101_ALUT (
.I0(CLBLM_R_X5Y102_SLICE_X6Y102_CO6),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(CLBLM_R_X7Y102_SLICE_X8Y102_BO5),
.I3(CLBLM_R_X5Y102_SLICE_X7Y102_AO5),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y101_SLICE_X7Y101_AO5),
.O6(CLBLM_R_X5Y101_SLICE_X7Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha220fbba5110f775)
  ) CLBLM_R_X5Y102_SLICE_X6Y102_DLUT (
.I0(CLBLM_R_X5Y102_SLICE_X6Y102_CO6),
.I1(CLBLM_R_X5Y101_SLICE_X6Y101_AO5),
.I2(CLBLM_R_X5Y102_SLICE_X7Y102_AO6),
.I3(CLBLM_R_X5Y102_SLICE_X6Y102_AO5),
.I4(CLBLM_R_X3Y104_SLICE_X3Y104_AO6),
.I5(CLBLL_L_X4Y104_SLICE_X4Y104_AO5),
.O5(CLBLM_R_X5Y102_SLICE_X6Y102_DO5),
.O6(CLBLM_R_X5Y102_SLICE_X6Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hed9921ffa599e1ff)
  ) CLBLM_R_X5Y102_SLICE_X6Y102_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_R_X5Y102_SLICE_X6Y102_CO5),
.O6(CLBLM_R_X5Y102_SLICE_X6Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h59a6a6599a65659a)
  ) CLBLM_R_X5Y102_SLICE_X6Y102_BLUT (
.I0(CLBLM_R_X3Y104_SLICE_X3Y104_AO6),
.I1(CLBLM_R_X5Y101_SLICE_X6Y101_AO5),
.I2(CLBLM_R_X5Y102_SLICE_X7Y102_AO6),
.I3(CLBLL_L_X4Y104_SLICE_X4Y104_AO5),
.I4(CLBLM_R_X5Y102_SLICE_X6Y102_CO6),
.I5(CLBLM_R_X5Y102_SLICE_X6Y102_AO5),
.O5(CLBLM_R_X5Y102_SLICE_X6Y102_BO5),
.O6(CLBLM_R_X5Y102_SLICE_X6Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h993f593fd1ff51ff)
  ) CLBLM_R_X5Y102_SLICE_X6Y102_ALUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y102_SLICE_X6Y102_AO5),
.O6(CLBLM_R_X5Y102_SLICE_X6Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfae8f5d4e8a0d450)
  ) CLBLM_R_X5Y102_SLICE_X7Y102_DLUT (
.I0(CLBLM_R_X7Y102_SLICE_X9Y102_AO6),
.I1(CLBLM_R_X7Y102_SLICE_X8Y102_BO5),
.I2(CLBLM_R_X7Y102_SLICE_X8Y102_CO5),
.I3(CLBLM_R_X5Y102_SLICE_X7Y102_AO5),
.I4(CLBLM_R_X7Y102_SLICE_X8Y102_DO6),
.I5(CLBLL_L_X4Y104_SLICE_X4Y104_AO5),
.O5(CLBLM_R_X5Y102_SLICE_X7Y102_DO5),
.O6(CLBLM_R_X5Y102_SLICE_X7Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc993366c3ccc3ccc)
  ) CLBLM_R_X5Y102_SLICE_X7Y102_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(CLBLM_R_X7Y102_SLICE_X8Y102_DO6),
.I2(CLBLM_R_X7Y102_SLICE_X8Y102_BO5),
.I3(CLBLM_R_X5Y102_SLICE_X7Y102_AO5),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(LIOB33_X0Y101_IOB_X0Y101_I),
.O5(CLBLM_R_X5Y102_SLICE_X7Y102_CO5),
.O6(CLBLM_R_X5Y102_SLICE_X7Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h17e8e817e81717e8)
  ) CLBLM_R_X5Y102_SLICE_X7Y102_BLUT (
.I0(CLBLM_R_X7Y102_SLICE_X8Y102_BO5),
.I1(CLBLL_L_X4Y104_SLICE_X4Y104_AO5),
.I2(CLBLM_R_X5Y102_SLICE_X7Y102_AO5),
.I3(CLBLM_R_X7Y102_SLICE_X8Y102_DO6),
.I4(CLBLM_R_X7Y102_SLICE_X9Y102_AO6),
.I5(CLBLM_R_X7Y102_SLICE_X8Y102_CO5),
.O5(CLBLM_R_X5Y102_SLICE_X7Y102_BO5),
.O6(CLBLM_R_X5Y102_SLICE_X7Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c66aa004cee0000)
  ) CLBLM_R_X5Y102_SLICE_X7Y102_ALUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y102_SLICE_X7Y102_AO5),
.O6(CLBLM_R_X5Y102_SLICE_X7Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fb31320ffff5fa0)
  ) CLBLM_R_X5Y103_SLICE_X6Y103_DLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLM_R_X5Y102_SLICE_X7Y102_CO6),
.I4(CLBLM_R_X5Y102_SLICE_X6Y102_DO6),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X5Y103_SLICE_X6Y103_DO5),
.O6(CLBLM_R_X5Y103_SLICE_X6Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h936c6c935fa0a05f)
  ) CLBLM_R_X5Y103_SLICE_X6Y103_CLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLM_R_X5Y102_SLICE_X7Y102_CO6),
.I4(CLBLM_R_X5Y102_SLICE_X6Y102_DO6),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X5Y103_SLICE_X6Y103_CO5),
.O6(CLBLM_R_X5Y103_SLICE_X6Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h78871ee18778e11e)
  ) CLBLM_R_X5Y103_SLICE_X6Y103_BLUT (
.I0(CLBLM_R_X5Y102_SLICE_X6Y102_DO6),
.I1(CLBLM_R_X5Y102_SLICE_X7Y102_BO6),
.I2(CLBLM_R_X7Y102_SLICE_X9Y102_BO6),
.I3(CLBLM_R_X5Y102_SLICE_X7Y102_DO6),
.I4(CLBLM_R_X5Y103_SLICE_X6Y103_AO6),
.I5(CLBLM_R_X5Y103_SLICE_X6Y103_AO5),
.O5(CLBLM_R_X5Y103_SLICE_X6Y103_BO5),
.O6(CLBLM_R_X5Y103_SLICE_X6Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000f0f00000)
  ) CLBLM_R_X5Y103_SLICE_X6Y103_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(1'b1),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y103_SLICE_X6Y103_AO5),
.O6(CLBLM_R_X5Y103_SLICE_X6Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y103_SLICE_X7Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y103_SLICE_X7Y103_DO5),
.O6(CLBLM_R_X5Y103_SLICE_X7Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y103_SLICE_X7Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y103_SLICE_X7Y103_CO5),
.O6(CLBLM_R_X5Y103_SLICE_X7Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y103_SLICE_X7Y103_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y103_SLICE_X7Y103_BO5),
.O6(CLBLM_R_X5Y103_SLICE_X7Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h9f60c03f3fc09f60)
  ) CLBLM_R_X5Y103_SLICE_X7Y103_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(CLBLM_R_X7Y102_SLICE_X9Y102_DO6),
.I4(CLBLM_R_X7Y102_SLICE_X8Y102_AO6),
.I5(CLBLM_R_X5Y101_SLICE_X7Y101_AO5),
.O5(CLBLM_R_X5Y103_SLICE_X7Y103_AO5),
.O6(CLBLM_R_X5Y103_SLICE_X7Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hce083b02ef8cbf23)
  ) CLBLM_R_X5Y104_SLICE_X6Y104_DLUT (
.I0(CLBLM_R_X5Y105_SLICE_X6Y105_AO6),
.I1(CLBLM_R_X7Y103_SLICE_X8Y103_AO6),
.I2(CLBLM_R_X5Y103_SLICE_X6Y103_DO6),
.I3(CLBLM_R_X7Y105_SLICE_X8Y105_AO6),
.I4(CLBLM_R_X5Y105_SLICE_X6Y105_AO5),
.I5(CLBLM_R_X5Y104_SLICE_X6Y104_BO6),
.O5(CLBLM_R_X5Y104_SLICE_X6Y104_DO5),
.O6(CLBLM_R_X5Y104_SLICE_X6Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9699333366963c3c)
  ) CLBLM_R_X5Y104_SLICE_X6Y104_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(CLBLM_R_X7Y103_SLICE_X8Y103_AO6),
.I2(CLBLM_R_X5Y103_SLICE_X6Y103_DO6),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(CLBLM_R_X5Y104_SLICE_X6Y104_BO6),
.O5(CLBLM_R_X5Y104_SLICE_X6Y104_CO5),
.O6(CLBLM_R_X5Y104_SLICE_X6Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7888877787777888)
  ) CLBLM_R_X5Y104_SLICE_X6Y104_BLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLM_R_X7Y102_SLICE_X9Y102_DO6),
.I5(CLBLM_R_X5Y102_SLICE_X7Y102_DO6),
.O5(CLBLM_R_X5Y104_SLICE_X6Y104_BO5),
.O6(CLBLM_R_X5Y104_SLICE_X6Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h9c3963c663c69c39)
  ) CLBLM_R_X5Y104_SLICE_X6Y104_ALUT (
.I0(CLBLM_R_X5Y103_SLICE_X6Y103_DO6),
.I1(CLBLM_R_X7Y103_SLICE_X8Y103_AO6),
.I2(CLBLM_R_X5Y105_SLICE_X6Y105_AO6),
.I3(CLBLM_R_X5Y104_SLICE_X6Y104_BO6),
.I4(CLBLM_R_X5Y105_SLICE_X6Y105_AO5),
.I5(CLBLM_R_X7Y105_SLICE_X8Y105_AO6),
.O5(CLBLM_R_X5Y104_SLICE_X6Y104_AO5),
.O6(CLBLM_R_X5Y104_SLICE_X6Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y104_SLICE_X7Y104_DO5),
.O6(CLBLM_R_X5Y104_SLICE_X7Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y104_SLICE_X7Y104_CO5),
.O6(CLBLM_R_X5Y104_SLICE_X7Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y104_SLICE_X7Y104_BO5),
.O6(CLBLM_R_X5Y104_SLICE_X7Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h965a69a566aa9955)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_ALUT (
.I0(CLBLM_R_X5Y103_SLICE_X6Y103_DO6),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(CLBLM_R_X5Y103_SLICE_X7Y103_AO6),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_R_X5Y104_SLICE_X7Y104_AO5),
.O6(CLBLM_R_X5Y104_SLICE_X7Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb2e8e8e822888888)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_DLUT (
.I0(CLBLL_L_X4Y104_SLICE_X5Y104_BO6),
.I1(CLBLM_R_X5Y101_SLICE_X6Y101_CO6),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_DO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3696c66693c36333)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_CLUT (
.I0(CLBLM_R_X5Y104_SLICE_X7Y104_AO6),
.I1(CLBLM_R_X5Y104_SLICE_X6Y104_CO6),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_R_X5Y105_SLICE_X6Y105_DO6),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_CO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9669969669699669)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_BLUT (
.I0(CLBLM_R_X5Y102_SLICE_X6Y102_DO6),
.I1(CLBLM_R_X5Y102_SLICE_X7Y102_BO6),
.I2(CLBLM_R_X5Y103_SLICE_X6Y103_AO6),
.I3(CLBLL_L_X4Y104_SLICE_X4Y104_CO6),
.I4(CLBLM_R_X5Y102_SLICE_X6Y102_BO6),
.I5(CLBLM_R_X3Y105_SLICE_X3Y105_AO5),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_BO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00f000f000)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(1'b1),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_AO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_DO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_CO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_BO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_AO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8ff8ff8808808800)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_DLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_R_X5Y104_SLICE_X6Y104_CO6),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLL_L_X4Y104_SLICE_X5Y104_DO6),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_DO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb44b4bb42dd2d22d)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_CLUT (
.I0(CLBLM_R_X5Y106_SLICE_X6Y106_AO6),
.I1(CLBLM_R_X5Y104_SLICE_X6Y104_AO6),
.I2(CLBLM_R_X5Y104_SLICE_X6Y104_DO6),
.I3(CLBLM_R_X5Y106_SLICE_X6Y106_AO5),
.I4(CLBLM_R_X7Y105_SLICE_X8Y105_BO6),
.I5(CLBLL_L_X4Y104_SLICE_X5Y104_DO6),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_CO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h936c5fa06c93a05f)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(CLBLM_R_X5Y104_SLICE_X6Y104_CO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLL_L_X4Y104_SLICE_X5Y104_DO6),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_BO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0aaaa0000)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(1'b1),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(1'b1),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_AO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_DO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_CO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_BO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_AO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33c3cc36996)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_DLUT (
.I0(CLBLL_L_X4Y107_SLICE_X5Y107_BO6),
.I1(CLBLM_R_X5Y106_SLICE_X6Y106_CO6),
.I2(CLBLM_R_X7Y107_SLICE_X8Y107_AO6),
.I3(CLBLM_R_X5Y107_SLICE_X6Y107_AO5),
.I4(CLBLM_R_X5Y107_SLICE_X6Y107_AO6),
.I5(CLBLM_R_X5Y106_SLICE_X6Y106_BO6),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_DO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he8b2c030fcf3e8b2)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_CLUT (
.I0(CLBLL_L_X4Y107_SLICE_X5Y107_BO6),
.I1(CLBLM_R_X5Y106_SLICE_X6Y106_CO6),
.I2(CLBLM_R_X7Y107_SLICE_X8Y107_AO6),
.I3(CLBLM_R_X5Y107_SLICE_X6Y107_AO5),
.I4(CLBLM_R_X5Y107_SLICE_X6Y107_AO6),
.I5(CLBLM_R_X5Y106_SLICE_X6Y106_BO6),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_CO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb2cf4dcf4d30b230)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(CLBLM_R_X5Y106_SLICE_X6Y106_BO6),
.I2(CLBLL_L_X4Y107_SLICE_X5Y107_BO6),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLM_R_X5Y106_SLICE_X6Y106_CO6),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_BO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00f000f000)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(1'b1),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_AO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_DO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_CO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_BO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_AO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffa8ffffffffff)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(CLBLM_R_X7Y109_SLICE_X8Y109_DO6),
.I4(CLBLL_L_X2Y107_SLICE_X1Y107_DO6),
.I5(CLBLM_R_X3Y106_SLICE_X2Y106_CO6),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_DO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_CLUT (
.I0(CLBLM_R_X7Y107_SLICE_X9Y107_BO6),
.I1(CLBLM_R_X7Y108_SLICE_X9Y108_CO6),
.I2(CLBLM_R_X7Y108_SLICE_X8Y108_AO6),
.I3(CLBLM_R_X5Y107_SLICE_X6Y107_CO6),
.I4(CLBLM_R_X5Y108_SLICE_X6Y108_DO6),
.I5(CLBLM_L_X8Y107_SLICE_X10Y107_BO6),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_CO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9669699669966996)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_BLUT (
.I0(CLBLM_R_X7Y108_SLICE_X8Y108_CO6),
.I1(CLBLM_R_X7Y107_SLICE_X9Y107_BO6),
.I2(CLBLM_R_X7Y108_SLICE_X9Y108_AO6),
.I3(CLBLM_L_X8Y107_SLICE_X10Y107_BO6),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_BO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2bb20330b22b3003)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_ALUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(CLBLM_R_X7Y108_SLICE_X8Y108_CO6),
.I2(CLBLM_R_X7Y108_SLICE_X9Y108_AO6),
.I3(CLBLM_R_X7Y107_SLICE_X9Y107_BO6),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLM_L_X8Y107_SLICE_X10Y107_BO6),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_AO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_DO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_CO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_BO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_AO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996696996966996)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_DLUT (
.I0(CLBLM_R_X7Y108_SLICE_X8Y108_CO6),
.I1(CLBLM_R_X5Y109_SLICE_X7Y109_AO6),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_CO6),
.I3(CLBLM_R_X5Y107_SLICE_X6Y107_CO6),
.I4(CLBLM_R_X7Y108_SLICE_X8Y108_AO6),
.I5(CLBLM_L_X8Y111_SLICE_X11Y111_AO6),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_DO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996a55ac33c0ff0)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(CLBLL_L_X4Y109_SLICE_X5Y109_BO6),
.I3(CLBLM_R_X7Y107_SLICE_X8Y107_CO6),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_CO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9996966666696999)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_BLUT (
.I0(CLBLM_R_X7Y109_SLICE_X8Y109_BO6),
.I1(CLBLM_R_X7Y108_SLICE_X8Y108_BO6),
.I2(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.I3(CLBLM_R_X5Y108_SLICE_X6Y108_BO6),
.I4(CLBLL_L_X4Y109_SLICE_X5Y109_BO6),
.I5(CLBLM_R_X5Y108_SLICE_X6Y108_AO6),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_BO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h80f8f880f880f880)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(CLBLL_L_X4Y109_SLICE_X5Y109_BO6),
.I3(CLBLM_R_X7Y107_SLICE_X8Y107_CO6),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_AO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_DO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_CO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_BO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0cc00cc00)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_AO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_DO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffdfffffffff)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_CLUT (
.I0(CLBLM_R_X5Y109_SLICE_X6Y109_BO6),
.I1(CLBLM_R_X5Y108_SLICE_X6Y108_CO6),
.I2(CLBLM_R_X3Y108_SLICE_X3Y108_DO6),
.I3(CLBLM_R_X7Y109_SLICE_X9Y109_AO6),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I5(CLBLL_L_X4Y109_SLICE_X5Y109_AO5),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_CO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffbffff)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_BLUT (
.I0(CLBLM_R_X3Y108_SLICE_X3Y108_DO6),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(CLBLM_L_X8Y110_SLICE_X11Y110_BO6),
.I3(CLBLL_L_X4Y110_SLICE_X5Y110_AO6),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(CLBLL_L_X4Y109_SLICE_X5Y109_AO5),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_BO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6668666666666666)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_ALUT (
.I0(CLBLM_R_X3Y110_SLICE_X2Y110_DO6),
.I1(CLBLM_R_X3Y110_SLICE_X2Y110_BO6),
.I2(CLBLM_L_X8Y104_SLICE_X10Y104_CO6),
.I3(CLBLM_R_X5Y110_SLICE_X6Y110_BO6),
.I4(CLBLM_L_X10Y110_SLICE_X13Y110_AO6),
.I5(CLBLM_R_X7Y104_SLICE_X8Y104_AO5),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_AO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_DO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_CO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2baf175f030f3fff)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_BLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(CLBLM_R_X5Y108_SLICE_X6Y108_AO6),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(CLBLM_R_X7Y108_SLICE_X9Y108_BO6),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_BO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h96693cc35aa5f00f)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(CLBLM_R_X5Y108_SLICE_X6Y108_AO6),
.I3(CLBLM_R_X7Y108_SLICE_X9Y108_BO6),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_AO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9699aa556696aaaa)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_DLUT (
.I0(CLBLM_R_X7Y111_SLICE_X9Y111_BO6),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(CLBLM_R_X5Y111_SLICE_X6Y111_BO6),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_DO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996a55a996655aa)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_CLUT (
.I0(CLBLM_L_X8Y109_SLICE_X10Y109_BO6),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_R_X7Y108_SLICE_X9Y108_CO6),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_CO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heac0bf3f80002a00)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_BLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(CLBLM_L_X8Y109_SLICE_X10Y109_BO6),
.I5(CLBLM_R_X7Y108_SLICE_X9Y108_CO6),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_BO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ff000000)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(1'b1),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_AO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_DO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_CO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_BO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_AO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8c0e80080000000)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_DLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_DO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9548e2c0e2486ac0)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(CLBLM_R_X5Y112_SLICE_X6Y112_DO6),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_CO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0202000bbb3a2a0)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_BLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_BO6),
.I5(CLBLM_R_X7Y113_SLICE_X8Y113_AO5),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_BO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000aaaa0000)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(1'b1),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(1'b1),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_AO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_DO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_CO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_BO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aa00aa00)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_AO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1a7050f0a0808000)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_DLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(CLBLM_R_X5Y112_SLICE_X6Y112_DO6),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_DO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h336333c663ccc6cc)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_CLUT (
.I0(CLBLM_R_X7Y112_SLICE_X8Y112_AO6),
.I1(CLBLM_R_X5Y113_SLICE_X6Y113_DO6),
.I2(CLBLM_R_X5Y113_SLICE_X7Y113_BO6),
.I3(CLBLM_R_X5Y112_SLICE_X6Y112_CO6),
.I4(CLBLM_R_X7Y110_SLICE_X8Y110_DO6),
.I5(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_CO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee808000c8800000)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_BLUT (
.I0(CLBLM_R_X5Y112_SLICE_X6Y112_DO6),
.I1(RIOB33_X105Y111_IOB_X1Y111_I),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_BO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h66669999b44b2dd2)
  ) CLBLM_R_X5Y113_SLICE_X6Y113_ALUT (
.I0(CLBLM_R_X7Y110_SLICE_X8Y110_DO6),
.I1(CLBLM_R_X5Y113_SLICE_X7Y113_BO6),
.I2(CLBLM_R_X5Y112_SLICE_X6Y112_CO6),
.I3(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.I4(CLBLM_R_X7Y112_SLICE_X8Y112_AO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X6Y113_AO5),
.O6(CLBLM_R_X5Y113_SLICE_X6Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcf0fdf4c000d040)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_DLUT (
.I0(CLBLM_R_X5Y114_SLICE_X7Y114_AO5),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_BO6),
.I2(CLBLM_R_X7Y110_SLICE_X8Y110_DO6),
.I3(CLBLM_R_X5Y113_SLICE_X7Y113_AO5),
.I4(CLBLM_R_X5Y115_SLICE_X6Y115_DO6),
.I5(CLBLM_R_X7Y112_SLICE_X8Y112_AO6),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_DO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heaeaea80ea808080)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_CLUT (
.I0(CLBLM_R_X5Y113_SLICE_X6Y113_BO6),
.I1(RIOB33_X105Y111_IOB_X1Y111_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(CLBLM_R_X5Y112_SLICE_X6Y112_CO6),
.I4(CLBLM_R_X5Y113_SLICE_X7Y113_DO6),
.I5(CLBLM_R_X7Y112_SLICE_X8Y112_DO6),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_CO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1337377f01131337)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_BLUT (
.I0(CLBLM_R_X7Y110_SLICE_X8Y110_AO5),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_BO6),
.I2(CLBLM_R_X7Y114_SLICE_X8Y114_DO6),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_BO6),
.I4(CLBLM_R_X5Y112_SLICE_X7Y112_AO6),
.I5(CLBLM_R_X5Y115_SLICE_X6Y115_CO6),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_BO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5555aaafaaaa000)
  ) CLBLM_R_X5Y113_SLICE_X7Y113_ALUT (
.I0(CLBLM_R_X7Y110_SLICE_X8Y110_AO5),
.I1(1'b1),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_BO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y113_SLICE_X7Y113_AO5),
.O6(CLBLM_R_X5Y113_SLICE_X7Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_DO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_CO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd0f4f4fd40d0d0f4)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_BLUT (
.I0(CLBLL_L_X4Y114_SLICE_X5Y114_CO6),
.I1(CLBLM_R_X7Y113_SLICE_X9Y113_AO5),
.I2(CLBLM_R_X7Y114_SLICE_X8Y114_AO6),
.I3(CLBLL_L_X4Y113_SLICE_X4Y113_AO6),
.I4(CLBLM_R_X7Y113_SLICE_X8Y113_CO6),
.I5(CLBLL_L_X4Y114_SLICE_X4Y114_BO5),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_BO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h93936c6cb3b32020)
  ) CLBLM_R_X5Y114_SLICE_X6Y114_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLM_R_X7Y113_SLICE_X9Y113_AO5),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(1'b1),
.I4(CLBLM_R_X7Y113_SLICE_X8Y113_CO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y114_SLICE_X6Y114_AO5),
.O6(CLBLM_R_X5Y114_SLICE_X6Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_DO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_CO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_BO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff00ff0000f000f)
  ) CLBLM_R_X5Y114_SLICE_X7Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X5Y113_SLICE_X7Y113_AO6),
.I3(CLBLM_R_X7Y114_SLICE_X8Y114_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y114_SLICE_X7Y114_AO5),
.O6(CLBLM_R_X5Y114_SLICE_X7Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h004000d040f0d0f0)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_DLUT (
.I0(CLBLM_R_X5Y115_SLICE_X6Y115_AO6),
.I1(CLBLL_L_X4Y115_SLICE_X5Y115_BO6),
.I2(CLBLM_R_X5Y114_SLICE_X7Y114_AO6),
.I3(CLBLM_R_X5Y115_SLICE_X6Y115_AO5),
.I4(CLBLM_R_X5Y116_SLICE_X6Y116_AO5),
.I5(CLBLM_R_X7Y114_SLICE_X8Y114_CO6),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_DO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h002b02bf02bf2bff)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_CLUT (
.I0(CLBLL_L_X4Y115_SLICE_X5Y115_BO6),
.I1(CLBLM_R_X5Y115_SLICE_X7Y115_AO5),
.I2(CLBLM_R_X7Y115_SLICE_X8Y115_CO6),
.I3(CLBLM_R_X7Y114_SLICE_X8Y114_CO6),
.I4(CLBLM_R_X5Y116_SLICE_X6Y116_AO5),
.I5(CLBLM_R_X7Y115_SLICE_X8Y115_BO5),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_CO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a5965a965a965a)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_BLUT (
.I0(CLBLM_L_X8Y114_SLICE_X10Y114_BO6),
.I1(LIOB33_X0Y113_IOB_X0Y113_I),
.I2(CLBLM_R_X7Y114_SLICE_X9Y114_DO6),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(LIOB33_X0Y115_IOB_X0Y115_I),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_BO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aaaaaafcc0c0c0)
  ) CLBLM_R_X5Y115_SLICE_X6Y115_ALUT (
.I0(CLBLM_R_X7Y115_SLICE_X8Y115_DO6),
.I1(CLBLM_R_X7Y115_SLICE_X8Y115_CO6),
.I2(CLBLM_R_X7Y115_SLICE_X8Y115_BO5),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y115_SLICE_X6Y115_AO5),
.O6(CLBLM_R_X5Y115_SLICE_X6Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_DO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc33cccc33cc33)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_BO6),
.I2(1'b1),
.I3(CLBLM_R_X5Y113_SLICE_X7Y113_AO5),
.I4(1'b1),
.I5(CLBLM_R_X5Y115_SLICE_X7Y115_BO6),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_CO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h071f1f7f0107071f)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_BLUT (
.I0(CLBLM_R_X5Y115_SLICE_X6Y115_AO5),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_AO6),
.I2(CLBLM_R_X5Y113_SLICE_X7Y113_AO6),
.I3(CLBLM_R_X7Y115_SLICE_X8Y115_CO5),
.I4(CLBLM_R_X5Y115_SLICE_X7Y115_AO6),
.I5(CLBLM_R_X5Y116_SLICE_X6Y116_CO6),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_BO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000c0c0c0c0)
  ) CLBLM_R_X5Y115_SLICE_X7Y115_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y115_SLICE_X7Y115_AO5),
.O6(CLBLM_R_X5Y115_SLICE_X7Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5aa5a55a5aa5a5)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_DLUT (
.I0(CLBLM_R_X5Y115_SLICE_X6Y115_BO6),
.I1(1'b1),
.I2(CLBLM_R_X7Y114_SLICE_X8Y114_BO6),
.I3(1'b1),
.I4(CLBLM_R_X5Y114_SLICE_X6Y114_BO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_DO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1301371337137f37)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_CLUT (
.I0(CLBLM_R_X5Y116_SLICE_X6Y116_AO6),
.I1(CLBLM_R_X5Y115_SLICE_X6Y115_AO6),
.I2(CLBLM_R_X7Y114_SLICE_X8Y114_BO6),
.I3(CLBLM_R_X5Y114_SLICE_X6Y114_BO6),
.I4(CLBLM_R_X7Y114_SLICE_X9Y114_DO6),
.I5(CLBLM_R_X7Y115_SLICE_X8Y115_BO6),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_CO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd42b42bd42bd2bd4)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_BLUT (
.I0(CLBLM_R_X5Y114_SLICE_X6Y114_BO6),
.I1(CLBLM_R_X7Y114_SLICE_X9Y114_DO6),
.I2(CLBLM_R_X7Y115_SLICE_X8Y115_BO6),
.I3(CLBLM_R_X5Y115_SLICE_X6Y115_AO6),
.I4(CLBLM_R_X5Y116_SLICE_X6Y116_AO6),
.I5(CLBLM_R_X7Y114_SLICE_X8Y114_BO6),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_BO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00e8c0e8c0)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(CLBLM_R_X7Y114_SLICE_X9Y114_DO6),
.I2(CLBLM_R_X7Y115_SLICE_X8Y115_BO6),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_AO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_DO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_CO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_BO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_AO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h15d52ae63300cc00)
  ) CLBLM_R_X7Y102_SLICE_X8Y102_DLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(RIOB33_X105Y113_IOB_X1Y113_I),
.O5(CLBLM_R_X7Y102_SLICE_X8Y102_DO5),
.O6(CLBLM_R_X7Y102_SLICE_X8Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00f000f000)
  ) CLBLM_R_X7Y102_SLICE_X8Y102_CLUT (
.I0(1'b1),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y102_SLICE_X8Y102_CO5),
.O6(CLBLM_R_X7Y102_SLICE_X8Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4ccc4040d3531f9f)
  ) CLBLM_R_X7Y102_SLICE_X8Y102_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y102_SLICE_X8Y102_BO5),
.O6(CLBLM_R_X7Y102_SLICE_X8Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3cf0f0dd445500)
  ) CLBLM_R_X7Y102_SLICE_X8Y102_ALUT (
.I0(CLBLM_L_X8Y102_SLICE_X10Y102_AO5),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(CLBLM_R_X7Y102_SLICE_X8Y102_DO6),
.I3(CLBLM_R_X7Y102_SLICE_X8Y102_BO6),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y102_SLICE_X8Y102_AO5),
.O6(CLBLM_R_X7Y102_SLICE_X8Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h699966695555a5a5)
  ) CLBLM_R_X7Y102_SLICE_X9Y102_DLUT (
.I0(CLBLM_R_X7Y103_SLICE_X9Y103_AO6),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(CLBLM_R_X7Y102_SLICE_X8Y102_BO6),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(CLBLM_L_X8Y102_SLICE_X10Y102_AO5),
.I5(LIOB33_X0Y101_IOB_X0Y101_I),
.O5(CLBLM_R_X7Y102_SLICE_X9Y102_DO5),
.O6(CLBLM_R_X7Y102_SLICE_X9Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h80ecc8feec80fec8)
  ) CLBLM_R_X7Y102_SLICE_X9Y102_CLUT (
.I0(CLBLM_R_X7Y102_SLICE_X9Y102_AO6),
.I1(CLBLM_R_X7Y102_SLICE_X8Y102_CO6),
.I2(CLBLM_R_X7Y102_SLICE_X8Y102_BO6),
.I3(CLBLM_R_X7Y102_SLICE_X9Y102_AO5),
.I4(CLBLM_L_X8Y102_SLICE_X10Y102_AO5),
.I5(CLBLM_R_X7Y103_SLICE_X9Y103_AO6),
.O5(CLBLM_R_X7Y102_SLICE_X9Y102_CO5),
.O6(CLBLM_R_X7Y102_SLICE_X9Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd22d4bb42dd2b44b)
  ) CLBLM_R_X7Y102_SLICE_X9Y102_BLUT (
.I0(CLBLM_L_X8Y102_SLICE_X10Y102_AO5),
.I1(CLBLM_R_X7Y102_SLICE_X8Y102_BO6),
.I2(CLBLM_R_X7Y102_SLICE_X8Y102_CO6),
.I3(CLBLM_R_X7Y103_SLICE_X9Y103_AO6),
.I4(CLBLM_R_X7Y102_SLICE_X9Y102_AO6),
.I5(CLBLM_R_X7Y102_SLICE_X9Y102_AO5),
.O5(CLBLM_R_X7Y102_SLICE_X9Y102_BO5),
.O6(CLBLM_R_X7Y102_SLICE_X9Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ff000000)
  ) CLBLM_R_X7Y102_SLICE_X9Y102_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(1'b1),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y102_SLICE_X9Y102_AO5),
.O6(CLBLM_R_X7Y102_SLICE_X9Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y103_SLICE_X8Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y103_SLICE_X8Y103_DO5),
.O6(CLBLM_R_X7Y103_SLICE_X8Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y103_SLICE_X8Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y103_SLICE_X8Y103_CO5),
.O6(CLBLM_R_X7Y103_SLICE_X8Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h696655a5996955a5)
  ) CLBLM_R_X7Y103_SLICE_X8Y103_BLUT (
.I0(CLBLM_L_X8Y103_SLICE_X11Y103_AO6),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(CLBLM_R_X7Y102_SLICE_X8Y102_AO5),
.I3(CLBLM_L_X8Y103_SLICE_X10Y103_AO5),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(RIOB33_X105Y101_IOB_X1Y102_I),
.O5(CLBLM_R_X7Y103_SLICE_X8Y103_BO5),
.O6(CLBLM_R_X7Y103_SLICE_X8Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h693c96c3c3693c96)
  ) CLBLM_R_X7Y103_SLICE_X8Y103_ALUT (
.I0(CLBLM_R_X5Y102_SLICE_X7Y102_DO6),
.I1(CLBLM_L_X8Y102_SLICE_X11Y102_BO6),
.I2(CLBLM_R_X7Y104_SLICE_X8Y104_AO6),
.I3(CLBLM_R_X7Y102_SLICE_X9Y102_BO6),
.I4(CLBLM_R_X7Y102_SLICE_X9Y102_CO6),
.I5(CLBLM_R_X5Y103_SLICE_X6Y103_AO5),
.O5(CLBLM_R_X7Y103_SLICE_X8Y103_AO5),
.O6(CLBLM_R_X7Y103_SLICE_X8Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y103_SLICE_X9Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y103_SLICE_X9Y103_DO5),
.O6(CLBLM_R_X7Y103_SLICE_X9Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y103_SLICE_X9Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y103_SLICE_X9Y103_CO5),
.O6(CLBLM_R_X7Y103_SLICE_X9Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y103_SLICE_X9Y103_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y103_SLICE_X9Y103_BO5),
.O6(CLBLM_R_X7Y103_SLICE_X9Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf999a5a509c9ffff)
  ) CLBLM_R_X7Y103_SLICE_X9Y103_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O5(CLBLM_R_X7Y103_SLICE_X9Y103_AO5),
.O6(CLBLM_R_X7Y103_SLICE_X9Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff87870087870000)
  ) CLBLM_R_X7Y104_SLICE_X8Y104_DLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(CLBLM_R_X7Y102_SLICE_X9Y102_DO6),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLM_R_X5Y102_SLICE_X7Y102_DO6),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_R_X7Y104_SLICE_X8Y104_DO5),
.O6(CLBLM_R_X7Y104_SLICE_X8Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf9f5905099550000)
  ) CLBLM_R_X7Y104_SLICE_X8Y104_CLUT (
.I0(CLBLM_R_X7Y103_SLICE_X8Y103_BO6),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLM_R_X7Y104_SLICE_X8Y104_DO6),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_R_X7Y104_SLICE_X8Y104_CO5),
.O6(CLBLM_R_X7Y104_SLICE_X8Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h935f6ca06ca0935f)
  ) CLBLM_R_X7Y104_SLICE_X8Y104_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(CLBLM_L_X8Y103_SLICE_X11Y103_AO6),
.I5(CLBLM_R_X7Y102_SLICE_X9Y102_CO6),
.O5(CLBLM_R_X7Y104_SLICE_X8Y104_BO5),
.O6(CLBLM_R_X7Y104_SLICE_X8Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f00005555000)
  ) CLBLM_R_X7Y104_SLICE_X8Y104_ALUT (
.I0(CLBLM_R_X7Y104_SLICE_X8Y104_DO6),
.I1(1'b1),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLM_R_X7Y103_SLICE_X8Y103_BO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y104_SLICE_X8Y104_AO5),
.O6(CLBLM_R_X7Y104_SLICE_X8Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y104_SLICE_X9Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y104_SLICE_X9Y104_DO5),
.O6(CLBLM_R_X7Y104_SLICE_X9Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y104_SLICE_X9Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y104_SLICE_X9Y104_CO5),
.O6(CLBLM_R_X7Y104_SLICE_X9Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h650fa6009af059ff)
  ) CLBLM_R_X7Y104_SLICE_X9Y104_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(CLBLM_L_X8Y104_SLICE_X11Y104_AO6),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(CLBLM_R_X7Y104_SLICE_X9Y104_AO6),
.I5(CLBLM_L_X10Y104_SLICE_X12Y104_AO6),
.O5(CLBLM_R_X7Y104_SLICE_X9Y104_BO5),
.O6(CLBLM_R_X7Y104_SLICE_X9Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbe3cfaf02800a000)
  ) CLBLM_R_X7Y104_SLICE_X9Y104_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(CLBLM_L_X8Y103_SLICE_X11Y103_AO6),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLM_R_X7Y102_SLICE_X9Y102_CO6),
.O5(CLBLM_R_X7Y104_SLICE_X9Y104_AO5),
.O6(CLBLM_R_X7Y104_SLICE_X9Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y105_SLICE_X8Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y105_SLICE_X8Y105_DO5),
.O6(CLBLM_R_X7Y105_SLICE_X8Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hec80b320fec8fb32)
  ) CLBLM_R_X7Y105_SLICE_X8Y105_CLUT (
.I0(CLBLM_R_X5Y105_SLICE_X6Y105_AO5),
.I1(CLBLM_L_X8Y103_SLICE_X10Y103_BO6),
.I2(CLBLM_R_X7Y104_SLICE_X8Y104_DO6),
.I3(CLBLM_R_X7Y106_SLICE_X8Y106_AO5),
.I4(CLBLM_L_X8Y105_SLICE_X10Y105_AO6),
.I5(CLBLM_R_X7Y104_SLICE_X8Y104_BO6),
.O5(CLBLM_R_X7Y105_SLICE_X8Y105_CO5),
.O6(CLBLM_R_X7Y105_SLICE_X8Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h96c33c96693cc369)
  ) CLBLM_R_X7Y105_SLICE_X8Y105_BLUT (
.I0(CLBLM_R_X7Y104_SLICE_X8Y104_DO6),
.I1(CLBLM_L_X8Y103_SLICE_X10Y103_BO6),
.I2(CLBLM_L_X8Y105_SLICE_X10Y105_AO6),
.I3(CLBLM_R_X7Y104_SLICE_X8Y104_BO6),
.I4(CLBLM_R_X5Y105_SLICE_X6Y105_AO5),
.I5(CLBLM_R_X7Y106_SLICE_X8Y106_AO5),
.O5(CLBLM_R_X7Y105_SLICE_X8Y105_BO5),
.O6(CLBLM_R_X7Y105_SLICE_X8Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0f0f00000)
  ) CLBLM_R_X7Y105_SLICE_X8Y105_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(1'b1),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(1'b1),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y105_SLICE_X8Y105_AO5),
.O6(CLBLM_R_X7Y105_SLICE_X8Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y105_SLICE_X9Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y105_SLICE_X9Y105_DO5),
.O6(CLBLM_R_X7Y105_SLICE_X9Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y105_SLICE_X9Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y105_SLICE_X9Y105_CO5),
.O6(CLBLM_R_X7Y105_SLICE_X9Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y105_SLICE_X9Y105_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y105_SLICE_X9Y105_BO5),
.O6(CLBLM_R_X7Y105_SLICE_X9Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he47d6c5f1b8293a0)
  ) CLBLM_R_X7Y105_SLICE_X9Y105_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_L_X8Y104_SLICE_X10Y104_CO6),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_R_X7Y104_SLICE_X8Y104_CO6),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(CLBLM_R_X7Y104_SLICE_X9Y104_BO6),
.O5(CLBLM_R_X7Y105_SLICE_X9Y105_AO5),
.O6(CLBLM_R_X7Y105_SLICE_X9Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4c13df7f134c7fdf)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_DLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_L_X8Y104_SLICE_X10Y104_CO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(CLBLM_R_X7Y106_SLICE_X8Y106_AO5),
.I4(CLBLM_R_X5Y104_SLICE_X6Y104_DO6),
.I5(CLBLM_R_X7Y104_SLICE_X8Y104_CO6),
.O5(CLBLM_R_X7Y106_SLICE_X8Y106_DO5),
.O6(CLBLM_R_X7Y106_SLICE_X8Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h96693cc36996c33c)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_L_X8Y104_SLICE_X10Y104_CO6),
.I2(CLBLM_R_X5Y104_SLICE_X6Y104_DO6),
.I3(CLBLM_R_X7Y106_SLICE_X8Y106_AO5),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_R_X7Y104_SLICE_X8Y104_CO6),
.O5(CLBLM_R_X7Y106_SLICE_X8Y106_CO5),
.O6(CLBLM_R_X7Y106_SLICE_X8Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc33c966996693cc3)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_BLUT (
.I0(CLBLM_R_X5Y104_SLICE_X6Y104_DO6),
.I1(CLBLM_L_X8Y106_SLICE_X11Y106_AO6),
.I2(CLBLM_R_X7Y105_SLICE_X8Y105_CO6),
.I3(CLBLM_L_X8Y104_SLICE_X10Y104_AO6),
.I4(CLBLM_R_X7Y105_SLICE_X8Y105_BO6),
.I5(CLBLM_R_X5Y106_SLICE_X6Y106_AO5),
.O5(CLBLM_R_X7Y106_SLICE_X8Y106_BO5),
.O6(CLBLM_R_X7Y106_SLICE_X8Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h96695aa5cccc0000)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_ALUT (
.I0(CLBLM_R_X5Y104_SLICE_X6Y104_DO6),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(CLBLM_L_X8Y104_SLICE_X10Y104_CO6),
.I3(CLBLM_R_X7Y104_SLICE_X8Y104_CO6),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y106_SLICE_X8Y106_AO5),
.O6(CLBLM_R_X7Y106_SLICE_X8Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y106_SLICE_X9Y106_DO5),
.O6(CLBLM_R_X7Y106_SLICE_X9Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y106_SLICE_X9Y106_CO5),
.O6(CLBLM_R_X7Y106_SLICE_X9Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y106_SLICE_X9Y106_BO5),
.O6(CLBLM_R_X7Y106_SLICE_X9Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h80008880a888ffa8)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_R_X7Y104_SLICE_X8Y104_CO6),
.I4(CLBLM_L_X8Y104_SLICE_X10Y104_CO6),
.I5(CLBLM_L_X8Y104_SLICE_X10Y104_AO6),
.O5(CLBLM_R_X7Y106_SLICE_X9Y106_AO5),
.O6(CLBLM_R_X7Y106_SLICE_X9Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdeee48885aaa0000)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_DLUT (
.I0(CLBLM_R_X7Y106_SLICE_X8Y106_AO6),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_R_X5Y106_SLICE_X6Y106_DO6),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLM_R_X7Y107_SLICE_X8Y107_DO5),
.O6(CLBLM_R_X7Y107_SLICE_X8Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha569695a5a9696a5)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_CLUT (
.I0(CLBLM_L_X8Y107_SLICE_X10Y107_BO6),
.I1(CLBLM_R_X7Y107_SLICE_X9Y107_AO6),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_BO6),
.I3(CLBLM_R_X7Y107_SLICE_X8Y107_AO5),
.I4(CLBLM_R_X7Y107_SLICE_X8Y107_DO6),
.I5(CLBLM_R_X7Y108_SLICE_X9Y108_AO6),
.O5(CLBLM_R_X7Y107_SLICE_X8Y107_CO5),
.O6(CLBLM_R_X7Y107_SLICE_X8Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2112a55a03300ff0)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(CLBLM_R_X7Y106_SLICE_X8Y106_AO6),
.I3(CLBLM_R_X5Y106_SLICE_X6Y106_DO6),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X7Y107_SLICE_X8Y107_BO5),
.O6(CLBLM_R_X7Y107_SLICE_X8Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00f000f000)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(1'b1),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y107_SLICE_X8Y107_AO5),
.O6(CLBLM_R_X7Y107_SLICE_X8Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8f707f80e51a15ea)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_DLUT (
.I0(CLBLM_R_X7Y104_SLICE_X8Y104_CO6),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLM_L_X8Y104_SLICE_X10Y104_AO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_L_X8Y104_SLICE_X10Y104_CO6),
.O5(CLBLM_R_X7Y107_SLICE_X9Y107_DO5),
.O6(CLBLM_R_X7Y107_SLICE_X9Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h96a55a96695aa569)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_CLUT (
.I0(CLBLM_R_X7Y108_SLICE_X9Y108_AO6),
.I1(CLBLM_R_X7Y106_SLICE_X8Y106_DO6),
.I2(CLBLM_L_X8Y108_SLICE_X10Y108_AO6),
.I3(CLBLM_R_X7Y109_SLICE_X8Y109_AO6),
.I4(CLBLM_R_X7Y107_SLICE_X9Y107_DO6),
.I5(CLBLM_L_X8Y107_SLICE_X10Y107_CO6),
.O5(CLBLM_R_X7Y107_SLICE_X9Y107_CO5),
.O6(CLBLM_R_X7Y107_SLICE_X9Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb7213f0321210303)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLM_R_X7Y106_SLICE_X8Y106_DO6),
.I2(CLBLM_R_X7Y105_SLICE_X9Y105_AO6),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X7Y107_SLICE_X9Y107_BO5),
.O6(CLBLM_R_X7Y107_SLICE_X9Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h96693cc36969c3c3)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLM_R_X7Y106_SLICE_X8Y106_DO6),
.I2(CLBLM_R_X7Y105_SLICE_X9Y105_AO6),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X7Y107_SLICE_X9Y107_AO5),
.O6(CLBLM_R_X7Y107_SLICE_X9Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_DO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7130f37117033f17)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_CLUT (
.I0(CLBLM_R_X5Y106_SLICE_X6Y106_DO6),
.I1(CLBLM_R_X7Y107_SLICE_X8Y107_AO5),
.I2(CLBLM_R_X7Y106_SLICE_X8Y106_BO6),
.I3(CLBLM_R_X7Y106_SLICE_X8Y106_CO6),
.I4(CLBLM_R_X5Y107_SLICE_X6Y107_AO5),
.I5(CLBLM_R_X7Y109_SLICE_X8Y109_AO6),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_CO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h965aa596aaaa55aa)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_BLUT (
.I0(CLBLM_L_X8Y108_SLICE_X10Y108_CO6),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(CLBLM_R_X7Y107_SLICE_X9Y107_BO6),
.I4(CLBLM_L_X8Y107_SLICE_X10Y107_BO6),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_BO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h956aa9566a9556a9)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_ALUT (
.I0(CLBLM_R_X7Y107_SLICE_X8Y107_AO5),
.I1(CLBLM_R_X5Y107_SLICE_X6Y107_AO5),
.I2(CLBLM_R_X5Y106_SLICE_X6Y106_DO6),
.I3(CLBLM_R_X7Y106_SLICE_X8Y106_BO6),
.I4(CLBLM_R_X7Y106_SLICE_X8Y106_CO6),
.I5(CLBLM_R_X7Y109_SLICE_X8Y109_AO6),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_AO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_DO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8eaf000c0a8e000c)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_CLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(CLBLM_R_X7Y107_SLICE_X9Y107_BO6),
.I2(CLBLM_L_X8Y108_SLICE_X10Y108_CO6),
.I3(CLBLM_L_X8Y107_SLICE_X10Y107_BO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_CO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h650c9af3a60c59f3)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(CLBLM_R_X7Y107_SLICE_X9Y107_BO6),
.I2(CLBLM_L_X8Y107_SLICE_X10Y107_BO6),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(CLBLM_L_X8Y108_SLICE_X10Y108_BO6),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_BO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00cc00cc00)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_AO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000008000)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_DLUT (
.I0(CLBLM_R_X7Y104_SLICE_X8Y104_AO5),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(CLBLM_R_X11Y106_SLICE_X14Y106_BO6),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_DO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc63939c6639c9c63)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_CLUT (
.I0(CLBLM_R_X7Y108_SLICE_X8Y108_BO6),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I2(CLBLM_R_X5Y108_SLICE_X6Y108_AO6),
.I3(CLBLM_R_X7Y108_SLICE_X9Y108_CO6),
.I4(CLBLM_R_X7Y109_SLICE_X8Y109_BO5),
.I5(CLBLM_R_X7Y109_SLICE_X8Y109_BO6),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_CO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0cc00cc00)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_BO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00f000f000)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_AO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00cc00cc00)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_DLUT (
.I0(1'b1),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(1'b1),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_DO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heafe80a8d5fd4054)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_CLUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_AO6),
.I1(CLBLM_R_X7Y108_SLICE_X9Y108_CO6),
.I2(CLBLM_R_X7Y109_SLICE_X8Y109_BO5),
.I3(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I4(CLBLM_R_X7Y109_SLICE_X9Y109_DO6),
.I5(CLBLM_L_X8Y109_SLICE_X10Y109_CO6),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_CO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6696996996996966)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_BLUT (
.I0(CLBLM_R_X7Y109_SLICE_X9Y109_DO6),
.I1(CLBLM_L_X8Y109_SLICE_X10Y109_CO6),
.I2(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.I3(CLBLM_R_X7Y109_SLICE_X8Y109_BO5),
.I4(CLBLM_R_X7Y111_SLICE_X8Y111_AO6),
.I5(CLBLM_R_X7Y108_SLICE_X9Y108_CO6),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_BO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h96d24488f0788888)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_ALUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(RIOB33_X105Y111_IOB_X1Y111_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(CLBLM_L_X8Y110_SLICE_X11Y110_DO6),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_AO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa88a880f8808800)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_DLUT (
.I0(RIOB33_X105Y107_IOB_X1Y108_I),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(CLBLM_R_X7Y110_SLICE_X9Y110_DO6),
.I3(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I4(CLBLM_R_X7Y111_SLICE_X9Y111_DO6),
.I5(LIOB33_X0Y113_IOB_X0Y113_I),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_DO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996969699666666)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_CLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I1(CLBLM_R_X7Y110_SLICE_X9Y110_CO6),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(LIOB33_X0Y113_IOB_X0Y113_I),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_CO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he817777717e88888)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_BLUT (
.I0(CLBLM_R_X7Y111_SLICE_X9Y111_DO6),
.I1(CLBLM_R_X7Y110_SLICE_X9Y110_DO6),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_BO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f00096966666)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_ALUT (
.I0(CLBLM_R_X7Y111_SLICE_X9Y111_DO6),
.I1(CLBLM_R_X7Y110_SLICE_X9Y110_DO6),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_AO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887887787787788)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_DLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(CLBLM_R_X7Y110_SLICE_X9Y110_AO5),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(CLBLM_R_X7Y110_SLICE_X9Y110_BO6),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_DO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7707700f8808800)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_CLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(CLBLM_R_X7Y110_SLICE_X9Y110_AO5),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(CLBLM_R_X7Y110_SLICE_X9Y110_BO6),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_CO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h462aa80022aa8000)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_BLUT (
.I0(RIOB33_X105Y111_IOB_X1Y111_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLM_L_X8Y110_SLICE_X11Y110_DO6),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_BO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h93936c6cecec8080)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_ALUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(CLBLM_L_X10Y110_SLICE_X13Y110_DO6),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(1'b1),
.I4(CLBLM_R_X7Y109_SLICE_X9Y109_AO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_AO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf9909090f5505050)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_DLUT (
.I0(CLBLM_L_X8Y111_SLICE_X10Y111_BO6),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_CO6),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_DO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996969669696996)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_CLUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_AO6),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_DO6),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_CO6),
.I3(CLBLM_R_X7Y108_SLICE_X9Y108_CO6),
.I4(CLBLM_R_X7Y109_SLICE_X8Y109_BO5),
.I5(CLBLM_L_X8Y110_SLICE_X10Y110_BO6),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_CO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a5965a965a965a)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_BLUT (
.I0(CLBLM_L_X8Y111_SLICE_X10Y111_CO6),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_BO6),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(RIOB33_X105Y101_IOB_X1Y102_I),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_BO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0aa00aa00)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(1'b1),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_AO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heca8e8a0c8808800)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_DLUT (
.I0(CLBLM_R_X7Y110_SLICE_X9Y110_AO6),
.I1(RIOB33_X105Y107_IOB_X1Y108_I),
.I2(CLBLM_R_X11Y111_SLICE_X14Y111_DO6),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(CLBLM_L_X10Y111_SLICE_X13Y111_CO6),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_DO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha956956a6a6a6a6a)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_CLUT (
.I0(CLBLM_R_X7Y110_SLICE_X9Y110_AO6),
.I1(CLBLM_L_X10Y111_SLICE_X13Y111_CO6),
.I2(CLBLM_R_X11Y111_SLICE_X14Y111_DO6),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(RIOB33_X105Y107_IOB_X1Y108_I),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_CO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93936c36c9c936)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_BLUT (
.I0(CLBLM_L_X8Y111_SLICE_X10Y111_CO6),
.I1(CLBLM_L_X8Y110_SLICE_X10Y110_AO6),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_AO6),
.I3(CLBLM_L_X10Y112_SLICE_X12Y112_BO6),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_AO6),
.I5(CLBLM_L_X8Y111_SLICE_X10Y111_DO6),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_BO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0995566aa)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_ALUT (
.I0(CLBLM_L_X8Y111_SLICE_X11Y111_DO6),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(CLBLM_L_X8Y111_SLICE_X11Y111_BO5),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_AO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb3ecffa02080a000)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_DLUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(CLBLM_R_X7Y112_SLICE_X8Y112_CO6),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(CLBLM_R_X7Y112_SLICE_X8Y112_BO6),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_DO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c7070f0e0800000)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_CLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_CO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6606600fcc0cc00)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_BLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_DO6),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(CLBLM_R_X7Y110_SLICE_X9Y110_CO6),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(RIOB33_X105Y109_IOB_X1Y110_I),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_BO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a95c03f956a3fc0)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(CLBLM_R_X7Y112_SLICE_X8Y112_BO6),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(CLBLM_R_X7Y112_SLICE_X8Y112_CO6),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_AO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1a70c0001a70c000)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_DLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_DO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfec0880080000000)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_CLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(CLBLM_L_X8Y110_SLICE_X11Y110_DO6),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_CO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffe8e800a000a000)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_BLUT (
.I0(CLBLM_L_X8Y111_SLICE_X11Y111_BO5),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(CLBLM_L_X8Y111_SLICE_X11Y111_DO6),
.I3(CLBLM_R_X7Y111_SLICE_X9Y111_CO6),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(RIOB33_X105Y107_IOB_X1Y107_I),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_BO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he11e55aa8778ff00)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_ALUT (
.I0(CLBLM_L_X8Y111_SLICE_X11Y111_DO6),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(CLBLM_R_X7Y111_SLICE_X9Y111_CO6),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(CLBLM_L_X8Y111_SLICE_X11Y111_BO5),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_AO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h936c6c936c93936c)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_DLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_R_X7Y111_SLICE_X8Y111_AO5),
.I4(CLBLM_R_X7Y109_SLICE_X9Y109_CO6),
.I5(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_DO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb3200000fb323030)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_CLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_AO6),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_CO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8778788777888877)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_L_X8Y112_SLICE_X11Y112_AO6),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_AO6),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_BO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c36cc66a55a55aa)
  ) CLBLM_R_X7Y113_SLICE_X8Y113_ALUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I1(CLBLM_L_X8Y113_SLICE_X10Y113_AO6),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLM_R_X7Y113_SLICE_X8Y113_BO6),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y113_SLICE_X8Y113_AO5),
.O6(CLBLM_R_X7Y113_SLICE_X8Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha220a000bab0b230)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y112_SLICE_X13Y112_DO6),
.I2(CLBLM_L_X8Y110_SLICE_X11Y110_AO5),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(CLBLM_L_X10Y113_SLICE_X12Y113_AO5),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_DO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc93636c9936c6c93)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_CLUT (
.I0(CLBLM_R_X7Y114_SLICE_X9Y114_AO6),
.I1(CLBLM_L_X10Y113_SLICE_X12Y113_CO6),
.I2(CLBLM_L_X10Y112_SLICE_X12Y112_CO6),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_AO5),
.I4(CLBLM_R_X7Y113_SLICE_X9Y113_BO5),
.I5(CLBLM_L_X10Y112_SLICE_X13Y112_CO6),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_CO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3cc33f0f00000)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y113_SLICE_X12Y113_AO5),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(CLBLM_L_X10Y112_SLICE_X13Y112_DO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_BO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f000005a5aaaaa)
  ) CLBLM_R_X7Y113_SLICE_X9Y113_ALUT (
.I0(CLBLM_L_X8Y113_SLICE_X10Y113_BO6),
.I1(1'b1),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(1'b1),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y113_SLICE_X9Y113_AO5),
.O6(CLBLM_R_X7Y113_SLICE_X9Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heaeac880c8808080)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_DLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_AO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(CLBLM_R_X7Y113_SLICE_X9Y113_DO6),
.I5(CLBLM_R_X7Y111_SLICE_X9Y111_AO5),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_DO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9595a66aa66a6a6a)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_CLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_AO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(CLBLM_R_X7Y113_SLICE_X9Y113_DO6),
.I5(CLBLM_R_X7Y111_SLICE_X9Y111_AO5),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_CO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h60f60066c0fc00cc)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(CLBLM_R_X7Y114_SLICE_X9Y114_BO6),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_L_X8Y113_SLICE_X10Y113_CO6),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_BO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c939393936c6c6c)
  ) CLBLM_R_X7Y114_SLICE_X8Y114_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLM_R_X7Y114_SLICE_X9Y114_BO6),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(CLBLM_L_X8Y113_SLICE_X10Y113_CO6),
.O5(CLBLM_R_X7Y114_SLICE_X8Y114_AO5),
.O6(CLBLM_R_X7Y114_SLICE_X8Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3b0b03033202000)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_DLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(CLBLM_R_X7Y113_SLICE_X9Y113_CO6),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(CLBLM_R_X7Y114_SLICE_X9Y114_AO5),
.I4(CLBLM_L_X8Y112_SLICE_X10Y112_DO6),
.I5(LIOB33_X0Y113_IOB_X0Y113_I),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_DO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha99533ff566acc00)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y112_SLICE_X12Y112_CO6),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(CLBLM_L_X10Y112_SLICE_X13Y112_CO6),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(CLBLM_L_X10Y113_SLICE_X12Y113_CO6),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_CO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he5151aea8f7f7080)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_BLUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_DO6),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(CLBLM_R_X7Y114_SLICE_X9Y114_CO6),
.I5(CLBLM_R_X7Y114_SLICE_X9Y114_AO5),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_BO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00993366cc)
  ) CLBLM_R_X7Y114_SLICE_X9Y114_ALUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(CLBLM_L_X10Y112_SLICE_X12Y112_CO6),
.I2(1'b1),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(CLBLM_L_X10Y112_SLICE_X13Y112_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y114_SLICE_X9Y114_AO5),
.O6(CLBLM_R_X7Y114_SLICE_X9Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc369966996c33c)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_DLUT (
.I0(CLBLM_R_X7Y115_SLICE_X8Y115_AO6),
.I1(CLBLM_R_X7Y111_SLICE_X9Y111_AO5),
.I2(CLBLM_R_X7Y113_SLICE_X9Y113_DO6),
.I3(CLBLM_R_X7Y115_SLICE_X8Y115_AO5),
.I4(CLBLM_L_X8Y114_SLICE_X10Y114_BO5),
.I5(CLBLM_L_X8Y114_SLICE_X10Y114_CO6),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_DO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h87788778f880f880)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y113_SLICE_X9Y113_DO6),
.I3(CLBLM_R_X7Y111_SLICE_X9Y111_AO5),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_CO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3cccccfaa0aa00)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_BLUT (
.I0(CLBLM_L_X8Y114_SLICE_X10Y114_BO5),
.I1(CLBLM_L_X8Y114_SLICE_X10Y114_BO6),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(CLBLM_L_X8Y114_SLICE_X10Y114_CO6),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_BO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000cccc0000)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_AO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_DO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_CO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_BO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_AO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y104_SLICE_X14Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y104_SLICE_X14Y104_DO5),
.O6(CLBLM_R_X11Y104_SLICE_X14Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y104_SLICE_X14Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y104_SLICE_X14Y104_CO5),
.O6(CLBLM_R_X11Y104_SLICE_X14Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y104_SLICE_X14Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y104_SLICE_X14Y104_BO5),
.O6(CLBLM_R_X11Y104_SLICE_X14Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf757775787d727d7)
  ) CLBLM_R_X11Y104_SLICE_X14Y104_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y104_SLICE_X14Y104_AO5),
.O6(CLBLM_R_X11Y104_SLICE_X14Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y104_SLICE_X15Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y104_SLICE_X15Y104_DO5),
.O6(CLBLM_R_X11Y104_SLICE_X15Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y104_SLICE_X15Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y104_SLICE_X15Y104_CO5),
.O6(CLBLM_R_X11Y104_SLICE_X15Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y104_SLICE_X15Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y104_SLICE_X15Y104_BO5),
.O6(CLBLM_R_X11Y104_SLICE_X15Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y104_SLICE_X15Y104_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y104_SLICE_X15Y104_AO5),
.O6(CLBLM_R_X11Y104_SLICE_X15Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h39c6c6399c63639c)
  ) CLBLM_R_X11Y105_SLICE_X14Y105_DLUT (
.I0(CLBLM_R_X7Y111_SLICE_X9Y111_AO6),
.I1(CLBLM_R_X11Y107_SLICE_X15Y107_AO5),
.I2(CLBLM_R_X11Y105_SLICE_X15Y105_AO6),
.I3(CLBLM_R_X11Y105_SLICE_X14Y105_AO5),
.I4(CLBLM_R_X11Y106_SLICE_X15Y106_BO6),
.I5(CLBLM_R_X11Y106_SLICE_X15Y106_AO5),
.O5(CLBLM_R_X11Y105_SLICE_X14Y105_DO5),
.O6(CLBLM_R_X11Y105_SLICE_X14Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6cc936c993c9c9c9)
  ) CLBLM_R_X11Y105_SLICE_X14Y105_CLUT (
.I0(CLBLM_R_X11Y105_SLICE_X14Y105_AO6),
.I1(CLBLM_R_X11Y105_SLICE_X15Y105_CO6),
.I2(CLBLM_L_X10Y104_SLICE_X13Y104_BO5),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(RIOB33_X105Y107_IOB_X1Y107_I),
.O5(CLBLM_R_X11Y105_SLICE_X14Y105_CO5),
.O6(CLBLM_R_X11Y105_SLICE_X14Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6fff666f06660006)
  ) CLBLM_R_X11Y105_SLICE_X14Y105_BLUT (
.I0(CLBLM_R_X11Y106_SLICE_X15Y106_BO6),
.I1(CLBLM_R_X11Y107_SLICE_X15Y107_AO5),
.I2(CLBLM_R_X11Y105_SLICE_X15Y105_AO6),
.I3(CLBLM_R_X11Y106_SLICE_X15Y106_AO5),
.I4(CLBLM_R_X7Y111_SLICE_X9Y111_AO6),
.I5(CLBLM_R_X11Y105_SLICE_X14Y105_AO5),
.O5(CLBLM_R_X11Y105_SLICE_X14Y105_BO5),
.O6(CLBLM_R_X11Y105_SLICE_X14Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa555555f000f000)
  ) CLBLM_R_X11Y105_SLICE_X14Y105_ALUT (
.I0(CLBLM_L_X10Y106_SLICE_X13Y106_AO6),
.I1(1'b1),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y105_SLICE_X14Y105_AO5),
.O6(CLBLM_R_X11Y105_SLICE_X14Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y105_SLICE_X15Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y105_SLICE_X15Y105_DO5),
.O6(CLBLM_R_X11Y105_SLICE_X15Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4bd2f0a5b42df0a5)
  ) CLBLM_R_X11Y105_SLICE_X15Y105_CLUT (
.I0(CLBLM_R_X11Y105_SLICE_X15Y105_AO6),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(CLBLM_R_X11Y106_SLICE_X15Y106_BO6),
.I3(CLBLM_R_X11Y106_SLICE_X15Y106_AO5),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(RIOB33_X105Y107_IOB_X1Y108_I),
.O5(CLBLM_R_X11Y105_SLICE_X15Y105_CO5),
.O6(CLBLM_R_X11Y105_SLICE_X15Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888a0a0a0a0)
  ) CLBLM_R_X11Y105_SLICE_X15Y105_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y105_SLICE_X15Y105_BO5),
.O6(CLBLM_R_X11Y105_SLICE_X15Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbf1f3f1f959f359f)
  ) CLBLM_R_X11Y105_SLICE_X15Y105_ALUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y105_SLICE_X15Y105_AO5),
.O6(CLBLM_R_X11Y105_SLICE_X15Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbd95426a173fe8c0)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_DLUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(CLBLM_R_X11Y106_SLICE_X15Y106_AO6),
.I2(CLBLM_R_X11Y107_SLICE_X14Y107_BO6),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(CLBLM_L_X12Y107_SLICE_X16Y107_AO6),
.I5(RIOB33_X105Y109_IOB_X1Y109_I),
.O5(CLBLM_R_X11Y106_SLICE_X14Y106_DO5),
.O6(CLBLM_R_X11Y106_SLICE_X14Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb222e888faaaa000)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_CLUT (
.I0(CLBLM_R_X11Y105_SLICE_X14Y105_BO6),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(CLBLM_R_X11Y106_SLICE_X14Y106_DO6),
.I5(RIOB33_X105Y107_IOB_X1Y108_I),
.O5(CLBLM_R_X11Y106_SLICE_X14Y106_CO5),
.O6(CLBLM_R_X11Y106_SLICE_X14Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h966669995aaaa555)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_BLUT (
.I0(CLBLM_R_X11Y106_SLICE_X14Y106_DO6),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(CLBLM_R_X11Y105_SLICE_X14Y105_BO6),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_R_X11Y106_SLICE_X14Y106_BO5),
.O6(CLBLM_R_X11Y106_SLICE_X14Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbf3f2a007fff153f)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y105_SLICE_X12Y105_AO6),
.I5(CLBLM_R_X11Y105_SLICE_X14Y105_CO6),
.O5(CLBLM_R_X11Y106_SLICE_X14Y106_AO5),
.O6(CLBLM_R_X11Y106_SLICE_X14Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y106_SLICE_X15Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y106_SLICE_X15Y106_DO5),
.O6(CLBLM_R_X11Y106_SLICE_X15Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y106_SLICE_X15Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y106_SLICE_X15Y106_CO5),
.O6(CLBLM_R_X11Y106_SLICE_X15Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hedc321ffa5c3a9ff)
  ) CLBLM_R_X11Y106_SLICE_X15Y106_BLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_R_X11Y106_SLICE_X15Y106_BO5),
.O6(CLBLM_R_X11Y106_SLICE_X15Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7030f0004cbcf000)
  ) CLBLM_R_X11Y106_SLICE_X15Y106_ALUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y106_SLICE_X15Y106_AO5),
.O6(CLBLM_R_X11Y106_SLICE_X15Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa569966996a55a)
  ) CLBLM_R_X11Y107_SLICE_X14Y107_DLUT (
.I0(CLBLM_R_X11Y107_SLICE_X15Y107_BO6),
.I1(CLBLM_R_X11Y107_SLICE_X15Y107_AO5),
.I2(CLBLM_L_X12Y107_SLICE_X16Y107_AO6),
.I3(CLBLM_R_X7Y110_SLICE_X8Y110_AO6),
.I4(CLBLM_R_X11Y106_SLICE_X15Y106_AO6),
.I5(CLBLM_R_X11Y107_SLICE_X14Y107_BO6),
.O5(CLBLM_R_X11Y107_SLICE_X14Y107_DO5),
.O6(CLBLM_R_X11Y107_SLICE_X14Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff5ade48de485a00)
  ) CLBLM_R_X11Y107_SLICE_X14Y107_CLUT (
.I0(CLBLM_R_X11Y107_SLICE_X15Y107_BO6),
.I1(CLBLM_R_X11Y107_SLICE_X15Y107_AO5),
.I2(CLBLM_L_X12Y107_SLICE_X16Y107_AO6),
.I3(CLBLM_R_X7Y110_SLICE_X8Y110_AO6),
.I4(CLBLM_R_X11Y106_SLICE_X15Y106_AO6),
.I5(CLBLM_R_X11Y107_SLICE_X14Y107_BO6),
.O5(CLBLM_R_X11Y107_SLICE_X14Y107_CO5),
.O6(CLBLM_R_X11Y107_SLICE_X14Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd05f2f5f7f005000)
  ) CLBLM_R_X11Y107_SLICE_X14Y107_BLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y107_SLICE_X14Y107_BO5),
.O6(CLBLM_R_X11Y107_SLICE_X14Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he8c0e8c069c369c3)
  ) CLBLM_R_X11Y107_SLICE_X14Y107_ALUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(CLBLM_R_X11Y106_SLICE_X14Y106_CO6),
.I2(CLBLM_R_X11Y107_SLICE_X15Y107_CO6),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y107_SLICE_X14Y107_AO5),
.O6(CLBLM_R_X11Y107_SLICE_X14Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfec8ec8088880000)
  ) CLBLM_R_X11Y107_SLICE_X15Y107_DLUT (
.I0(CLBLM_R_X11Y107_SLICE_X15Y107_AO6),
.I1(CLBLM_L_X10Y107_SLICE_X12Y107_AO6),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLM_R_X11Y107_SLICE_X15Y107_BO5),
.I5(RIOB33_X105Y107_IOB_X1Y108_I),
.O5(CLBLM_R_X11Y107_SLICE_X15Y107_DO5),
.O6(CLBLM_R_X11Y107_SLICE_X15Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc936936c55aaff00)
  ) CLBLM_R_X11Y107_SLICE_X15Y107_CLUT (
.I0(CLBLM_R_X11Y107_SLICE_X15Y107_AO6),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(CLBLM_L_X10Y107_SLICE_X12Y107_AO6),
.I4(CLBLM_R_X11Y107_SLICE_X15Y107_BO5),
.I5(RIOB33_X105Y107_IOB_X1Y108_I),
.O5(CLBLM_R_X11Y107_SLICE_X15Y107_CO5),
.O6(CLBLM_R_X11Y107_SLICE_X15Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc0033ffcc00)
  ) CLBLM_R_X11Y107_SLICE_X15Y107_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(1'b1),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(CLBLM_L_X12Y107_SLICE_X16Y107_AO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y107_SLICE_X15Y107_BO5),
.O6(CLBLM_R_X11Y107_SLICE_X15Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee888888ff000000)
  ) CLBLM_R_X11Y107_SLICE_X15Y107_ALUT (
.I0(CLBLM_R_X11Y106_SLICE_X15Y106_AO6),
.I1(CLBLM_R_X11Y107_SLICE_X14Y107_BO6),
.I2(1'b1),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y107_SLICE_X15Y107_AO5),
.O6(CLBLM_R_X11Y107_SLICE_X15Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc396963c3c6969c3)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_DLUT (
.I0(CLBLM_R_X11Y106_SLICE_X14Y106_CO6),
.I1(CLBLM_R_X11Y108_SLICE_X15Y108_AO5),
.I2(CLBLM_R_X11Y105_SLICE_X15Y105_BO6),
.I3(CLBLM_R_X11Y107_SLICE_X15Y107_CO6),
.I4(CLBLM_L_X10Y108_SLICE_X13Y108_AO6),
.I5(CLBLM_R_X11Y108_SLICE_X14Y108_BO6),
.O5(CLBLM_R_X11Y108_SLICE_X14Y108_DO5),
.O6(CLBLM_R_X11Y108_SLICE_X14Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3b2b230fce8e8c0)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_CLUT (
.I0(CLBLM_R_X11Y106_SLICE_X14Y106_CO6),
.I1(CLBLM_R_X11Y108_SLICE_X15Y108_AO5),
.I2(CLBLM_R_X11Y105_SLICE_X15Y105_BO6),
.I3(CLBLM_R_X11Y107_SLICE_X15Y107_CO6),
.I4(CLBLM_L_X10Y108_SLICE_X13Y108_AO6),
.I5(CLBLM_R_X11Y108_SLICE_X14Y108_BO6),
.O5(CLBLM_R_X11Y108_SLICE_X14Y108_CO5),
.O6(CLBLM_R_X11Y108_SLICE_X14Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h36c9c9366c93936c)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_BLUT (
.I0(CLBLM_R_X11Y107_SLICE_X14Y107_CO6),
.I1(CLBLM_L_X10Y107_SLICE_X12Y107_BO6),
.I2(CLBLM_L_X8Y111_SLICE_X11Y111_BO6),
.I3(CLBLM_L_X10Y108_SLICE_X12Y108_DO6),
.I4(CLBLM_R_X11Y110_SLICE_X15Y110_AO6),
.I5(CLBLM_L_X10Y107_SLICE_X12Y107_AO6),
.O5(CLBLM_R_X11Y108_SLICE_X14Y108_BO5),
.O6(CLBLM_R_X11Y108_SLICE_X14Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5559a6a9a6a5aaa)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_ALUT (
.I0(CLBLM_R_X11Y108_SLICE_X14Y108_BO6),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(CLBLM_R_X11Y106_SLICE_X14Y106_CO6),
.I5(CLBLM_R_X11Y107_SLICE_X15Y107_CO6),
.O5(CLBLM_R_X11Y108_SLICE_X14Y108_AO5),
.O6(CLBLM_R_X11Y108_SLICE_X14Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc366966696cc3ccc)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_DLUT (
.I0(CLBLM_R_X11Y110_SLICE_X15Y110_AO6),
.I1(CLBLM_L_X12Y108_SLICE_X16Y108_BO6),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(CLBLM_L_X10Y107_SLICE_X12Y107_BO6),
.O5(CLBLM_R_X11Y108_SLICE_X15Y108_DO5),
.O6(CLBLM_R_X11Y108_SLICE_X15Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996996696966666)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_CLUT (
.I0(CLBLM_L_X10Y107_SLICE_X12Y107_BO6),
.I1(CLBLM_R_X11Y110_SLICE_X15Y110_BO6),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_R_X11Y108_SLICE_X15Y108_CO5),
.O6(CLBLM_R_X11Y108_SLICE_X15Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc8c8c0c0808000)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(CLBLM_L_X10Y107_SLICE_X12Y107_BO6),
.I4(CLBLM_R_X11Y110_SLICE_X15Y110_AO6),
.I5(CLBLM_L_X12Y108_SLICE_X16Y108_BO6),
.O5(CLBLM_R_X11Y108_SLICE_X15Y108_BO5),
.O6(CLBLM_R_X11Y108_SLICE_X15Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h95956a6ac0c0c0c0)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_ALUT (
.I0(CLBLM_R_X11Y107_SLICE_X15Y107_DO6),
.I1(RIOB33_X105Y107_IOB_X1Y108_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(1'b1),
.I4(CLBLM_R_X11Y108_SLICE_X15Y108_CO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y108_SLICE_X15Y108_AO5),
.O6(CLBLM_R_X11Y108_SLICE_X15Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd42b2bd4af50af50)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_DLUT (
.I0(CLBLM_R_X11Y106_SLICE_X14Y106_AO6),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(CLBLM_L_X10Y109_SLICE_X13Y109_AO5),
.I3(CLBLM_L_X10Y108_SLICE_X13Y108_CO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_R_X11Y109_SLICE_X14Y109_DO5),
.O6(CLBLM_R_X11Y109_SLICE_X14Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c69c39669c3963c)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_CLUT (
.I0(CLBLM_L_X10Y108_SLICE_X12Y108_AO6),
.I1(CLBLM_R_X11Y110_SLICE_X14Y110_AO5),
.I2(CLBLM_R_X11Y109_SLICE_X15Y109_BO6),
.I3(CLBLM_R_X11Y108_SLICE_X14Y108_CO6),
.I4(CLBLM_R_X11Y110_SLICE_X15Y110_CO6),
.I5(CLBLM_R_X11Y109_SLICE_X15Y109_AO6),
.O5(CLBLM_R_X11Y109_SLICE_X14Y109_CO5),
.O6(CLBLM_R_X11Y109_SLICE_X14Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0c8e0c8e000000)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_L_X10Y109_SLICE_X13Y109_AO5),
.I2(CLBLM_R_X11Y106_SLICE_X14Y106_AO6),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_L_X10Y108_SLICE_X13Y108_CO6),
.O5(CLBLM_R_X11Y109_SLICE_X14Y109_BO5),
.O6(CLBLM_R_X11Y109_SLICE_X14Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h96f0a53c5af0963c)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y109_SLICE_X13Y109_AO5),
.I2(CLBLM_L_X10Y109_SLICE_X13Y109_BO6),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(CLBLM_R_X11Y106_SLICE_X14Y106_AO6),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_R_X11Y109_SLICE_X14Y109_AO5),
.O6(CLBLM_R_X11Y109_SLICE_X14Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y109_SLICE_X15Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y109_SLICE_X15Y109_DO5),
.O6(CLBLM_R_X11Y109_SLICE_X15Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y109_SLICE_X15Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y109_SLICE_X15Y109_CO5),
.O6(CLBLM_R_X11Y109_SLICE_X15Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe80ec80c8808080)
  ) CLBLM_R_X11Y109_SLICE_X15Y109_BLUT (
.I0(CLBLM_R_X11Y107_SLICE_X15Y107_DO6),
.I1(CLBLM_R_X11Y108_SLICE_X15Y108_DO6),
.I2(CLBLM_R_X11Y108_SLICE_X15Y108_CO6),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_R_X11Y109_SLICE_X15Y109_BO5),
.O6(CLBLM_R_X11Y109_SLICE_X15Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc96693cc36666ccc)
  ) CLBLM_R_X11Y109_SLICE_X15Y109_ALUT (
.I0(CLBLM_R_X11Y107_SLICE_X15Y107_DO6),
.I1(CLBLM_R_X11Y108_SLICE_X15Y108_DO6),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(CLBLM_R_X11Y108_SLICE_X15Y108_CO6),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_R_X11Y109_SLICE_X15Y109_AO5),
.O6(CLBLM_R_X11Y109_SLICE_X15Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2c48684040c0c0c0)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_DLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(RIOB33_X105Y111_IOB_X1Y111_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLM_L_X12Y110_SLICE_X17Y110_AO6),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_R_X11Y110_SLICE_X14Y110_DO5),
.O6(CLBLM_R_X11Y110_SLICE_X14Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeeaa88088008800)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_CLUT (
.I0(CLBLM_L_X12Y110_SLICE_X17Y110_BO6),
.I1(CLBLM_R_X11Y110_SLICE_X15Y110_CO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(CLBLM_R_X11Y109_SLICE_X15Y109_BO6),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(RIOB33_X105Y107_IOB_X1Y108_I),
.O5(CLBLM_R_X11Y110_SLICE_X14Y110_CO5),
.O6(CLBLM_R_X11Y110_SLICE_X14Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h993c963c96cc66cc)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(CLBLM_L_X12Y110_SLICE_X17Y110_BO6),
.I2(CLBLM_R_X11Y110_SLICE_X15Y110_CO6),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_R_X11Y109_SLICE_X15Y109_BO6),
.O5(CLBLM_R_X11Y110_SLICE_X14Y110_BO5),
.O6(CLBLM_R_X11Y110_SLICE_X14Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc33c0ff0cccc0000)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y107_IOB_X1Y108_I),
.I2(CLBLM_R_X11Y110_SLICE_X15Y110_CO6),
.I3(CLBLM_R_X11Y109_SLICE_X15Y109_BO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y110_SLICE_X14Y110_AO5),
.O6(CLBLM_R_X11Y110_SLICE_X14Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h505aaa000aaa0000)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_DLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(1'b1),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(CLBLM_L_X12Y110_SLICE_X17Y110_AO6),
.O5(CLBLM_R_X11Y110_SLICE_X15Y110_DO5),
.O6(CLBLM_R_X11Y110_SLICE_X15Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a95956a956a956a)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_CLUT (
.I0(CLBLM_R_X11Y108_SLICE_X15Y108_BO6),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_L_X12Y110_SLICE_X16Y110_DO6),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_R_X11Y110_SLICE_X15Y110_CO5),
.O6(CLBLM_R_X11Y110_SLICE_X15Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4488a200aa00aa00)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_BLUT (
.I0(RIOB33_X105Y111_IOB_X1Y111_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y109_IOB_X1Y110_I),
.O5(CLBLM_R_X11Y110_SLICE_X15Y110_BO5),
.O6(CLBLM_R_X11Y110_SLICE_X15Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3fc03fc05a5aaaaa)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_ALUT (
.I0(CLBLM_L_X12Y110_SLICE_X16Y110_DO6),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(CLBLM_R_X11Y110_SLICE_X15Y110_BO6),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y110_SLICE_X15Y110_AO5),
.O6(CLBLM_R_X11Y110_SLICE_X15Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfce8e8c0a000a000)
  ) CLBLM_R_X11Y111_SLICE_X14Y111_DLUT (
.I0(CLBLM_L_X12Y110_SLICE_X16Y110_AO6),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(CLBLM_R_X11Y111_SLICE_X15Y111_AO6),
.I3(CLBLM_R_X11Y110_SLICE_X14Y110_CO6),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(RIOB33_X105Y107_IOB_X1Y108_I),
.O5(CLBLM_R_X11Y111_SLICE_X14Y111_DO5),
.O6(CLBLM_R_X11Y111_SLICE_X14Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h11373f7f153f7fff)
  ) CLBLM_R_X11Y111_SLICE_X14Y111_CLUT (
.I0(CLBLM_R_X11Y110_SLICE_X14Y110_AO6),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(CLBLM_L_X10Y107_SLICE_X13Y107_DO6),
.I4(CLBLM_R_X11Y110_SLICE_X14Y110_BO6),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLM_R_X11Y111_SLICE_X14Y111_CO5),
.O6(CLBLM_R_X11Y111_SLICE_X14Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h56a5a9a56a559555)
  ) CLBLM_R_X11Y111_SLICE_X14Y111_BLUT (
.I0(CLBLM_R_X11Y110_SLICE_X14Y110_BO6),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(CLBLM_R_X11Y110_SLICE_X14Y110_AO6),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(CLBLM_L_X10Y107_SLICE_X13Y107_DO6),
.O5(CLBLM_R_X11Y111_SLICE_X14Y111_BO5),
.O6(CLBLM_R_X11Y111_SLICE_X14Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1e3c78f0993366cc)
  ) CLBLM_R_X11Y111_SLICE_X14Y111_ALUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(CLBLM_R_X11Y110_SLICE_X14Y110_CO6),
.I2(CLBLM_R_X11Y111_SLICE_X15Y111_AO6),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(CLBLM_L_X12Y110_SLICE_X16Y110_AO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y111_SLICE_X14Y111_AO5),
.O6(CLBLM_R_X11Y111_SLICE_X14Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y111_SLICE_X15Y111_DO5),
.O6(CLBLM_R_X11Y111_SLICE_X15Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y111_SLICE_X15Y111_CO5),
.O6(CLBLM_R_X11Y111_SLICE_X15Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y111_SLICE_X15Y111_BO5),
.O6(CLBLM_R_X11Y111_SLICE_X15Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999966696669666)
  ) CLBLM_R_X11Y111_SLICE_X15Y111_ALUT (
.I0(CLBLM_R_X11Y110_SLICE_X15Y110_DO6),
.I1(CLBLM_L_X12Y110_SLICE_X16Y110_CO6),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLM_R_X11Y111_SLICE_X15Y111_AO5),
.O6(CLBLM_R_X11Y111_SLICE_X15Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y101_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y101_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y102_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y102_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y103_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y103_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y104_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y104_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y105_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y105_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y106_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y106_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y107_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y107_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y108_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y108_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y109_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y109_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y110_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y110_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y111_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y111_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y112_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y112_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y113_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y113_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y114_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y114_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y115_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y115_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y116_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y116_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y117_IOB_X0Y117_IBUF (
.I(LIOB33_X0Y117_IOB_X0Y117_IPAD),
.O(LIOB33_X0Y117_IOB_X0Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y118_OBUF (
.I(CLBLL_L_X2Y111_SLICE_X0Y111_AO5),
.O(LIOB33_X0Y117_IOB_X0Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUF (
.I(CLBLL_L_X2Y110_SLICE_X0Y110_AO5),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUF (
.I(CLBLL_L_X2Y110_SLICE_X0Y110_CO5),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUF (
.I(CLBLL_L_X2Y109_SLICE_X0Y109_AO5),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUF (
.I(CLBLL_L_X2Y110_SLICE_X0Y110_BO6),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUF (
.I(CLBLL_L_X2Y109_SLICE_X0Y109_DO6),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(CLBLL_L_X2Y110_SLICE_X0Y110_BO5),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y125_OBUF (
.I(CLBLL_L_X2Y109_SLICE_X0Y109_AO6),
.O(LIOB33_X0Y125_IOB_X0Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y126_OBUF (
.I(CLBLL_L_X2Y108_SLICE_X1Y108_BO6),
.O(LIOB33_X0Y125_IOB_X0Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y127_OBUF (
.I(CLBLL_L_X2Y111_SLICE_X0Y111_BO5),
.O(LIOB33_X0Y127_IOB_X0Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y128_OBUF (
.I(CLBLL_L_X2Y111_SLICE_X1Y111_AO6),
.O(LIOB33_X0Y127_IOB_X0Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y129_OBUF (
.I(CLBLL_L_X2Y111_SLICE_X1Y111_BO6),
.O(LIOB33_X0Y129_IOB_X0Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y130_OBUF (
.I(CLBLL_L_X2Y111_SLICE_X0Y111_BO6),
.O(LIOB33_X0Y129_IOB_X0Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y131_OBUF (
.I(CLBLM_R_X3Y111_SLICE_X2Y111_AO5),
.O(LIOB33_X0Y131_IOB_X0Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y132_OBUF (
.I(CLBLL_L_X2Y111_SLICE_X1Y111_AO5),
.O(LIOB33_X0Y131_IOB_X0Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y133_OBUF (
.I(CLBLM_R_X5Y110_SLICE_X6Y110_AO6),
.O(LIOB33_X0Y133_IOB_X0Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y134_OBUF (
.I(1'b0),
.O(LIOB33_X0Y133_IOB_X0Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y135_OBUF (
.I(CLBLM_R_X3Y112_SLICE_X3Y112_BO5),
.O(LIOB33_X0Y135_IOB_X0Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUF (
.I(CLBLM_R_X3Y112_SLICE_X3Y112_CO6),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUF (
.I(CLBLL_L_X4Y114_SLICE_X4Y114_AO6),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUF (
.I(CLBLL_L_X4Y114_SLICE_X4Y114_BO6),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUF (
.I(CLBLL_L_X4Y114_SLICE_X5Y114_AO5),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUF (
.I(CLBLL_L_X4Y114_SLICE_X5Y114_AO6),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y141_OBUF (
.I(CLBLM_R_X5Y116_SLICE_X6Y116_DO6),
.O(LIOB33_X0Y141_IOB_X0Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y142_OBUF (
.I(CLBLM_R_X5Y116_SLICE_X6Y116_BO6),
.O(LIOB33_X0Y141_IOB_X0Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y143_IOB_X0Y143_OBUF (
.I(CLBLL_L_X4Y115_SLICE_X5Y115_AO6),
.O(LIOB33_X0Y143_IOB_X0Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y145_OBUF (
.I(CLBLM_R_X5Y115_SLICE_X7Y115_CO6),
.O(LIOB33_X0Y145_IOB_X0Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y146_OBUF (
.I(CLBLM_R_X5Y113_SLICE_X6Y113_AO6),
.O(LIOB33_X0Y145_IOB_X0Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y147_OBUF (
.I(CLBLM_R_X5Y113_SLICE_X6Y113_AO5),
.O(LIOB33_X0Y147_IOB_X0Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y148_OBUF (
.I(CLBLM_R_X5Y113_SLICE_X7Y113_CO6),
.O(LIOB33_X0Y147_IOB_X0Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y100_IOB_X0Y100_IBUF (
.I(LIOB33_SING_X0Y100_IOB_X0Y100_IPAD),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_OBUF (
.I(CLBLM_R_X5Y113_SLICE_X6Y113_CO6),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y101_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y102_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y103_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y104_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y105_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y105_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y106_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y107_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y108_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y109_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y110_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y111_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y112_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y113_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y100_IOB_X1Y100_IBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_IPAD),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_I)
  );
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A = CLBLL_L_X2Y105_SLICE_X0Y105_AO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B = CLBLL_L_X2Y105_SLICE_X0Y105_BO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C = CLBLL_L_X2Y105_SLICE_X0Y105_CO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D = CLBLL_L_X2Y105_SLICE_X0Y105_DO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_AMUX = CLBLL_L_X2Y105_SLICE_X0Y105_AO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A = CLBLL_L_X2Y105_SLICE_X1Y105_AO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B = CLBLL_L_X2Y105_SLICE_X1Y105_BO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C = CLBLL_L_X2Y105_SLICE_X1Y105_CO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D = CLBLL_L_X2Y105_SLICE_X1Y105_DO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_AMUX = CLBLL_L_X2Y105_SLICE_X1Y105_AO5;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A = CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B = CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C = CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D = CLBLL_L_X2Y106_SLICE_X0Y106_DO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_AMUX = CLBLL_L_X2Y106_SLICE_X0Y106_AO5;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_BMUX = CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A = CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B = CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C = CLBLL_L_X2Y106_SLICE_X1Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D = CLBLL_L_X2Y106_SLICE_X1Y106_DO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_AMUX = CLBLL_L_X2Y106_SLICE_X1Y106_AO5;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_BMUX = CLBLL_L_X2Y106_SLICE_X1Y106_BO5;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_DMUX = CLBLL_L_X2Y106_SLICE_X1Y106_DO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B = CLBLL_L_X2Y107_SLICE_X0Y107_BO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C = CLBLL_L_X2Y107_SLICE_X0Y107_CO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D = CLBLL_L_X2Y107_SLICE_X0Y107_DO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_AMUX = CLBLL_L_X2Y107_SLICE_X0Y107_AO5;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A = CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B = CLBLL_L_X2Y107_SLICE_X1Y107_BO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C = CLBLL_L_X2Y107_SLICE_X1Y107_CO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D = CLBLL_L_X2Y107_SLICE_X1Y107_DO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_AMUX = CLBLL_L_X2Y107_SLICE_X1Y107_AO5;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A = CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B = CLBLL_L_X2Y108_SLICE_X0Y108_BO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C = CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D = CLBLL_L_X2Y108_SLICE_X0Y108_DO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_AMUX = CLBLL_L_X2Y108_SLICE_X0Y108_AO5;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_BMUX = CLBLL_L_X2Y108_SLICE_X0Y108_BO5;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A = CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B = CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C = CLBLL_L_X2Y108_SLICE_X1Y108_CO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D = CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_AMUX = CLBLL_L_X2Y108_SLICE_X1Y108_AO5;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A = CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B = CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C = CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D = CLBLL_L_X2Y109_SLICE_X0Y109_DO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_AMUX = CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A = CLBLL_L_X2Y109_SLICE_X1Y109_AO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B = CLBLL_L_X2Y109_SLICE_X1Y109_BO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C = CLBLL_L_X2Y109_SLICE_X1Y109_CO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D = CLBLL_L_X2Y109_SLICE_X1Y109_DO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A = CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B = CLBLL_L_X2Y110_SLICE_X0Y110_BO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C = CLBLL_L_X2Y110_SLICE_X0Y110_CO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D = CLBLL_L_X2Y110_SLICE_X0Y110_DO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_AMUX = CLBLL_L_X2Y110_SLICE_X0Y110_AO5;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_BMUX = CLBLL_L_X2Y110_SLICE_X0Y110_BO5;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_CMUX = CLBLL_L_X2Y110_SLICE_X0Y110_CO5;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A = CLBLL_L_X2Y110_SLICE_X1Y110_AO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B = CLBLL_L_X2Y110_SLICE_X1Y110_BO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C = CLBLL_L_X2Y110_SLICE_X1Y110_CO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D = CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A = CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B = CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C = CLBLL_L_X2Y111_SLICE_X0Y111_CO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D = CLBLL_L_X2Y111_SLICE_X0Y111_DO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_AMUX = CLBLL_L_X2Y111_SLICE_X0Y111_AO5;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_BMUX = CLBLL_L_X2Y111_SLICE_X0Y111_BO5;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A = CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B = CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C = CLBLL_L_X2Y111_SLICE_X1Y111_CO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D = CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_AMUX = CLBLL_L_X2Y111_SLICE_X1Y111_AO5;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A = CLBLL_L_X4Y104_SLICE_X4Y104_AO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B = CLBLL_L_X4Y104_SLICE_X4Y104_BO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C = CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D = CLBLL_L_X4Y104_SLICE_X4Y104_DO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_AMUX = CLBLL_L_X4Y104_SLICE_X4Y104_AO5;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A = CLBLL_L_X4Y104_SLICE_X5Y104_AO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B = CLBLL_L_X4Y104_SLICE_X5Y104_BO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C = CLBLL_L_X4Y104_SLICE_X5Y104_CO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D = CLBLL_L_X4Y104_SLICE_X5Y104_DO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A = CLBLL_L_X4Y105_SLICE_X4Y105_AO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B = CLBLL_L_X4Y105_SLICE_X4Y105_BO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C = CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D = CLBLL_L_X4Y105_SLICE_X4Y105_DO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A = CLBLL_L_X4Y105_SLICE_X5Y105_AO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C = CLBLL_L_X4Y105_SLICE_X5Y105_CO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D = CLBLL_L_X4Y105_SLICE_X5Y105_DO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_AMUX = CLBLL_L_X4Y105_SLICE_X5Y105_AO5;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_BMUX = CLBLL_L_X4Y105_SLICE_X5Y105_BO5;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A = CLBLL_L_X4Y106_SLICE_X4Y106_AO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B = CLBLL_L_X4Y106_SLICE_X4Y106_BO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C = CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D = CLBLL_L_X4Y106_SLICE_X4Y106_DO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_AMUX = CLBLL_L_X4Y106_SLICE_X4Y106_AO5;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A = CLBLL_L_X4Y106_SLICE_X5Y106_AO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B = CLBLL_L_X4Y106_SLICE_X5Y106_BO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C = CLBLL_L_X4Y106_SLICE_X5Y106_CO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D = CLBLL_L_X4Y106_SLICE_X5Y106_DO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A = CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B = CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C = CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D = CLBLL_L_X4Y107_SLICE_X4Y107_DO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_AMUX = CLBLL_L_X4Y107_SLICE_X4Y107_AO5;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_BMUX = CLBLL_L_X4Y107_SLICE_X4Y107_BO5;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A = CLBLL_L_X4Y107_SLICE_X5Y107_AO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B = CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C = CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D = CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B = CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D = CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A = CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B = CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C = CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D = CLBLL_L_X4Y108_SLICE_X5Y108_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A = CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B = CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_AMUX = CLBLL_L_X4Y109_SLICE_X4Y109_AO5;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_BMUX = CLBLL_L_X4Y109_SLICE_X4Y109_BO5;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A = CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B = CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C = CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D = CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_AMUX = CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_BMUX = CLBLL_L_X4Y109_SLICE_X5Y109_BO5;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A = CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B = CLBLL_L_X4Y110_SLICE_X4Y110_BO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C = CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D = CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_AMUX = CLBLL_L_X4Y110_SLICE_X4Y110_AO5;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A = CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B = CLBLL_L_X4Y110_SLICE_X5Y110_BO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C = CLBLL_L_X4Y110_SLICE_X5Y110_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D = CLBLL_L_X4Y110_SLICE_X5Y110_DO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A = CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B = CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C = CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A = CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B = CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D = CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A = CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B = CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D = CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_AMUX = CLBLL_L_X4Y112_SLICE_X4Y112_AO5;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A = CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C = CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D = CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A = CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D = CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_AMUX = CLBLL_L_X4Y113_SLICE_X4Y113_AO5;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A = CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C = CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D = CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A = CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B = CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C = CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D = CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_AMUX = CLBLL_L_X4Y114_SLICE_X4Y114_AO5;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_BMUX = CLBLL_L_X4Y114_SLICE_X4Y114_BO5;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_CMUX = CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A = CLBLL_L_X4Y114_SLICE_X5Y114_AO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B = CLBLL_L_X4Y114_SLICE_X5Y114_BO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C = CLBLL_L_X4Y114_SLICE_X5Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D = CLBLL_L_X4Y114_SLICE_X5Y114_DO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_AMUX = CLBLL_L_X4Y114_SLICE_X5Y114_AO5;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_CMUX = CLBLL_L_X4Y114_SLICE_X5Y114_CO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A = CLBLL_L_X4Y115_SLICE_X4Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B = CLBLL_L_X4Y115_SLICE_X4Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C = CLBLL_L_X4Y115_SLICE_X4Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D = CLBLL_L_X4Y115_SLICE_X4Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A = CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B = CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C = CLBLL_L_X4Y115_SLICE_X5Y115_CO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D = CLBLL_L_X4Y115_SLICE_X5Y115_DO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_AMUX = CLBLL_L_X4Y115_SLICE_X5Y115_AO5;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_A = CLBLM_L_X8Y102_SLICE_X10Y102_AO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_B = CLBLM_L_X8Y102_SLICE_X10Y102_BO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_C = CLBLM_L_X8Y102_SLICE_X10Y102_CO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_D = CLBLM_L_X8Y102_SLICE_X10Y102_DO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_AMUX = CLBLM_L_X8Y102_SLICE_X10Y102_AO5;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_A = CLBLM_L_X8Y102_SLICE_X11Y102_AO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_B = CLBLM_L_X8Y102_SLICE_X11Y102_BO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_C = CLBLM_L_X8Y102_SLICE_X11Y102_CO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_D = CLBLM_L_X8Y102_SLICE_X11Y102_DO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_AMUX = CLBLM_L_X8Y102_SLICE_X11Y102_AO5;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A = CLBLM_L_X8Y103_SLICE_X10Y103_AO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B = CLBLM_L_X8Y103_SLICE_X10Y103_BO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C = CLBLM_L_X8Y103_SLICE_X10Y103_CO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D = CLBLM_L_X8Y103_SLICE_X10Y103_DO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_AMUX = CLBLM_L_X8Y103_SLICE_X10Y103_AO5;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A = CLBLM_L_X8Y103_SLICE_X11Y103_AO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B = CLBLM_L_X8Y103_SLICE_X11Y103_BO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C = CLBLM_L_X8Y103_SLICE_X11Y103_CO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D = CLBLM_L_X8Y103_SLICE_X11Y103_DO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A = CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B = CLBLM_L_X8Y104_SLICE_X10Y104_BO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C = CLBLM_L_X8Y104_SLICE_X10Y104_CO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D = CLBLM_L_X8Y104_SLICE_X10Y104_DO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A = CLBLM_L_X8Y104_SLICE_X11Y104_AO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B = CLBLM_L_X8Y104_SLICE_X11Y104_BO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C = CLBLM_L_X8Y104_SLICE_X11Y104_CO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D = CLBLM_L_X8Y104_SLICE_X11Y104_DO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A = CLBLM_L_X8Y105_SLICE_X10Y105_AO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B = CLBLM_L_X8Y105_SLICE_X10Y105_BO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C = CLBLM_L_X8Y105_SLICE_X10Y105_CO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D = CLBLM_L_X8Y105_SLICE_X10Y105_DO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_AMUX = CLBLM_L_X8Y105_SLICE_X10Y105_AO5;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A = CLBLM_L_X8Y105_SLICE_X11Y105_AO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B = CLBLM_L_X8Y105_SLICE_X11Y105_BO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C = CLBLM_L_X8Y105_SLICE_X11Y105_CO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D = CLBLM_L_X8Y105_SLICE_X11Y105_DO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A = CLBLM_L_X8Y106_SLICE_X10Y106_AO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B = CLBLM_L_X8Y106_SLICE_X10Y106_BO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C = CLBLM_L_X8Y106_SLICE_X10Y106_CO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D = CLBLM_L_X8Y106_SLICE_X10Y106_DO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A = CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B = CLBLM_L_X8Y106_SLICE_X11Y106_BO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C = CLBLM_L_X8Y106_SLICE_X11Y106_CO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D = CLBLM_L_X8Y106_SLICE_X11Y106_DO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_AMUX = CLBLM_L_X8Y106_SLICE_X11Y106_AO5;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A = CLBLM_L_X8Y107_SLICE_X10Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B = CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C = CLBLM_L_X8Y107_SLICE_X10Y107_CO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D = CLBLM_L_X8Y107_SLICE_X10Y107_DO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_AMUX = CLBLM_L_X8Y107_SLICE_X10Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A = CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B = CLBLM_L_X8Y107_SLICE_X11Y107_BO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C = CLBLM_L_X8Y107_SLICE_X11Y107_CO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D = CLBLM_L_X8Y107_SLICE_X11Y107_DO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_AMUX = CLBLM_L_X8Y107_SLICE_X11Y107_AO5;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A = CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B = CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C = CLBLM_L_X8Y108_SLICE_X10Y108_CO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D = CLBLM_L_X8Y108_SLICE_X10Y108_DO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_AMUX = CLBLM_L_X8Y108_SLICE_X10Y108_AO5;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A = CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B = CLBLM_L_X8Y108_SLICE_X11Y108_BO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C = CLBLM_L_X8Y108_SLICE_X11Y108_CO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D = CLBLM_L_X8Y108_SLICE_X11Y108_DO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A = CLBLM_L_X8Y109_SLICE_X10Y109_AO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B = CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C = CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D = CLBLM_L_X8Y109_SLICE_X10Y109_DO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A = CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B = CLBLM_L_X8Y109_SLICE_X11Y109_BO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C = CLBLM_L_X8Y109_SLICE_X11Y109_CO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D = CLBLM_L_X8Y109_SLICE_X11Y109_DO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_AMUX = CLBLM_L_X8Y109_SLICE_X11Y109_AO5;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A = CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_AMUX = CLBLM_L_X8Y110_SLICE_X10Y110_AO5;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_BMUX = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A = CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B = CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D = CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_AMUX = CLBLM_L_X8Y110_SLICE_X11Y110_AO5;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A = CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B = CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D = CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A = CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B = CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D = CLBLM_L_X8Y111_SLICE_X11Y111_DO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_AMUX = CLBLM_L_X8Y111_SLICE_X11Y111_AO5;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_BMUX = CLBLM_L_X8Y111_SLICE_X11Y111_BO5;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A = CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B = CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C = CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D = CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A = CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B = CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C = CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D = CLBLM_L_X8Y112_SLICE_X11Y112_DO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_AMUX = CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B = CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C = CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_AMUX = CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_BMUX = CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A = CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B = CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C = CLBLM_L_X8Y113_SLICE_X11Y113_CO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D = CLBLM_L_X8Y113_SLICE_X11Y113_DO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A = CLBLM_L_X8Y114_SLICE_X10Y114_AO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B = CLBLM_L_X8Y114_SLICE_X10Y114_BO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C = CLBLM_L_X8Y114_SLICE_X10Y114_CO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D = CLBLM_L_X8Y114_SLICE_X10Y114_DO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_AMUX = CLBLM_L_X8Y114_SLICE_X10Y114_AO5;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_BMUX = CLBLM_L_X8Y114_SLICE_X10Y114_BO5;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A = CLBLM_L_X8Y114_SLICE_X11Y114_AO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B = CLBLM_L_X8Y114_SLICE_X11Y114_BO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C = CLBLM_L_X8Y114_SLICE_X11Y114_CO6;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D = CLBLM_L_X8Y114_SLICE_X11Y114_DO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A = CLBLM_L_X10Y103_SLICE_X12Y103_AO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B = CLBLM_L_X10Y103_SLICE_X12Y103_BO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C = CLBLM_L_X10Y103_SLICE_X12Y103_CO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D = CLBLM_L_X10Y103_SLICE_X12Y103_DO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_AMUX = CLBLM_L_X10Y103_SLICE_X12Y103_AO5;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_BMUX = CLBLM_L_X10Y103_SLICE_X12Y103_BO5;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_CMUX = CLBLM_L_X10Y103_SLICE_X12Y103_CO5;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A = CLBLM_L_X10Y103_SLICE_X13Y103_AO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B = CLBLM_L_X10Y103_SLICE_X13Y103_BO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C = CLBLM_L_X10Y103_SLICE_X13Y103_CO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D = CLBLM_L_X10Y103_SLICE_X13Y103_DO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_AMUX = CLBLM_L_X10Y103_SLICE_X13Y103_AO5;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A = CLBLM_L_X10Y104_SLICE_X12Y104_AO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C = CLBLM_L_X10Y104_SLICE_X12Y104_CO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D = CLBLM_L_X10Y104_SLICE_X12Y104_DO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_DMUX = CLBLM_L_X10Y104_SLICE_X12Y104_DO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A = CLBLM_L_X10Y104_SLICE_X13Y104_AO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B = CLBLM_L_X10Y104_SLICE_X13Y104_BO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C = CLBLM_L_X10Y104_SLICE_X13Y104_CO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D = CLBLM_L_X10Y104_SLICE_X13Y104_DO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_AMUX = CLBLM_L_X10Y104_SLICE_X13Y104_AO5;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_BMUX = CLBLM_L_X10Y104_SLICE_X13Y104_BO5;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_CMUX = CLBLM_L_X10Y104_SLICE_X13Y104_CO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A = CLBLM_L_X10Y105_SLICE_X12Y105_AO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B = CLBLM_L_X10Y105_SLICE_X12Y105_BO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C = CLBLM_L_X10Y105_SLICE_X12Y105_CO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D = CLBLM_L_X10Y105_SLICE_X12Y105_DO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_CMUX = CLBLM_L_X10Y105_SLICE_X12Y105_CO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_DMUX = CLBLM_L_X10Y105_SLICE_X12Y105_DO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A = CLBLM_L_X10Y105_SLICE_X13Y105_AO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B = CLBLM_L_X10Y105_SLICE_X13Y105_BO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C = CLBLM_L_X10Y105_SLICE_X13Y105_CO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D = CLBLM_L_X10Y105_SLICE_X13Y105_DO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A = CLBLM_L_X10Y106_SLICE_X12Y106_AO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C = CLBLM_L_X10Y106_SLICE_X12Y106_CO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D = CLBLM_L_X10Y106_SLICE_X12Y106_DO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A = CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B = CLBLM_L_X10Y106_SLICE_X13Y106_BO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C = CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D = CLBLM_L_X10Y106_SLICE_X13Y106_DO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A = CLBLM_L_X10Y107_SLICE_X12Y107_AO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B = CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C = CLBLM_L_X10Y107_SLICE_X12Y107_CO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D = CLBLM_L_X10Y107_SLICE_X12Y107_DO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A = CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B = CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C = CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D = CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_AMUX = CLBLM_L_X10Y107_SLICE_X13Y107_AO5;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A = CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B = CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C = CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D = CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_AMUX = CLBLM_L_X10Y108_SLICE_X12Y108_AO5;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A = CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B = CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C = CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D = CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_AMUX = CLBLM_L_X10Y108_SLICE_X13Y108_AO5;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_BMUX = CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A = CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C = CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_AMUX = CLBLM_L_X10Y109_SLICE_X12Y109_AO5;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A = CLBLM_L_X10Y109_SLICE_X13Y109_AO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B = CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D = CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_AMUX = CLBLM_L_X10Y109_SLICE_X13Y109_AO5;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A = CLBLM_L_X10Y110_SLICE_X12Y110_AO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B = CLBLM_L_X10Y110_SLICE_X12Y110_BO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C = CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D = CLBLM_L_X10Y110_SLICE_X12Y110_DO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_AMUX = CLBLM_L_X10Y110_SLICE_X12Y110_AO5;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A = CLBLM_L_X10Y110_SLICE_X13Y110_AO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B = CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C = CLBLM_L_X10Y110_SLICE_X13Y110_CO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D = CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_AMUX = CLBLM_L_X10Y110_SLICE_X13Y110_AO5;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_DMUX = CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A = CLBLM_L_X10Y111_SLICE_X12Y111_AO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B = CLBLM_L_X10Y111_SLICE_X12Y111_BO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C = CLBLM_L_X10Y111_SLICE_X12Y111_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D = CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A = CLBLM_L_X10Y111_SLICE_X13Y111_AO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B = CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C = CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D = CLBLM_L_X10Y111_SLICE_X13Y111_DO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_AMUX = CLBLM_L_X10Y111_SLICE_X13Y111_AO5;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_BMUX = CLBLM_L_X10Y111_SLICE_X13Y111_BO5;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_DMUX = CLBLM_L_X10Y111_SLICE_X13Y111_DO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A = CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B = CLBLM_L_X10Y112_SLICE_X12Y112_BO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C = CLBLM_L_X10Y112_SLICE_X12Y112_CO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D = CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_AMUX = CLBLM_L_X10Y112_SLICE_X12Y112_AO5;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A = CLBLM_L_X10Y112_SLICE_X13Y112_AO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B = CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C = CLBLM_L_X10Y112_SLICE_X13Y112_CO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D = CLBLM_L_X10Y112_SLICE_X13Y112_DO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_AMUX = CLBLM_L_X10Y112_SLICE_X13Y112_AO5;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A = CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B = CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C = CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D = CLBLM_L_X10Y113_SLICE_X12Y113_DO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_AMUX = CLBLM_L_X10Y113_SLICE_X12Y113_AO5;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A = CLBLM_L_X10Y113_SLICE_X13Y113_AO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B = CLBLM_L_X10Y113_SLICE_X13Y113_BO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C = CLBLM_L_X10Y113_SLICE_X13Y113_CO6;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D = CLBLM_L_X10Y113_SLICE_X13Y113_DO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A = CLBLM_L_X12Y107_SLICE_X16Y107_AO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B = CLBLM_L_X12Y107_SLICE_X16Y107_BO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C = CLBLM_L_X12Y107_SLICE_X16Y107_CO6;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D = CLBLM_L_X12Y107_SLICE_X16Y107_DO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A = CLBLM_L_X12Y107_SLICE_X17Y107_AO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B = CLBLM_L_X12Y107_SLICE_X17Y107_BO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C = CLBLM_L_X12Y107_SLICE_X17Y107_CO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D = CLBLM_L_X12Y107_SLICE_X17Y107_DO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A = CLBLM_L_X12Y108_SLICE_X16Y108_AO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B = CLBLM_L_X12Y108_SLICE_X16Y108_BO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C = CLBLM_L_X12Y108_SLICE_X16Y108_CO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D = CLBLM_L_X12Y108_SLICE_X16Y108_DO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A = CLBLM_L_X12Y108_SLICE_X17Y108_AO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B = CLBLM_L_X12Y108_SLICE_X17Y108_BO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C = CLBLM_L_X12Y108_SLICE_X17Y108_CO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D = CLBLM_L_X12Y108_SLICE_X17Y108_DO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A = CLBLM_L_X12Y109_SLICE_X16Y109_AO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B = CLBLM_L_X12Y109_SLICE_X16Y109_BO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C = CLBLM_L_X12Y109_SLICE_X16Y109_CO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D = CLBLM_L_X12Y109_SLICE_X16Y109_DO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A = CLBLM_L_X12Y109_SLICE_X17Y109_AO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B = CLBLM_L_X12Y109_SLICE_X17Y109_BO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C = CLBLM_L_X12Y109_SLICE_X17Y109_CO6;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D = CLBLM_L_X12Y109_SLICE_X17Y109_DO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A = CLBLM_L_X12Y110_SLICE_X16Y110_AO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B = CLBLM_L_X12Y110_SLICE_X16Y110_BO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C = CLBLM_L_X12Y110_SLICE_X16Y110_CO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D = CLBLM_L_X12Y110_SLICE_X16Y110_DO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A = CLBLM_L_X12Y110_SLICE_X17Y110_AO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B = CLBLM_L_X12Y110_SLICE_X17Y110_BO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C = CLBLM_L_X12Y110_SLICE_X17Y110_CO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D = CLBLM_L_X12Y110_SLICE_X17Y110_DO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_CMUX = CLBLM_L_X12Y110_SLICE_X17Y110_CO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A = CLBLM_R_X3Y103_SLICE_X2Y103_AO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B = CLBLM_R_X3Y103_SLICE_X2Y103_BO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C = CLBLM_R_X3Y103_SLICE_X2Y103_CO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D = CLBLM_R_X3Y103_SLICE_X2Y103_DO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A = CLBLM_R_X3Y103_SLICE_X3Y103_AO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B = CLBLM_R_X3Y103_SLICE_X3Y103_BO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C = CLBLM_R_X3Y103_SLICE_X3Y103_CO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D = CLBLM_R_X3Y103_SLICE_X3Y103_DO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A = CLBLM_R_X3Y104_SLICE_X2Y104_AO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B = CLBLM_R_X3Y104_SLICE_X2Y104_BO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C = CLBLM_R_X3Y104_SLICE_X2Y104_CO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D = CLBLM_R_X3Y104_SLICE_X2Y104_DO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_AMUX = CLBLM_R_X3Y104_SLICE_X2Y104_AO5;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_BMUX = CLBLM_R_X3Y104_SLICE_X2Y104_BO5;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_CMUX = CLBLM_R_X3Y104_SLICE_X2Y104_CO5;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A = CLBLM_R_X3Y104_SLICE_X3Y104_AO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B = CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C = CLBLM_R_X3Y104_SLICE_X3Y104_CO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D = CLBLM_R_X3Y104_SLICE_X3Y104_DO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_AMUX = CLBLM_R_X3Y104_SLICE_X3Y104_AO5;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_BMUX = CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A = CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B = CLBLM_R_X3Y105_SLICE_X2Y105_BO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C = CLBLM_R_X3Y105_SLICE_X2Y105_CO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D = CLBLM_R_X3Y105_SLICE_X2Y105_DO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_AMUX = CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A = CLBLM_R_X3Y105_SLICE_X3Y105_AO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B = CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C = CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D = CLBLM_R_X3Y105_SLICE_X3Y105_DO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_AMUX = CLBLM_R_X3Y105_SLICE_X3Y105_AO5;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A = CLBLM_R_X3Y106_SLICE_X2Y106_AO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B = CLBLM_R_X3Y106_SLICE_X2Y106_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C = CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D = CLBLM_R_X3Y106_SLICE_X2Y106_DO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A = CLBLM_R_X3Y106_SLICE_X3Y106_AO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B = CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C = CLBLM_R_X3Y106_SLICE_X3Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D = CLBLM_R_X3Y106_SLICE_X3Y106_DO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_AMUX = CLBLM_R_X3Y106_SLICE_X3Y106_AO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A = CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B = CLBLM_R_X3Y107_SLICE_X2Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C = CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D = CLBLM_R_X3Y107_SLICE_X2Y107_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A = CLBLM_R_X3Y107_SLICE_X3Y107_AO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B = CLBLM_R_X3Y107_SLICE_X3Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C = CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D = CLBLM_R_X3Y107_SLICE_X3Y107_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_AMUX = CLBLM_R_X3Y107_SLICE_X3Y107_AO5;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_BMUX = CLBLM_R_X3Y107_SLICE_X3Y107_BO5;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A = CLBLM_R_X3Y108_SLICE_X2Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B = CLBLM_R_X3Y108_SLICE_X2Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C = CLBLM_R_X3Y108_SLICE_X2Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D = CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_AMUX = CLBLM_R_X3Y108_SLICE_X2Y108_AO5;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_CMUX = CLBLM_R_X3Y108_SLICE_X2Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A = CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B = CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C = CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A = CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B = CLBLM_R_X3Y109_SLICE_X2Y109_BO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D = CLBLM_R_X3Y109_SLICE_X2Y109_DO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_AMUX = CLBLM_R_X3Y109_SLICE_X2Y109_AO5;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A = CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B = CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C = CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D = CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_AMUX = CLBLM_R_X3Y109_SLICE_X3Y109_AO5;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_BMUX = CLBLM_R_X3Y109_SLICE_X3Y109_BO5;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_CMUX = CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A = CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C = CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_AMUX = CLBLM_R_X3Y110_SLICE_X2Y110_AO5;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_BMUX = CLBLM_R_X3Y110_SLICE_X2Y110_BO5;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B = CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C = CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_AMUX = CLBLM_R_X3Y110_SLICE_X3Y110_AO5;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A = CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B = CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D = CLBLM_R_X3Y111_SLICE_X2Y111_DO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_AMUX = CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A = CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B = CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C = CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_AMUX = CLBLM_R_X3Y111_SLICE_X3Y111_AO5;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A = CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B = CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C = CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D = CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A = CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C = CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D = CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_AMUX = CLBLM_R_X3Y112_SLICE_X3Y112_AO5;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_BMUX = CLBLM_R_X3Y112_SLICE_X3Y112_BO5;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_A = CLBLM_R_X5Y101_SLICE_X6Y101_AO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_B = CLBLM_R_X5Y101_SLICE_X6Y101_BO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_C = CLBLM_R_X5Y101_SLICE_X6Y101_CO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_D = CLBLM_R_X5Y101_SLICE_X6Y101_DO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_AMUX = CLBLM_R_X5Y101_SLICE_X6Y101_AO5;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_A = CLBLM_R_X5Y101_SLICE_X7Y101_AO6;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_B = CLBLM_R_X5Y101_SLICE_X7Y101_BO6;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_C = CLBLM_R_X5Y101_SLICE_X7Y101_CO6;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_D = CLBLM_R_X5Y101_SLICE_X7Y101_DO6;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_AMUX = CLBLM_R_X5Y101_SLICE_X7Y101_AO5;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_A = CLBLM_R_X5Y102_SLICE_X6Y102_AO6;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_B = CLBLM_R_X5Y102_SLICE_X6Y102_BO6;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_C = CLBLM_R_X5Y102_SLICE_X6Y102_CO6;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_D = CLBLM_R_X5Y102_SLICE_X6Y102_DO6;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_AMUX = CLBLM_R_X5Y102_SLICE_X6Y102_AO5;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_A = CLBLM_R_X5Y102_SLICE_X7Y102_AO6;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_B = CLBLM_R_X5Y102_SLICE_X7Y102_BO6;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_C = CLBLM_R_X5Y102_SLICE_X7Y102_CO6;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_D = CLBLM_R_X5Y102_SLICE_X7Y102_DO6;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_AMUX = CLBLM_R_X5Y102_SLICE_X7Y102_AO5;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_A = CLBLM_R_X5Y103_SLICE_X6Y103_AO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_B = CLBLM_R_X5Y103_SLICE_X6Y103_BO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_C = CLBLM_R_X5Y103_SLICE_X6Y103_CO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_D = CLBLM_R_X5Y103_SLICE_X6Y103_DO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_AMUX = CLBLM_R_X5Y103_SLICE_X6Y103_AO5;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_A = CLBLM_R_X5Y103_SLICE_X7Y103_AO6;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_B = CLBLM_R_X5Y103_SLICE_X7Y103_BO6;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_C = CLBLM_R_X5Y103_SLICE_X7Y103_CO6;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_D = CLBLM_R_X5Y103_SLICE_X7Y103_DO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A = CLBLM_R_X5Y104_SLICE_X6Y104_AO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B = CLBLM_R_X5Y104_SLICE_X6Y104_BO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C = CLBLM_R_X5Y104_SLICE_X6Y104_CO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D = CLBLM_R_X5Y104_SLICE_X6Y104_DO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A = CLBLM_R_X5Y104_SLICE_X7Y104_AO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B = CLBLM_R_X5Y104_SLICE_X7Y104_BO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C = CLBLM_R_X5Y104_SLICE_X7Y104_CO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D = CLBLM_R_X5Y104_SLICE_X7Y104_DO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A = CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B = CLBLM_R_X5Y105_SLICE_X6Y105_BO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C = CLBLM_R_X5Y105_SLICE_X6Y105_CO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D = CLBLM_R_X5Y105_SLICE_X6Y105_DO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_AMUX = CLBLM_R_X5Y105_SLICE_X6Y105_AO5;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_DMUX = CLBLM_R_X5Y105_SLICE_X6Y105_DO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A = CLBLM_R_X5Y105_SLICE_X7Y105_AO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B = CLBLM_R_X5Y105_SLICE_X7Y105_BO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C = CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D = CLBLM_R_X5Y105_SLICE_X7Y105_DO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A = CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B = CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C = CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D = CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_AMUX = CLBLM_R_X5Y106_SLICE_X6Y106_AO5;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A = CLBLM_R_X5Y106_SLICE_X7Y106_AO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B = CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C = CLBLM_R_X5Y106_SLICE_X7Y106_CO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D = CLBLM_R_X5Y106_SLICE_X7Y106_DO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A = CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C = CLBLM_R_X5Y107_SLICE_X6Y107_CO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D = CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_AMUX = CLBLM_R_X5Y107_SLICE_X6Y107_AO5;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A = CLBLM_R_X5Y107_SLICE_X7Y107_AO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C = CLBLM_R_X5Y107_SLICE_X7Y107_CO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D = CLBLM_R_X5Y107_SLICE_X7Y107_DO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A = CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B = CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C = CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D = CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A = CLBLM_R_X5Y108_SLICE_X7Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B = CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C = CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D = CLBLM_R_X5Y108_SLICE_X7Y108_DO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A = CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B = CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C = CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D = CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A = CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B = CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C = CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D = CLBLM_R_X5Y109_SLICE_X7Y109_DO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_AMUX = CLBLM_R_X5Y109_SLICE_X7Y109_AO5;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B = CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D = CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A = CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B = CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C = CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D = CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B = CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C = CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_AMUX = CLBLM_R_X5Y111_SLICE_X6Y111_AO5;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A = CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B = CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C = CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A = CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B = CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C = CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D = CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_AMUX = CLBLM_R_X5Y112_SLICE_X6Y112_AO5;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A = CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B = CLBLM_R_X5Y112_SLICE_X7Y112_BO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C = CLBLM_R_X5Y112_SLICE_X7Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D = CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B = CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D = CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_AMUX = CLBLM_R_X5Y113_SLICE_X6Y113_AO5;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A = CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B = CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C = CLBLM_R_X5Y113_SLICE_X7Y113_CO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D = CLBLM_R_X5Y113_SLICE_X7Y113_DO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_AMUX = CLBLM_R_X5Y113_SLICE_X7Y113_AO5;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_BMUX = CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A = CLBLM_R_X5Y114_SLICE_X6Y114_AO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B = CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C = CLBLM_R_X5Y114_SLICE_X6Y114_CO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D = CLBLM_R_X5Y114_SLICE_X6Y114_DO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_AMUX = CLBLM_R_X5Y114_SLICE_X6Y114_AO5;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A = CLBLM_R_X5Y114_SLICE_X7Y114_AO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B = CLBLM_R_X5Y114_SLICE_X7Y114_BO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C = CLBLM_R_X5Y114_SLICE_X7Y114_CO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D = CLBLM_R_X5Y114_SLICE_X7Y114_DO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_AMUX = CLBLM_R_X5Y114_SLICE_X7Y114_AO5;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A = CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B = CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C = CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D = CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_AMUX = CLBLM_R_X5Y115_SLICE_X6Y115_AO5;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A = CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B = CLBLM_R_X5Y115_SLICE_X7Y115_BO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D = CLBLM_R_X5Y115_SLICE_X7Y115_DO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_AMUX = CLBLM_R_X5Y115_SLICE_X7Y115_AO5;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A = CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B = CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C = CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_AMUX = CLBLM_R_X5Y116_SLICE_X6Y116_AO5;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A = CLBLM_R_X5Y116_SLICE_X7Y116_AO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B = CLBLM_R_X5Y116_SLICE_X7Y116_BO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C = CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_A = CLBLM_R_X7Y102_SLICE_X8Y102_AO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_B = CLBLM_R_X7Y102_SLICE_X8Y102_BO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_C = CLBLM_R_X7Y102_SLICE_X8Y102_CO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_D = CLBLM_R_X7Y102_SLICE_X8Y102_DO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_AMUX = CLBLM_R_X7Y102_SLICE_X8Y102_AO5;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_BMUX = CLBLM_R_X7Y102_SLICE_X8Y102_BO5;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_CMUX = CLBLM_R_X7Y102_SLICE_X8Y102_CO5;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_A = CLBLM_R_X7Y102_SLICE_X9Y102_AO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_B = CLBLM_R_X7Y102_SLICE_X9Y102_BO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_C = CLBLM_R_X7Y102_SLICE_X9Y102_CO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_D = CLBLM_R_X7Y102_SLICE_X9Y102_DO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_AMUX = CLBLM_R_X7Y102_SLICE_X9Y102_AO5;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_CMUX = CLBLM_R_X7Y102_SLICE_X9Y102_CO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A = CLBLM_R_X7Y103_SLICE_X8Y103_AO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B = CLBLM_R_X7Y103_SLICE_X8Y103_BO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C = CLBLM_R_X7Y103_SLICE_X8Y103_CO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D = CLBLM_R_X7Y103_SLICE_X8Y103_DO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A = CLBLM_R_X7Y103_SLICE_X9Y103_AO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B = CLBLM_R_X7Y103_SLICE_X9Y103_BO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C = CLBLM_R_X7Y103_SLICE_X9Y103_CO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D = CLBLM_R_X7Y103_SLICE_X9Y103_DO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A = CLBLM_R_X7Y104_SLICE_X8Y104_AO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B = CLBLM_R_X7Y104_SLICE_X8Y104_BO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C = CLBLM_R_X7Y104_SLICE_X8Y104_CO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D = CLBLM_R_X7Y104_SLICE_X8Y104_DO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_AMUX = CLBLM_R_X7Y104_SLICE_X8Y104_AO5;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_BMUX = CLBLM_R_X7Y104_SLICE_X8Y104_BO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A = CLBLM_R_X7Y104_SLICE_X9Y104_AO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B = CLBLM_R_X7Y104_SLICE_X9Y104_BO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C = CLBLM_R_X7Y104_SLICE_X9Y104_CO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D = CLBLM_R_X7Y104_SLICE_X9Y104_DO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A = CLBLM_R_X7Y105_SLICE_X8Y105_AO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B = CLBLM_R_X7Y105_SLICE_X8Y105_BO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C = CLBLM_R_X7Y105_SLICE_X8Y105_CO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D = CLBLM_R_X7Y105_SLICE_X8Y105_DO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_AMUX = CLBLM_R_X7Y105_SLICE_X8Y105_AO5;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A = CLBLM_R_X7Y105_SLICE_X9Y105_AO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B = CLBLM_R_X7Y105_SLICE_X9Y105_BO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C = CLBLM_R_X7Y105_SLICE_X9Y105_CO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D = CLBLM_R_X7Y105_SLICE_X9Y105_DO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A = CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B = CLBLM_R_X7Y106_SLICE_X8Y106_BO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C = CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D = CLBLM_R_X7Y106_SLICE_X8Y106_DO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_AMUX = CLBLM_R_X7Y106_SLICE_X8Y106_AO5;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A = CLBLM_R_X7Y106_SLICE_X9Y106_AO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B = CLBLM_R_X7Y106_SLICE_X9Y106_BO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C = CLBLM_R_X7Y106_SLICE_X9Y106_CO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D = CLBLM_R_X7Y106_SLICE_X9Y106_DO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A = CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B = CLBLM_R_X7Y107_SLICE_X8Y107_BO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C = CLBLM_R_X7Y107_SLICE_X8Y107_CO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D = CLBLM_R_X7Y107_SLICE_X8Y107_DO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_AMUX = CLBLM_R_X7Y107_SLICE_X8Y107_AO5;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A = CLBLM_R_X7Y107_SLICE_X9Y107_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B = CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C = CLBLM_R_X7Y107_SLICE_X9Y107_CO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D = CLBLM_R_X7Y107_SLICE_X9Y107_DO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_AMUX = CLBLM_R_X7Y107_SLICE_X9Y107_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_BMUX = CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B = CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C = CLBLM_R_X7Y108_SLICE_X8Y108_CO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D = CLBLM_R_X7Y108_SLICE_X8Y108_DO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A = CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B = CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C = CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D = CLBLM_R_X7Y108_SLICE_X9Y108_DO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_AMUX = CLBLM_R_X7Y108_SLICE_X9Y108_AO5;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A = CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B = CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C = CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D = CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_AMUX = CLBLM_R_X7Y109_SLICE_X8Y109_AO5;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_BMUX = CLBLM_R_X7Y109_SLICE_X8Y109_BO5;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A = CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B = CLBLM_R_X7Y109_SLICE_X9Y109_BO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C = CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D = CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A = CLBLM_R_X7Y110_SLICE_X8Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B = CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D = CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_AMUX = CLBLM_R_X7Y110_SLICE_X8Y110_AO5;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A = CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B = CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C = CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D = CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_AMUX = CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A = CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C = CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_AMUX = CLBLM_R_X7Y111_SLICE_X8Y111_AO5;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B = CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C = CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D = CLBLM_R_X7Y111_SLICE_X9Y111_DO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_AMUX = CLBLM_R_X7Y111_SLICE_X9Y111_AO5;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B = CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C = CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A = CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A = CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C = CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_AMUX = CLBLM_R_X7Y113_SLICE_X8Y113_AO5;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A = CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B = CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_AMUX = CLBLM_R_X7Y113_SLICE_X9Y113_AO5;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_BMUX = CLBLM_R_X7Y113_SLICE_X9Y113_BO5;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A = CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B = CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C = CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D = CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A = CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B = CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C = CLBLM_R_X7Y114_SLICE_X9Y114_CO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D = CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_AMUX = CLBLM_R_X7Y114_SLICE_X9Y114_AO5;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_CMUX = CLBLM_R_X7Y114_SLICE_X9Y114_CO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A = CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B = CLBLM_R_X7Y115_SLICE_X8Y115_BO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C = CLBLM_R_X7Y115_SLICE_X8Y115_CO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D = CLBLM_R_X7Y115_SLICE_X8Y115_DO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_AMUX = CLBLM_R_X7Y115_SLICE_X8Y115_AO5;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_BMUX = CLBLM_R_X7Y115_SLICE_X8Y115_BO5;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_CMUX = CLBLM_R_X7Y115_SLICE_X8Y115_CO5;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A = CLBLM_R_X7Y115_SLICE_X9Y115_AO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B = CLBLM_R_X7Y115_SLICE_X9Y115_BO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C = CLBLM_R_X7Y115_SLICE_X9Y115_CO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D = CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_A = CLBLM_R_X11Y104_SLICE_X14Y104_AO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_B = CLBLM_R_X11Y104_SLICE_X14Y104_BO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_C = CLBLM_R_X11Y104_SLICE_X14Y104_CO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_D = CLBLM_R_X11Y104_SLICE_X14Y104_DO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_AMUX = CLBLM_R_X11Y104_SLICE_X14Y104_AO5;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_A = CLBLM_R_X11Y104_SLICE_X15Y104_AO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_B = CLBLM_R_X11Y104_SLICE_X15Y104_BO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_C = CLBLM_R_X11Y104_SLICE_X15Y104_CO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_D = CLBLM_R_X11Y104_SLICE_X15Y104_DO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A = CLBLM_R_X11Y105_SLICE_X14Y105_AO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B = CLBLM_R_X11Y105_SLICE_X14Y105_BO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C = CLBLM_R_X11Y105_SLICE_X14Y105_CO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D = CLBLM_R_X11Y105_SLICE_X14Y105_DO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_AMUX = CLBLM_R_X11Y105_SLICE_X14Y105_AO5;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A = CLBLM_R_X11Y105_SLICE_X15Y105_AO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B = CLBLM_R_X11Y105_SLICE_X15Y105_BO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C = CLBLM_R_X11Y105_SLICE_X15Y105_CO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D = CLBLM_R_X11Y105_SLICE_X15Y105_DO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_AMUX = CLBLM_R_X11Y105_SLICE_X15Y105_AO5;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_BMUX = CLBLM_R_X11Y105_SLICE_X15Y105_BO5;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A = CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B = CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C = CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D = CLBLM_R_X11Y106_SLICE_X14Y106_DO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_AMUX = CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A = CLBLM_R_X11Y106_SLICE_X15Y106_AO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B = CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C = CLBLM_R_X11Y106_SLICE_X15Y106_CO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D = CLBLM_R_X11Y106_SLICE_X15Y106_DO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_AMUX = CLBLM_R_X11Y106_SLICE_X15Y106_AO5;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A = CLBLM_R_X11Y107_SLICE_X14Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B = CLBLM_R_X11Y107_SLICE_X14Y107_BO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C = CLBLM_R_X11Y107_SLICE_X14Y107_CO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D = CLBLM_R_X11Y107_SLICE_X14Y107_DO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_AMUX = CLBLM_R_X11Y107_SLICE_X14Y107_AO5;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_BMUX = CLBLM_R_X11Y107_SLICE_X14Y107_BO5;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A = CLBLM_R_X11Y107_SLICE_X15Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B = CLBLM_R_X11Y107_SLICE_X15Y107_BO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C = CLBLM_R_X11Y107_SLICE_X15Y107_CO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D = CLBLM_R_X11Y107_SLICE_X15Y107_DO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_AMUX = CLBLM_R_X11Y107_SLICE_X15Y107_AO5;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_BMUX = CLBLM_R_X11Y107_SLICE_X15Y107_BO5;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_CMUX = CLBLM_R_X11Y107_SLICE_X15Y107_CO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A = CLBLM_R_X11Y108_SLICE_X14Y108_AO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B = CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C = CLBLM_R_X11Y108_SLICE_X14Y108_CO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D = CLBLM_R_X11Y108_SLICE_X14Y108_DO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_BMUX = CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A = CLBLM_R_X11Y108_SLICE_X15Y108_AO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B = CLBLM_R_X11Y108_SLICE_X15Y108_BO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C = CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D = CLBLM_R_X11Y108_SLICE_X15Y108_DO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_AMUX = CLBLM_R_X11Y108_SLICE_X15Y108_AO5;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_CMUX = CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A = CLBLM_R_X11Y109_SLICE_X14Y109_AO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B = CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C = CLBLM_R_X11Y109_SLICE_X14Y109_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D = CLBLM_R_X11Y109_SLICE_X14Y109_DO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A = CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B = CLBLM_R_X11Y109_SLICE_X15Y109_BO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C = CLBLM_R_X11Y109_SLICE_X15Y109_CO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D = CLBLM_R_X11Y109_SLICE_X15Y109_DO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_BMUX = CLBLM_R_X11Y109_SLICE_X15Y109_BO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A = CLBLM_R_X11Y110_SLICE_X14Y110_AO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B = CLBLM_R_X11Y110_SLICE_X14Y110_BO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C = CLBLM_R_X11Y110_SLICE_X14Y110_CO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D = CLBLM_R_X11Y110_SLICE_X14Y110_DO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_AMUX = CLBLM_R_X11Y110_SLICE_X14Y110_AO5;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A = CLBLM_R_X11Y110_SLICE_X15Y110_AO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B = CLBLM_R_X11Y110_SLICE_X15Y110_BO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C = CLBLM_R_X11Y110_SLICE_X15Y110_CO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D = CLBLM_R_X11Y110_SLICE_X15Y110_DO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_AMUX = CLBLM_R_X11Y110_SLICE_X15Y110_AO5;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_CMUX = CLBLM_R_X11Y110_SLICE_X15Y110_CO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A = CLBLM_R_X11Y111_SLICE_X14Y111_AO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B = CLBLM_R_X11Y111_SLICE_X14Y111_BO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C = CLBLM_R_X11Y111_SLICE_X14Y111_CO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D = CLBLM_R_X11Y111_SLICE_X14Y111_DO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_AMUX = CLBLM_R_X11Y111_SLICE_X14Y111_AO5;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A = CLBLM_R_X11Y111_SLICE_X15Y111_AO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B = CLBLM_R_X11Y111_SLICE_X15Y111_BO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C = CLBLM_R_X11Y111_SLICE_X15Y111_CO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D = CLBLM_R_X11Y111_SLICE_X15Y111_DO6;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_O = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_O = LIOB33_X0Y101_IOB_X0Y101_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_O = LIOB33_X0Y103_IOB_X0Y104_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_O = LIOB33_X0Y103_IOB_X0Y103_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_O = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_O = LIOB33_X0Y105_IOB_X0Y105_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_O = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_O = LIOB33_X0Y109_IOB_X0Y109_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_O = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_O = LIOB33_X0Y111_IOB_X0Y111_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_O = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_O = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_O = LIOB33_X0Y117_IOB_X0Y117_I;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_OQ = CLBLL_L_X2Y111_SLICE_X0Y111_AO5;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = CLBLL_L_X2Y110_SLICE_X0Y110_BO6;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = CLBLL_L_X2Y110_SLICE_X0Y110_BO5;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = CLBLL_L_X2Y109_SLICE_X0Y109_DO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_OQ = CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_OQ = CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_OQ = CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_OQ = CLBLL_L_X2Y111_SLICE_X0Y111_BO5;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_OQ = CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_OQ = CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_OQ = 1'b0;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_OQ = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_OQ = CLBLM_R_X3Y112_SLICE_X3Y112_BO5;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = CLBLL_L_X4Y114_SLICE_X5Y114_AO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = CLBLL_L_X4Y114_SLICE_X5Y114_AO5;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_OQ = CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_OQ = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_OQ = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_OQ = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_OQ = CLBLM_R_X5Y113_SLICE_X7Y113_CO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_OQ = CLBLM_R_X5Y113_SLICE_X6Y113_AO5;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_TQ = 1'b1;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_O = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O = LIOB33_X0Y107_IOB_X0Y107_I;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = CLBLL_L_X2Y110_SLICE_X0Y110_CO5;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = CLBLL_L_X2Y110_SLICE_X0Y110_AO5;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ = CLBLL_L_X2Y111_SLICE_X1Y111_AO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ = CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ = CLBLL_L_X4Y115_SLICE_X5Y115_AO5;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ = CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O = LIOB33_X0Y113_IOB_X0Y113_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C6 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D1 = CLBLM_L_X10Y103_SLICE_X12Y103_CO5;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D2 = CLBLM_R_X11Y104_SLICE_X14Y104_AO5;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D3 = CLBLM_L_X10Y103_SLICE_X12Y103_AO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D4 = CLBLM_L_X10Y103_SLICE_X12Y103_AO5;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D5 = CLBLM_L_X8Y102_SLICE_X11Y102_AO5;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D6 = CLBLM_L_X10Y104_SLICE_X12Y104_DO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign LIOB33_X0Y147_IOB_X0Y147_O = CLBLM_R_X5Y113_SLICE_X6Y113_AO5;
  assign LIOB33_X0Y147_IOB_X0Y148_O = CLBLM_R_X5Y113_SLICE_X7Y113_CO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A6 = CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A2 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A5 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A6 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B1 = CLBLM_R_X11Y105_SLICE_X15Y105_AO5;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B2 = CLBLM_L_X10Y104_SLICE_X12Y104_DO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B5 = CLBLM_R_X11Y104_SLICE_X14Y104_AO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B6 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C1 = CLBLM_L_X10Y103_SLICE_X12Y103_AO5;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C2 = CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C3 = CLBLM_R_X11Y105_SLICE_X15Y105_AO5;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C4 = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C5 = CLBLM_L_X10Y104_SLICE_X13Y104_AO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C6 = CLBLM_R_X11Y104_SLICE_X14Y104_AO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B3 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D1 = CLBLM_L_X10Y104_SLICE_X13Y104_AO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D2 = CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D3 = CLBLM_R_X11Y104_SLICE_X14Y104_AO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D4 = CLBLM_R_X11Y105_SLICE_X15Y105_AO5;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D5 = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D6 = CLBLM_L_X10Y103_SLICE_X12Y103_AO5;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B4 = 1'b1;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A1 = CLBLM_L_X10Y103_SLICE_X12Y103_DO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A2 = CLBLM_L_X8Y102_SLICE_X11Y102_CO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A3 = CLBLM_L_X10Y104_SLICE_X13Y104_CO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A4 = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A5 = CLBLM_L_X10Y103_SLICE_X12Y103_BO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A6 = CLBLM_L_X10Y103_SLICE_X12Y103_BO5;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B1 = CLBLM_L_X10Y104_SLICE_X12Y104_DO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B2 = CLBLM_L_X10Y103_SLICE_X12Y103_AO5;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B3 = CLBLM_L_X10Y103_SLICE_X12Y103_AO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B4 = CLBLM_R_X11Y104_SLICE_X14Y104_AO5;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B5 = CLBLM_L_X10Y103_SLICE_X12Y103_CO5;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B6 = CLBLM_L_X8Y102_SLICE_X11Y102_AO5;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C1 = CLBLM_L_X10Y103_SLICE_X12Y103_CO5;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C5 = CLBLM_L_X10Y104_SLICE_X12Y104_DO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C6 = CLBLM_R_X11Y104_SLICE_X14Y104_AO5;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D2 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D4 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B2 = CLBLM_L_X10Y103_SLICE_X12Y103_BO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B3 = CLBLM_R_X7Y104_SLICE_X8Y104_AO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B4 = CLBLM_R_X7Y102_SLICE_X9Y102_CO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A1 = CLBLM_R_X11Y105_SLICE_X15Y105_AO5;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A3 = CLBLM_R_X11Y104_SLICE_X14Y104_AO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A5 = CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A6 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B1 = CLBLM_L_X8Y103_SLICE_X10Y103_DO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B2 = CLBLM_L_X10Y105_SLICE_X12Y105_DO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B3 = CLBLM_L_X10Y105_SLICE_X12Y105_CO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B4 = CLBLM_L_X10Y109_SLICE_X12Y109_AO5;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B5 = CLBLM_R_X11Y105_SLICE_X15Y105_BO5;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B6 = CLBLM_L_X8Y105_SLICE_X10Y105_AO5;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C1 = CLBLM_L_X10Y105_SLICE_X13Y105_AO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C2 = CLBLM_L_X10Y103_SLICE_X13Y103_AO5;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C6 = CLBLM_L_X10Y104_SLICE_X13Y104_BO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D1 = CLBLM_R_X11Y105_SLICE_X15Y105_BO5;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D2 = CLBLM_L_X10Y105_SLICE_X12Y105_CO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D3 = CLBLM_L_X10Y105_SLICE_X12Y105_DO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D4 = CLBLM_L_X8Y105_SLICE_X10Y105_AO5;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D5 = CLBLM_L_X8Y103_SLICE_X10Y103_DO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D6 = CLBLM_L_X10Y109_SLICE_X12Y109_AO5;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A3 = CLBLM_L_X10Y105_SLICE_X13Y105_AO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A5 = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B1 = CLBLM_L_X8Y103_SLICE_X10Y103_DO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B4 = CLBLM_L_X10Y105_SLICE_X12Y105_DO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B5 = CLBLM_L_X10Y105_SLICE_X12Y105_CO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C1 = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C2 = CLBLM_L_X10Y105_SLICE_X13Y105_AO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D1 = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D2 = CLBLM_L_X10Y103_SLICE_X12Y103_BO5;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D3 = CLBLM_L_X10Y104_SLICE_X13Y104_AO5;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D4 = CLBLM_L_X10Y104_SLICE_X13Y104_CO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D5 = CLBLM_R_X11Y105_SLICE_X14Y105_DO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D6 = CLBLM_L_X10Y104_SLICE_X13Y104_DO6;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_A1 = CLBLM_R_X5Y102_SLICE_X6Y102_CO6;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_A2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_A3 = CLBLM_R_X7Y102_SLICE_X8Y102_BO5;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_B5 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A6 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B1 = CLBLM_L_X10Y106_SLICE_X13Y106_DO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B2 = CLBLM_L_X10Y109_SLICE_X12Y109_AO5;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B3 = CLBLM_L_X10Y108_SLICE_X13Y108_AO5;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B4 = CLBLM_L_X10Y106_SLICE_X12Y106_DO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B5 = CLBLM_L_X10Y105_SLICE_X12Y105_AO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B6 = CLBLM_L_X10Y107_SLICE_X13Y107_AO5;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C1 = CLBLM_L_X10Y105_SLICE_X12Y105_AO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C2 = CLBLM_L_X10Y107_SLICE_X13Y107_AO5;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C3 = CLBLM_L_X10Y109_SLICE_X12Y109_AO5;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C4 = CLBLM_L_X10Y108_SLICE_X13Y108_AO5;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C5 = CLBLM_L_X10Y106_SLICE_X13Y106_DO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C6 = CLBLM_L_X10Y106_SLICE_X12Y106_DO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D1 = CLBLM_R_X11Y105_SLICE_X14Y105_BO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D2 = CLBLM_L_X10Y104_SLICE_X13Y104_AO5;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D3 = CLBLM_R_X11Y107_SLICE_X14Y107_DO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D4 = CLBLM_L_X10Y104_SLICE_X13Y104_DO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D5 = CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D6 = CLBLM_R_X11Y105_SLICE_X14Y105_DO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A1 = CLBLM_R_X11Y105_SLICE_X14Y105_CO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A3 = CLBLM_L_X10Y105_SLICE_X12Y105_AO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B1 = CLBLM_L_X10Y104_SLICE_X13Y104_DO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B6 = CLBLM_R_X11Y105_SLICE_X15Y105_CO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C1 = CLBLM_L_X10Y105_SLICE_X12Y105_AO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C2 = CLBLM_L_X10Y109_SLICE_X12Y109_AO5;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C3 = CLBLM_L_X10Y108_SLICE_X13Y108_AO5;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C4 = CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C5 = CLBLM_L_X10Y106_SLICE_X12Y106_DO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C6 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D3 = CLBLM_L_X10Y104_SLICE_X13Y104_DO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D4 = CLBLM_R_X11Y105_SLICE_X15Y105_CO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C2 = CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C3 = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C4 = CLBLL_L_X4Y109_SLICE_X4Y109_AO5;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A1 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A3 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A6 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C1 = CLBLM_R_X11Y111_SLICE_X14Y111_BO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B1 = CLBLM_L_X10Y107_SLICE_X12Y107_AO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B2 = CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B3 = CLBLM_R_X11Y105_SLICE_X14Y105_BO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B4 = CLBLM_R_X11Y107_SLICE_X14Y107_CO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B5 = CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B6 = CLBLM_R_X11Y107_SLICE_X14Y107_DO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C1 = CLBLM_R_X11Y108_SLICE_X15Y108_AO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C2 = CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C6 = CLBLM_R_X11Y107_SLICE_X14Y107_AO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D1 = CLBLM_R_X11Y108_SLICE_X15Y108_AO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D2 = CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D6 = CLBLM_R_X11Y107_SLICE_X14Y107_AO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A1 = CLBLM_L_X10Y110_SLICE_X13Y110_AO5;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A3 = CLBLM_R_X11Y107_SLICE_X14Y107_BO5;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A6 = CLBLM_L_X10Y107_SLICE_X12Y107_CO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B1 = CLBLM_L_X10Y110_SLICE_X13Y110_AO5;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B3 = CLBLM_R_X11Y107_SLICE_X14Y107_BO5;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B6 = CLBLM_L_X10Y107_SLICE_X12Y107_CO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C6 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D1 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D2 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D3 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D4 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D5 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D6 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_T1 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B2 = CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B3 = CLBLM_L_X10Y111_SLICE_X13Y111_AO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A2 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A4 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A5 = CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A6 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A1 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A2 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A6 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C1 = CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B1 = CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B2 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B3 = CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B4 = CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B5 = CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B6 = CLBLM_L_X10Y108_SLICE_X13Y108_AO5;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C2 = CLBLM_R_X11Y110_SLICE_X15Y110_BO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C1 = CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C2 = CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C3 = CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C4 = CLBLM_L_X10Y108_SLICE_X13Y108_AO5;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C5 = CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C6 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D1 = CLBLM_L_X10Y109_SLICE_X13Y109_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D2 = CLBLM_R_X11Y107_SLICE_X14Y107_AO5;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D3 = CLBLM_R_X11Y108_SLICE_X14Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D6 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A1 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A5 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A6 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B1 = CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B2 = CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B3 = CLBLM_R_X11Y108_SLICE_X14Y108_DO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B4 = CLBLM_R_X11Y108_SLICE_X14Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B5 = CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B6 = CLBLM_L_X10Y108_SLICE_X12Y108_AO5;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C1 = CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C2 = CLBLM_L_X8Y106_SLICE_X11Y106_AO5;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C3 = CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C4 = CLBLM_L_X10Y108_SLICE_X12Y108_AO5;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C5 = CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C6 = CLBLM_R_X11Y108_SLICE_X14Y108_DO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D1 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D2 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D3 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D4 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D6 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A1 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A4 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A6 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B1 = CLBLM_R_X5Y101_SLICE_X6Y101_AO5;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B2 = CLBLM_R_X3Y104_SLICE_X2Y104_AO5;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B3 = CLBLM_R_X3Y103_SLICE_X3Y103_AO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B4 = CLBLM_R_X5Y102_SLICE_X6Y102_AO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B5 = CLBLL_L_X4Y104_SLICE_X4Y104_AO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B6 = CLBLM_R_X3Y104_SLICE_X2Y104_BO5;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C1 = CLBLL_L_X4Y104_SLICE_X4Y104_AO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C2 = CLBLM_R_X3Y103_SLICE_X3Y103_AO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C3 = CLBLM_R_X5Y101_SLICE_X6Y101_AO5;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C4 = CLBLM_R_X3Y104_SLICE_X2Y104_BO5;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C5 = CLBLM_R_X3Y104_SLICE_X2Y104_AO5;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C6 = CLBLM_R_X5Y102_SLICE_X6Y102_AO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D3 = CLBLM_R_X5Y101_SLICE_X6Y101_BO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D4 = CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B6 = CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A1 = CLBLL_L_X4Y105_SLICE_X5Y105_BO5;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A2 = CLBLM_R_X5Y103_SLICE_X6Y103_CO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A3 = CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A4 = CLBLL_L_X4Y104_SLICE_X5Y104_BO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A5 = CLBLM_R_X5Y103_SLICE_X6Y103_BO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A6 = CLBLL_L_X4Y105_SLICE_X5Y105_AO5;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B4 = CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B6 = CLBLM_R_X5Y101_SLICE_X6Y101_BO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C1 = CLBLM_R_X5Y103_SLICE_X6Y103_BO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C2 = CLBLM_R_X5Y103_SLICE_X6Y103_CO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C6 = CLBLL_L_X4Y104_SLICE_X5Y104_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C4 = CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D1 = CLBLM_R_X5Y103_SLICE_X6Y103_BO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D2 = CLBLM_R_X5Y103_SLICE_X6Y103_CO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D3 = CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D4 = CLBLL_L_X4Y105_SLICE_X5Y105_AO5;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D5 = CLBLL_L_X4Y105_SLICE_X5Y105_BO5;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D6 = CLBLL_L_X4Y104_SLICE_X5Y104_BO6;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_D = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_D = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A2 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A4 = CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A5 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A6 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B2 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B4 = CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B5 = CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B6 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C2 = CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C5 = CLBLM_R_X11Y108_SLICE_X14Y108_AO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D2 = CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D5 = CLBLM_R_X11Y108_SLICE_X14Y108_AO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A1 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A2 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A6 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B1 = CLBLM_R_X7Y109_SLICE_X8Y109_AO5;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B2 = CLBLM_R_X11Y109_SLICE_X14Y109_DO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B3 = CLBLM_L_X8Y108_SLICE_X11Y108_DO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B4 = CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B5 = CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B6 = CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C1 = CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C2 = CLBLM_L_X8Y108_SLICE_X11Y108_DO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C3 = CLBLM_R_X11Y109_SLICE_X14Y109_DO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C4 = CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C5 = CLBLM_R_X7Y109_SLICE_X8Y109_AO5;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C6 = CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D1 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D2 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D3 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D4 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D5 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D6 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A1 = CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A2 = CLBLM_R_X5Y105_SLICE_X6Y105_BO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A6 = CLBLL_L_X4Y104_SLICE_X4Y104_DO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B1 = CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B2 = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B3 = CLBLL_L_X4Y105_SLICE_X5Y105_AO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B4 = CLBLL_L_X4Y105_SLICE_X5Y105_AO5;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B5 = CLBLM_R_X5Y105_SLICE_X6Y105_BO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B6 = CLBLL_L_X4Y104_SLICE_X4Y104_DO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C1 = CLBLM_R_X5Y105_SLICE_X6Y105_BO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C2 = CLBLL_L_X4Y105_SLICE_X5Y105_AO5;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C3 = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C4 = CLBLL_L_X4Y104_SLICE_X4Y104_DO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C5 = CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C6 = CLBLL_L_X4Y105_SLICE_X5Y105_AO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D1 = CLBLM_R_X3Y104_SLICE_X3Y104_DO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D3 = CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A1 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A5 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A6 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B1 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B3 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B6 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C2 = CLBLL_L_X4Y105_SLICE_X5Y105_DO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C3 = CLBLL_L_X4Y105_SLICE_X4Y105_DO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C4 = CLBLL_L_X4Y104_SLICE_X5Y104_CO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D1 = CLBLM_R_X5Y101_SLICE_X6Y101_CO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D6 = CLBLL_L_X4Y104_SLICE_X5Y104_BO6;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A3 = CLBLM_L_X8Y104_SLICE_X11Y104_AO6;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B4 = CLBLM_R_X7Y104_SLICE_X9Y104_AO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B5 = CLBLM_L_X8Y105_SLICE_X10Y105_AO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B6 = CLBLM_R_X7Y105_SLICE_X8Y105_AO5;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A2 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A6 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B1 = CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B5 = CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C1 = CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C3 = CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D2 = CLBLM_R_X11Y110_SLICE_X14Y110_DO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D4 = CLBLM_L_X10Y111_SLICE_X13Y111_DO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A2 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A3 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A6 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B1 = CLBLM_L_X10Y110_SLICE_X12Y110_DO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B2 = CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B3 = CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B4 = CLBLM_L_X10Y111_SLICE_X12Y111_BO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B5 = CLBLM_L_X10Y110_SLICE_X12Y110_AO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B6 = CLBLM_L_X10Y110_SLICE_X12Y110_AO5;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C1 = CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C2 = CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C3 = CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C4 = CLBLM_L_X10Y112_SLICE_X12Y112_AO5;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C5 = CLBLM_L_X10Y112_SLICE_X13Y112_AO5;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C6 = CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A3 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A5 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A6 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D1 = CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D2 = CLBLM_L_X10Y112_SLICE_X12Y112_AO5;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D3 = CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B2 = CLBLM_R_X3Y106_SLICE_X3Y106_CO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B3 = CLBLM_R_X3Y107_SLICE_X3Y107_DO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B6 = CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C1 = CLBLL_L_X4Y104_SLICE_X5Y104_AO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C2 = CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C3 = CLBLL_L_X4Y106_SLICE_X4Y106_AO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C4 = CLBLL_L_X4Y106_SLICE_X4Y106_AO5;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C5 = CLBLM_R_X3Y106_SLICE_X2Y106_DO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C6 = CLBLL_L_X4Y105_SLICE_X4Y105_BO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D1 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D2 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D3 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D4 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D5 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D6 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_A1 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_A2 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_A3 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_A4 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_A5 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_A6 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A1 = CLBLL_L_X4Y104_SLICE_X5Y104_DO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A2 = CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A3 = CLBLL_L_X4Y106_SLICE_X4Y106_AO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A4 = CLBLM_R_X5Y104_SLICE_X6Y104_AO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A5 = CLBLL_L_X4Y104_SLICE_X5Y104_AO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A6 = CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_A1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_B1 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_B2 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B1 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B2 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B3 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B4 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B5 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B6 = 1'b1;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_A3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_C1 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C1 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C2 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C3 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C4 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C5 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C6 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_D1 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_D2 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_D3 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_D4 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_D5 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_D6 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D1 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D2 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D3 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D4 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D5 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D6 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_A2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_A3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_A4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_A5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_A6 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_B1 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_B2 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_B3 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_B4 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_B5 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_B6 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_C1 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_C2 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_C3 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_C4 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_C5 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_C6 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_D1 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_D2 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_D3 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_D4 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_D5 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_D6 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D5 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A2 = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A4 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A5 = CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A6 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D6 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B1 = CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B3 = CLBLM_R_X11Y110_SLICE_X14Y110_AO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B4 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B6 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C2 = CLBLM_R_X11Y110_SLICE_X14Y110_DO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C6 = CLBLM_L_X10Y111_SLICE_X13Y111_DO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D1 = CLBLM_L_X12Y110_SLICE_X16Y110_CO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D4 = CLBLM_R_X11Y110_SLICE_X15Y110_DO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A2 = CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A3 = CLBLM_L_X10Y111_SLICE_X13Y111_AO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A6 = CLBLM_L_X10Y111_SLICE_X12Y111_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B1 = CLBLM_L_X10Y112_SLICE_X13Y112_AO5;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B2 = CLBLM_L_X10Y111_SLICE_X13Y111_BO5;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B3 = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B4 = CLBLM_R_X11Y109_SLICE_X14Y109_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B5 = CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B6 = CLBLM_R_X7Y108_SLICE_X9Y108_AO5;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C1 = CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C4 = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C6 = CLBLM_R_X11Y109_SLICE_X14Y109_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A1 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A5 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D1 = CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A6 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D2 = CLBLM_R_X7Y108_SLICE_X9Y108_AO5;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D4 = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B1 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B5 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B6 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D3 = CLBLM_L_X10Y111_SLICE_X13Y111_BO5;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D5 = CLBLM_L_X10Y112_SLICE_X13Y112_AO5;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D6 = CLBLM_R_X11Y109_SLICE_X14Y109_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C1 = CLBLL_L_X4Y105_SLICE_X4Y105_AO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C3 = CLBLM_R_X3Y106_SLICE_X2Y106_DO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_A5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D1 = CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D2 = CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D3 = CLBLM_R_X3Y106_SLICE_X3Y106_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D4 = CLBLL_L_X4Y107_SLICE_X4Y107_AO5;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D5 = CLBLM_R_X3Y107_SLICE_X3Y107_DO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D6 = CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A4 = CLBLL_L_X4Y104_SLICE_X5Y104_CO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A6 = CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A6 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B2 = CLBLL_L_X4Y104_SLICE_X5Y104_CO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B6 = CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B4 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B6 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C3 = CLBLM_R_X5Y105_SLICE_X6Y105_CO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C6 = CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C3 = CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C4 = CLBLM_R_X11Y106_SLICE_X15Y106_AO5;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C6 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D1 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D2 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D3 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D1 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D2 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D3 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D4 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D5 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D6 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D4 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D5 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A1 = CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C1 = CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A2 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A6 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B1 = CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B2 = CLBLM_R_X11Y107_SLICE_X15Y107_AO5;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B3 = CLBLM_R_X11Y105_SLICE_X15Y105_AO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B4 = CLBLM_R_X11Y106_SLICE_X15Y106_AO5;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B5 = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B6 = CLBLM_R_X11Y105_SLICE_X14Y105_AO5;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C1 = CLBLM_R_X11Y105_SLICE_X14Y105_AO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C2 = CLBLM_R_X11Y105_SLICE_X15Y105_CO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C3 = CLBLM_L_X10Y104_SLICE_X13Y104_BO5;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C6 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D1 = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D2 = CLBLM_R_X11Y107_SLICE_X15Y107_AO5;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D3 = CLBLM_R_X11Y105_SLICE_X15Y105_AO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D4 = CLBLM_R_X11Y105_SLICE_X14Y105_AO5;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D5 = CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D6 = CLBLM_R_X11Y106_SLICE_X15Y106_AO5;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A1 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A3 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_A6 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B3 = CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B4 = CLBLM_L_X10Y111_SLICE_X12Y111_BO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B5 = CLBLM_L_X10Y111_SLICE_X13Y111_AO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_B6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_A1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_A2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_A3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C4 = CLBLM_L_X10Y111_SLICE_X13Y111_AO5;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_A4 = 1'b1;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_A5 = 1'b1;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_A6 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_C2 = CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_B1 = CLBLM_L_X10Y103_SLICE_X12Y103_AO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_B2 = CLBLM_R_X7Y102_SLICE_X9Y102_AO5;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_B3 = CLBLM_L_X8Y102_SLICE_X10Y102_AO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D1 = CLBLM_R_X11Y111_SLICE_X14Y111_BO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_B4 = CLBLM_L_X10Y103_SLICE_X12Y103_CO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D2 = CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D4 = CLBLM_L_X10Y111_SLICE_X13Y111_AO5;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_B5 = CLBLM_L_X8Y102_SLICE_X11Y102_AO6;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X10Y112_SLICE_X13Y112_D6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_B6 = CLBLM_L_X10Y103_SLICE_X13Y103_BO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_C1 = CLBLM_L_X8Y102_SLICE_X11Y102_AO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_C2 = CLBLM_L_X8Y102_SLICE_X10Y102_AO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_C3 = CLBLM_L_X10Y103_SLICE_X12Y103_CO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_C4 = CLBLM_L_X10Y103_SLICE_X12Y103_AO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_C5 = CLBLM_L_X10Y103_SLICE_X13Y103_BO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_C6 = CLBLM_R_X7Y102_SLICE_X9Y102_AO5;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A2 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A3 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_A6 = 1'b1;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_D1 = 1'b1;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_D2 = 1'b1;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_D3 = 1'b1;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_D4 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B5 = CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_D5 = 1'b1;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_D6 = 1'b1;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B6 = CLBLM_L_X10Y112_SLICE_X12Y112_AO5;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C1 = CLBLM_L_X10Y111_SLICE_X13Y111_AO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_B4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C4 = CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_C6 = CLBLM_L_X10Y111_SLICE_X12Y111_BO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_A1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_A2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_A3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_A4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_A5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_A6 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A2 = CLBLL_L_X4Y105_SLICE_X5Y105_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D1 = CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D2 = CLBLM_L_X10Y111_SLICE_X13Y111_AO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D3 = CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D4 = CLBLM_L_X10Y112_SLICE_X12Y112_AO5;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y112_SLICE_X12Y112_D6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B1 = CLBLL_L_X4Y107_SLICE_X5Y107_AO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B5 = CLBLL_L_X4Y106_SLICE_X5Y106_AO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B6 = CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_C4 = 1'b1;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_C5 = 1'b1;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_C6 = 1'b1;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_D1 = 1'b1;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_D2 = 1'b1;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_D3 = 1'b1;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_D4 = 1'b1;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_D5 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D1 = CLBLL_L_X4Y106_SLICE_X5Y106_AO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D2 = CLBLL_L_X4Y107_SLICE_X5Y107_AO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D3 = CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D4 = CLBLL_L_X4Y107_SLICE_X4Y107_AO5;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D5 = CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D6 = CLBLL_L_X4Y107_SLICE_X4Y107_BO5;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_D6 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A2 = CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A4 = CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A5 = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B5 = CLBLL_L_X4Y105_SLICE_X5Y105_CO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B6 = CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C1 = CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C5 = CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C6 = CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C1 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C2 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C3 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C4 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C5 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A6 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C6 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D1 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D2 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D3 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D4 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D5 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D6 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D4 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D5 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D6 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D3 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A5 = CLBLM_L_X10Y105_SLICE_X12Y105_AO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A6 = CLBLM_R_X11Y105_SLICE_X14Y105_CO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B1 = CLBLM_R_X11Y106_SLICE_X14Y106_DO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B5 = CLBLM_R_X11Y105_SLICE_X14Y105_BO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C1 = CLBLM_R_X11Y105_SLICE_X14Y105_BO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C5 = CLBLM_R_X11Y106_SLICE_X14Y106_DO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C6 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D2 = CLBLM_R_X11Y106_SLICE_X15Y106_AO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D3 = CLBLM_R_X11Y107_SLICE_X14Y107_BO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D5 = CLBLM_L_X12Y107_SLICE_X16Y107_AO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D6 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C1 = CLBLM_R_X11Y111_SLICE_X14Y111_BO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C3 = CLBLM_R_X11Y111_SLICE_X14Y111_AO5;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C4 = CLBLM_L_X10Y112_SLICE_X13Y112_AO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C5 = CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C6 = CLBLM_R_X11Y111_SLICE_X14Y111_CO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A2 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A3 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A4 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A5 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_A6 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B2 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B3 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B4 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B5 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_B6 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C2 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C3 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C4 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C5 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_C6 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A2 = CLBLM_L_X10Y103_SLICE_X13Y103_BO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A5 = CLBLM_L_X8Y102_SLICE_X10Y102_AO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B2 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A6 = CLBLM_L_X10Y103_SLICE_X12Y103_CO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B5 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D2 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D3 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D4 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D5 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X13Y113_D6 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B6 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C1 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C2 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C3 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C4 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C5 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C6 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A1 = CLBLM_R_X11Y111_SLICE_X14Y111_AO5;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A2 = CLBLM_R_X11Y111_SLICE_X14Y111_CO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_A5 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B1 = CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B2 = CLBLM_L_X10Y110_SLICE_X12Y110_AO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B3 = CLBLM_L_X10Y112_SLICE_X13Y112_AO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B4 = CLBLM_L_X10Y111_SLICE_X12Y111_BO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D1 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D2 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D3 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B5 = CLBLM_R_X11Y111_SLICE_X14Y111_BO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_B6 = CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D5 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D6 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A3 = CLBLM_L_X8Y102_SLICE_X10Y102_AO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A4 = CLBLM_R_X7Y103_SLICE_X9Y103_AO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A5 = CLBLM_L_X10Y103_SLICE_X12Y103_CO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A5 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A6 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_C2 = CLBLM_L_X10Y113_SLICE_X12Y113_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B2 = CLBLL_L_X4Y109_SLICE_X5Y109_BO5;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B5 = CLBLM_L_X8Y102_SLICE_X11Y102_BO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B6 = CLBLM_L_X8Y102_SLICE_X11Y102_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B3 = CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B1 = CLBLM_L_X10Y103_SLICE_X12Y103_DO6;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D3 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C1 = CLBLM_L_X8Y103_SLICE_X10Y103_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C1 = CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B6 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D1 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D2 = 1'b1;
  assign CLBLM_L_X10Y113_SLICE_X12Y113_D4 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C4 = CLBLM_L_X10Y103_SLICE_X13Y103_AO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C5 = CLBLM_L_X10Y104_SLICE_X12Y104_CO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C5 = CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C6 = CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D1 = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D2 = CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D3 = CLBLL_L_X4Y109_SLICE_X5Y109_BO5;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D4 = CLBLL_L_X4Y109_SLICE_X4Y109_AO5;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D5 = CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D4 = CLBLM_L_X8Y102_SLICE_X11Y102_CO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D5 = CLBLM_L_X10Y104_SLICE_X12Y104_CO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D6 = CLBLM_R_X3Y109_SLICE_X3Y109_BO5;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A3 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A5 = CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A6 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A1 = CLBLM_R_X11Y106_SLICE_X15Y106_AO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A2 = CLBLM_R_X11Y107_SLICE_X14Y107_BO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A3 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B2 = CLBLM_R_X5Y107_SLICE_X6Y107_CO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B3 = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B3 = CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B4 = CLBLM_L_X10Y112_SLICE_X12Y112_BO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C1 = CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C2 = CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C3 = CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C4 = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C5 = CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C6 = CLBLM_R_X5Y107_SLICE_X6Y107_CO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B3 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B5 = CLBLM_L_X12Y107_SLICE_X16Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B6 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C1 = CLBLM_R_X11Y107_SLICE_X15Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D1 = CLBLL_L_X4Y109_SLICE_X5Y109_BO5;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D2 = CLBLL_L_X4Y109_SLICE_X4Y109_AO5;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D3 = CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D4 = CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D5 = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D6 = CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D1 = CLBLM_R_X11Y107_SLICE_X15Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D2 = CLBLM_L_X10Y107_SLICE_X12Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D5 = CLBLM_R_X11Y107_SLICE_X15Y107_BO5;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D6 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A2 = CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A3 = CLBLM_R_X11Y107_SLICE_X15Y107_CO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A5 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A6 = 1'b1;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_D = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B6 = 1'b1;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_D = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C1 = CLBLM_R_X11Y107_SLICE_X15Y107_BO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C2 = CLBLM_R_X11Y107_SLICE_X15Y107_AO5;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C3 = CLBLM_L_X12Y107_SLICE_X16Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C4 = CLBLM_R_X7Y110_SLICE_X8Y110_AO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C5 = CLBLM_R_X11Y106_SLICE_X15Y106_AO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C6 = CLBLM_R_X11Y107_SLICE_X14Y107_BO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D1 = CLBLM_R_X11Y107_SLICE_X15Y107_BO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D2 = CLBLM_R_X11Y107_SLICE_X15Y107_AO5;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D3 = CLBLM_L_X12Y107_SLICE_X16Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D4 = CLBLM_R_X7Y110_SLICE_X8Y110_AO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D5 = CLBLM_R_X11Y106_SLICE_X15Y106_AO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D6 = CLBLM_R_X11Y107_SLICE_X14Y107_BO6;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D1 = CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D3 = CLBLM_R_X11Y111_SLICE_X14Y111_DO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A1 = CLBLM_L_X10Y104_SLICE_X12Y104_CO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A5 = CLBLM_L_X8Y102_SLICE_X11Y102_CO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B1 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B2 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B3 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B4 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B5 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B6 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C1 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C2 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C3 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C4 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C5 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C6 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D1 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D2 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D3 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D4 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D5 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D6 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A1 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A4 = CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A5 = CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A4 = CLBLM_R_X7Y104_SLICE_X9Y104_AO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A5 = CLBLM_L_X8Y105_SLICE_X10Y105_AO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A6 = CLBLM_R_X7Y105_SLICE_X8Y105_AO5;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_A6 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A1 = CLBLM_L_X8Y105_SLICE_X10Y105_AO5;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A2 = CLBLM_L_X10Y104_SLICE_X12Y104_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B2 = CLBLL_L_X4Y109_SLICE_X4Y109_BO5;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B4 = CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B3 = CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B5 = CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B6 = CLBLM_R_X3Y109_SLICE_X3Y109_BO5;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_B1 = CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B1 = CLBLM_L_X8Y105_SLICE_X10Y105_AO5;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B2 = CLBLM_L_X10Y104_SLICE_X12Y104_AO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B3 = CLBLM_L_X8Y104_SLICE_X11Y104_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C3 = CLBLL_L_X4Y112_SLICE_X4Y112_AO5;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C6 = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C5 = CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C6 = CLBLM_R_X7Y104_SLICE_X9Y104_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C2 = CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_C4 = CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C2 = CLBLM_L_X8Y103_SLICE_X10Y103_CO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D1 = CLBLL_L_X4Y110_SLICE_X4Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D2 = CLBLM_R_X3Y109_SLICE_X3Y109_BO5;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D3 = CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D4 = CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D5 = CLBLL_L_X4Y109_SLICE_X4Y109_BO5;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D2 = CLBLM_L_X8Y103_SLICE_X10Y103_CO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y110_SLICE_X4Y110_D6 = CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D6 = CLBLM_R_X7Y104_SLICE_X9Y104_AO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A2 = CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A3 = CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_A6 = CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B1 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B2 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B3 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B4 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B5 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_B6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D5 = CLBLM_R_X5Y115_SLICE_X6Y115_DO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D6 = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A1 = CLBLM_R_X11Y107_SLICE_X15Y107_DO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C1 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C2 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C3 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C4 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C5 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_C6 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B4 = CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B5 = CLBLM_R_X11Y110_SLICE_X15Y110_AO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B6 = CLBLM_L_X12Y108_SLICE_X16Y108_BO6;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D1 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D2 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D3 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D4 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D5 = 1'b1;
  assign CLBLL_L_X4Y110_SLICE_X5Y110_D6 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D1 = CLBLM_R_X11Y110_SLICE_X15Y110_AO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D2 = CLBLM_L_X12Y108_SLICE_X16Y108_BO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D6 = CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A1 = CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A5 = CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A6 = CLBLM_R_X11Y107_SLICE_X15Y107_CO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B1 = CLBLM_R_X11Y107_SLICE_X14Y107_CO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B2 = CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B3 = CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B4 = CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B5 = CLBLM_R_X11Y110_SLICE_X15Y110_AO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B6 = CLBLM_L_X10Y107_SLICE_X12Y107_AO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C1 = CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C2 = CLBLM_R_X11Y108_SLICE_X15Y108_AO5;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C3 = CLBLM_R_X11Y105_SLICE_X15Y105_BO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D3 = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C4 = CLBLM_R_X11Y107_SLICE_X15Y107_CO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C5 = CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C6 = CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D1 = CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D2 = CLBLM_R_X11Y108_SLICE_X15Y108_AO5;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D3 = CLBLM_R_X11Y105_SLICE_X15Y105_BO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D4 = CLBLM_R_X11Y107_SLICE_X15Y107_CO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D5 = CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D6 = CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C5 = CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C6 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A1 = CLBLM_L_X8Y103_SLICE_X10Y103_DO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A6 = CLBLM_L_X10Y105_SLICE_X13Y105_CO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B1 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B2 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B3 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B4 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B5 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B6 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C1 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C2 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C3 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C4 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C5 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C6 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D1 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D2 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D3 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D4 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D5 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D6 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A1 = CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A5 = CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A1 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A5 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A6 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B1 = CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B1 = CLBLM_L_X8Y104_SLICE_X10Y104_DO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C2 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C3 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B4 = CLBLM_L_X10Y105_SLICE_X12Y105_BO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B6 = CLBLM_L_X8Y105_SLICE_X10Y105_CO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C1 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C2 = CLBLM_L_X10Y105_SLICE_X13Y105_CO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C3 = CLBLM_L_X8Y103_SLICE_X10Y103_DO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D1 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D2 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D3 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D4 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D5 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D6 = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_D = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D1 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D2 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D3 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D4 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D5 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D6 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A1 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A2 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A3 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A4 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A5 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A6 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B1 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B2 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B3 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B4 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B5 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B6 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A1 = CLBLM_R_X11Y107_SLICE_X15Y107_DO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A2 = CLBLM_R_X11Y108_SLICE_X15Y108_DO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C1 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C2 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C3 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C4 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C5 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C6 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A5 = CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B1 = CLBLM_R_X11Y107_SLICE_X15Y107_DO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B2 = CLBLM_R_X11Y108_SLICE_X15Y108_DO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B3 = CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D1 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D2 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D3 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D4 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D5 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D6 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C1 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C2 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C3 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C4 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C5 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C6 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D1 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D2 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D3 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D4 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D5 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A2 = CLBLM_L_X10Y109_SLICE_X13Y109_AO5;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A3 = CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A5 = CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B2 = CLBLM_L_X10Y109_SLICE_X13Y109_AO5;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B3 = CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B6 = CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C1 = CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C2 = CLBLM_R_X11Y110_SLICE_X14Y110_AO5;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C3 = CLBLM_R_X11Y109_SLICE_X15Y109_BO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C4 = CLBLM_R_X11Y108_SLICE_X14Y108_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C5 = CLBLM_R_X11Y110_SLICE_X15Y110_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C6 = CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D1 = CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D3 = CLBLM_L_X10Y109_SLICE_X13Y109_AO5;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D4 = CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_D = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_D = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A1 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A2 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A6 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B3 = CLBLM_L_X8Y105_SLICE_X11Y105_AO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B4 = CLBLM_L_X10Y106_SLICE_X12Y106_AO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B6 = CLBLM_L_X10Y106_SLICE_X12Y106_CO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C1 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C2 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C3 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C4 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C5 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C6 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D5 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A4 = CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A5 = CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A6 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D2 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D3 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A1 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A2 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A3 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A4 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A5 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C1 = CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C2 = CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B1 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B2 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B3 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B4 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B5 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D1 = CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D2 = CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C1 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C2 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C3 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C4 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C5 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C6 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D1 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D2 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D3 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D4 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D5 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A1 = CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A2 = CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A6 = CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B2 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B3 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B4 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B5 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B6 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B3 = CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C2 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C3 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C4 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C5 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C6 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A1 = CLBLM_L_X12Y110_SLICE_X16Y110_DO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A4 = CLBLM_R_X11Y110_SLICE_X15Y110_BO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D2 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D3 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D4 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D5 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D6 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B6 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C1 = CLBLM_R_X11Y108_SLICE_X15Y108_BO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C4 = CLBLM_L_X12Y110_SLICE_X16Y110_DO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D2 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D6 = CLBLM_L_X12Y110_SLICE_X17Y110_AO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A1 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A2 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C4 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A3 = CLBLM_R_X11Y110_SLICE_X15Y110_CO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A4 = CLBLM_R_X11Y109_SLICE_X15Y109_BO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A6 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C5 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C6 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B2 = CLBLM_L_X12Y110_SLICE_X17Y110_BO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B3 = CLBLM_R_X11Y110_SLICE_X15Y110_CO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B6 = CLBLM_R_X11Y109_SLICE_X15Y109_BO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C1 = CLBLM_L_X12Y110_SLICE_X17Y110_BO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C2 = CLBLM_R_X11Y110_SLICE_X15Y110_CO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C4 = CLBLM_R_X11Y109_SLICE_X15Y109_BO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C6 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D2 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D4 = CLBLM_L_X12Y110_SLICE_X17Y110_AO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A3 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A5 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A6 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B3 = CLBLM_L_X8Y104_SLICE_X10Y104_BO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B6 = CLBLM_L_X10Y105_SLICE_X12Y105_BO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C1 = CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C2 = CLBLM_L_X8Y104_SLICE_X10Y104_BO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C3 = CLBLM_L_X10Y105_SLICE_X13Y105_BO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C4 = CLBLM_L_X8Y107_SLICE_X11Y107_AO5;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C5 = CLBLM_L_X10Y105_SLICE_X13Y105_DO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C6 = CLBLM_L_X10Y106_SLICE_X13Y106_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A6 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D1 = CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D4 = CLBLM_L_X8Y107_SLICE_X11Y107_AO5;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B2 = CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B3 = CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B6 = CLBLM_R_X7Y109_SLICE_X9Y109_BO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D5 = CLBLM_L_X10Y105_SLICE_X13Y105_DO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C1 = CLBLL_L_X4Y110_SLICE_X4Y110_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C2 = CLBLM_R_X7Y113_SLICE_X8Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C3 = CLBLM_R_X3Y112_SLICE_X3Y112_AO5;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C4 = CLBLL_L_X4Y113_SLICE_X4Y113_AO5;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C5 = CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C6 = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A3 = CLBLM_L_X8Y104_SLICE_X10Y104_BO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A6 = CLBLM_L_X10Y105_SLICE_X12Y105_BO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B3 = CLBLM_R_X7Y106_SLICE_X9Y106_AO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D2 = CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D3 = CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D4 = CLBLM_R_X7Y109_SLICE_X9Y109_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D6 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C1 = CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C2 = CLBLM_L_X10Y105_SLICE_X13Y105_BO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C3 = CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C4 = CLBLM_L_X8Y104_SLICE_X10Y104_BO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C5 = CLBLM_R_X7Y105_SLICE_X8Y105_CO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C6 = CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D1 = CLBLM_R_X7Y106_SLICE_X9Y106_AO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D2 = CLBLM_L_X8Y105_SLICE_X10Y105_BO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C6 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A1 = CLBLM_R_X11Y110_SLICE_X15Y110_DO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A2 = CLBLM_L_X12Y110_SLICE_X16Y110_CO6;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_A6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D6 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B1 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B2 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B3 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B4 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B5 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_B6 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C1 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C2 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C3 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C4 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C5 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_C6 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D1 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D2 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D3 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D4 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D5 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X15Y111_D6 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A2 = CLBLM_R_X11Y110_SLICE_X14Y110_CO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A3 = CLBLM_R_X11Y111_SLICE_X15Y111_AO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A5 = CLBLM_L_X12Y110_SLICE_X16Y110_AO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_A6 = 1'b1;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B1 = CLBLM_R_X11Y110_SLICE_X14Y110_BO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B3 = CLBLM_R_X11Y110_SLICE_X14Y110_AO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_B6 = CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C1 = CLBLM_R_X11Y110_SLICE_X14Y110_AO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C4 = CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C5 = CLBLM_R_X11Y110_SLICE_X14Y110_BO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_C6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D1 = CLBLM_L_X12Y110_SLICE_X16Y110_AO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D3 = CLBLM_R_X11Y111_SLICE_X15Y111_AO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D4 = CLBLM_R_X11Y110_SLICE_X14Y110_CO6;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X11Y111_SLICE_X14Y111_D6 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A1 = CLBLM_L_X10Y106_SLICE_X12Y106_CO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A2 = CLBLM_L_X10Y105_SLICE_X13Y105_DO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B3 = CLBLM_L_X8Y107_SLICE_X11Y107_BO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B4 = CLBLM_L_X8Y106_SLICE_X11Y106_BO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B6 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C1 = CLBLM_L_X8Y106_SLICE_X11Y106_BO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C6 = CLBLM_L_X8Y107_SLICE_X11Y107_BO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A1 = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A2 = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A3 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A4 = 1'b1;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A5 = CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_A6 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B1 = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B2 = CLBLL_L_X4Y114_SLICE_X5Y114_BO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B3 = CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D5 = CLBLM_L_X10Y106_SLICE_X12Y106_CO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B4 = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B5 = CLBLL_L_X4Y114_SLICE_X4Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_B6 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C3 = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C4 = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_C6 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A1 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A4 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A6 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B2 = CLBLM_R_X7Y106_SLICE_X9Y106_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B3 = CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B4 = CLBLM_L_X8Y107_SLICE_X10Y107_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B5 = CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B6 = CLBLM_L_X8Y108_SLICE_X10Y108_AO5;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B1 = CLBLM_L_X8Y107_SLICE_X11Y107_BO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D3 = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D4 = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y114_SLICE_X4Y114_D6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C1 = CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C2 = CLBLM_L_X8Y109_SLICE_X11Y109_AO5;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C3 = CLBLM_L_X8Y107_SLICE_X11Y107_CO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C4 = CLBLM_L_X8Y108_SLICE_X10Y108_AO5;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C5 = CLBLM_R_X7Y106_SLICE_X9Y106_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C6 = CLBLM_L_X8Y107_SLICE_X10Y107_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D1 = CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D2 = CLBLM_L_X8Y109_SLICE_X11Y109_AO5;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D3 = CLBLM_L_X8Y107_SLICE_X11Y107_CO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D4 = CLBLM_L_X8Y108_SLICE_X10Y108_AO5;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D5 = CLBLM_R_X7Y106_SLICE_X9Y106_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D6 = CLBLM_L_X8Y107_SLICE_X10Y107_AO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A1 = CLBLM_R_X5Y114_SLICE_X6Y114_AO5;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A2 = CLBLM_R_X5Y114_SLICE_X6Y114_AO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A3 = CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A4 = CLBLL_L_X4Y114_SLICE_X4Y114_BO5;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A5 = CLBLL_L_X4Y114_SLICE_X5Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_A6 = 1'b1;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_D = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_D = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B2 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B4 = CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_B6 = CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A6 = CLBLM_L_X8Y111_SLICE_X11Y111_BO5;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C2 = CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_C6 = CLBLM_R_X7Y113_SLICE_X8Y113_AO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D1 = CLBLM_R_X5Y114_SLICE_X6Y114_AO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D2 = CLBLL_L_X4Y114_SLICE_X4Y114_AO5;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D3 = CLBLL_L_X4Y114_SLICE_X4Y114_DO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D4 = CLBLL_L_X4Y114_SLICE_X5Y114_CO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D5 = CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  assign CLBLL_L_X4Y114_SLICE_X5Y114_D6 = CLBLL_L_X4Y114_SLICE_X5Y114_BO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_A1 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_A2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_A3 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_A5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_A6 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_B1 = CLBLM_L_X8Y102_SLICE_X10Y102_AO5;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_B2 = CLBLM_R_X7Y102_SLICE_X8Y102_BO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_B3 = CLBLM_R_X7Y102_SLICE_X8Y102_CO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_B4 = CLBLM_R_X7Y103_SLICE_X9Y103_AO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_B5 = CLBLM_R_X7Y102_SLICE_X9Y102_AO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_B6 = CLBLM_R_X7Y102_SLICE_X9Y102_AO5;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_C1 = CLBLM_R_X7Y102_SLICE_X9Y102_AO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_C2 = CLBLM_R_X7Y102_SLICE_X8Y102_CO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_C3 = CLBLM_R_X7Y102_SLICE_X8Y102_BO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_C4 = CLBLM_R_X7Y102_SLICE_X9Y102_AO5;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_C5 = CLBLM_L_X8Y102_SLICE_X10Y102_AO5;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_C6 = CLBLM_R_X7Y103_SLICE_X9Y103_AO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_D1 = CLBLM_R_X7Y103_SLICE_X9Y103_AO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_D2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_D3 = CLBLM_R_X7Y102_SLICE_X8Y102_BO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_D4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_D5 = CLBLM_L_X8Y102_SLICE_X10Y102_AO5;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_D6 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_A1 = CLBLM_L_X8Y102_SLICE_X10Y102_AO5;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_A2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_A3 = CLBLM_R_X7Y102_SLICE_X8Y102_DO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_A4 = CLBLM_R_X7Y102_SLICE_X8Y102_BO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_A6 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_B1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_B2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_B3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_B4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_B5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_B6 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_C1 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_C2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_C3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_C4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_C5 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_C6 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_D1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_D2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_D3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_D4 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_D5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_D6 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D4 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A2 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A3 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A6 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B2 = CLBLM_L_X8Y108_SLICE_X11Y108_DO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B4 = CLBLM_R_X11Y109_SLICE_X14Y109_AO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A2 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A3 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C6 = CLBLM_R_X11Y109_SLICE_X14Y109_AO6;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_A6 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C2 = CLBLM_L_X8Y108_SLICE_X11Y108_DO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B2 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B4 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B5 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D5 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D6 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_B6 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C2 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_C6 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A1 = CLBLM_R_X7Y109_SLICE_X8Y109_AO5;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A2 = CLBLM_L_X8Y107_SLICE_X11Y107_BO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A3 = CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A4 = CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A5 = CLBLM_L_X8Y107_SLICE_X11Y107_DO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A6 = CLBLM_L_X8Y108_SLICE_X10Y108_AO5;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D2 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X4Y115_D6 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B1 = CLBLM_L_X8Y107_SLICE_X10Y107_DO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B2 = CLBLM_L_X8Y109_SLICE_X11Y109_BO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B3 = CLBLM_L_X8Y108_SLICE_X11Y108_CO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B4 = CLBLM_L_X8Y108_SLICE_X11Y108_BO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B5 = CLBLM_L_X8Y109_SLICE_X11Y109_AO5;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B6 = CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C1 = CLBLM_L_X8Y109_SLICE_X10Y109_AO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C2 = CLBLM_L_X8Y110_SLICE_X10Y110_AO5;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C3 = CLBLM_L_X8Y108_SLICE_X10Y108_DO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C4 = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C5 = CLBLM_L_X8Y109_SLICE_X10Y109_DO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C6 = CLBLM_R_X5Y109_SLICE_X7Y109_AO5;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B4 = CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D1 = CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D2 = CLBLM_L_X8Y108_SLICE_X10Y108_AO5;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D3 = CLBLM_L_X8Y107_SLICE_X11Y107_DO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D4 = CLBLM_L_X8Y107_SLICE_X11Y107_BO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D5 = CLBLM_R_X7Y109_SLICE_X8Y109_AO5;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A1 = CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A2 = CLBLM_R_X5Y115_SLICE_X6Y115_AO5;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A3 = CLBLM_R_X5Y114_SLICE_X7Y114_AO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A4 = CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_A6 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D6 = CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B1 = CLBLL_L_X4Y114_SLICE_X5Y114_DO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B2 = CLBLM_R_X5Y114_SLICE_X6Y114_AO5;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B4 = CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B5 = CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_B6 = CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C2 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_C6 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C2 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D1 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D2 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D3 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D4 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D5 = 1'b1;
  assign CLBLL_L_X4Y115_SLICE_X5Y115_D6 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D5 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D6 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A6 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B1 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B2 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B3 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B4 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B5 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B6 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C1 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C2 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C3 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C4 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C5 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C6 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D4 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D1 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D2 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D3 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D4 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D5 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D6 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A1 = CLBLM_R_X5Y102_SLICE_X7Y102_DO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A2 = CLBLM_L_X8Y102_SLICE_X11Y102_BO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A3 = CLBLM_R_X7Y104_SLICE_X8Y104_AO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A4 = CLBLM_R_X7Y102_SLICE_X9Y102_BO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A5 = CLBLM_R_X7Y102_SLICE_X9Y102_CO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A6 = CLBLM_R_X5Y103_SLICE_X6Y103_AO5;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B1 = CLBLM_L_X8Y103_SLICE_X11Y103_AO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B3 = CLBLM_R_X7Y102_SLICE_X8Y102_AO5;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B4 = CLBLM_L_X8Y103_SLICE_X10Y103_AO5;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B6 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D4 = CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C1 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C2 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C3 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C4 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C5 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C6 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D6 = CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D1 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D2 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D3 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D4 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D5 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D6 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B6 = CLBLL_L_X4Y114_SLICE_X4Y114_BO5;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C4 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A1 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A3 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A6 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B3 = CLBLM_R_X11Y109_SLICE_X14Y109_AO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B4 = CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B6 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C1 = CLBLM_R_X7Y107_SLICE_X8Y107_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C2 = CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C5 = CLBLM_L_X10Y111_SLICE_X13Y111_AO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C6 = CLBLM_R_X11Y110_SLICE_X15Y110_DO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D1 = CLBLM_L_X12Y110_SLICE_X17Y110_AO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D6 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A1 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A3 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B1 = CLBLM_L_X8Y108_SLICE_X11Y108_BO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B2 = CLBLM_L_X8Y109_SLICE_X11Y109_BO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B4 = CLBLM_L_X8Y108_SLICE_X10Y108_DO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B5 = CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C1 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C2 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C3 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C4 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D1 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D2 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D3 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D4 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D6 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A3 = CLBLM_L_X8Y103_SLICE_X11Y103_AO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A6 = CLBLM_R_X7Y102_SLICE_X9Y102_CO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B3 = CLBLM_L_X8Y104_SLICE_X11Y104_AO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B5 = CLBLM_R_X7Y104_SLICE_X9Y104_AO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B6 = CLBLM_L_X10Y104_SLICE_X12Y104_AO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C1 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C2 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C3 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C4 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C5 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C6 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D1 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D2 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D3 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D4 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D5 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D6 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A1 = CLBLM_R_X7Y104_SLICE_X8Y104_DO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A2 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A5 = CLBLM_R_X7Y103_SLICE_X8Y103_BO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A6 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B5 = CLBLM_L_X8Y103_SLICE_X11Y103_AO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B6 = CLBLM_R_X7Y102_SLICE_X9Y102_CO6;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_D = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_D = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C1 = CLBLM_R_X7Y103_SLICE_X8Y103_BO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C5 = CLBLM_R_X7Y104_SLICE_X8Y104_DO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D3 = CLBLM_R_X7Y102_SLICE_X9Y102_DO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D5 = CLBLM_R_X5Y102_SLICE_X7Y102_DO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A1 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A3 = CLBLM_R_X11Y111_SLICE_X14Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B1 = CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B3 = CLBLM_R_X11Y111_SLICE_X14Y111_DO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C2 = CLBLM_R_X11Y111_SLICE_X14Y111_AO5;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C4 = CLBLM_R_X11Y111_SLICE_X14Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C5 = CLBLM_R_X11Y111_SLICE_X14Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C6 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D2 = CLBLM_R_X11Y111_SLICE_X14Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D4 = CLBLM_L_X8Y111_SLICE_X11Y111_AO5;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D6 = CLBLM_R_X11Y111_SLICE_X14Y111_AO5;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A1 = CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A3 = CLBLM_L_X8Y109_SLICE_X10Y109_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A4 = CLBLM_L_X10Y110_SLICE_X13Y110_CO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A6 = CLBLM_L_X8Y109_SLICE_X11Y109_CO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B1 = CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B2 = CLBLM_L_X8Y108_SLICE_X11Y108_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B3 = CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B4 = CLBLM_L_X10Y110_SLICE_X13Y110_CO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B5 = CLBLM_L_X8Y109_SLICE_X11Y109_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B6 = CLBLM_L_X8Y109_SLICE_X11Y109_CO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C1 = CLBLM_L_X8Y109_SLICE_X11Y109_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C2 = CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C3 = CLBLM_L_X8Y108_SLICE_X11Y108_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C4 = CLBLM_L_X8Y108_SLICE_X10Y108_DO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D1 = CLBLM_L_X8Y109_SLICE_X10Y109_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D4 = CLBLM_L_X10Y110_SLICE_X13Y110_CO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D5 = CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D6 = CLBLM_L_X8Y109_SLICE_X11Y109_CO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B3 = CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B5 = CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B6 = CLBLL_L_X4Y110_SLICE_X4Y110_AO5;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D5 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A2 = CLBLM_L_X8Y104_SLICE_X10Y104_CO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A4 = CLBLM_R_X7Y104_SLICE_X8Y104_CO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A6 = CLBLM_R_X7Y104_SLICE_X9Y104_BO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D6 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B1 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B2 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B3 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B4 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B5 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B6 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C1 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C2 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C3 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C4 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C5 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C6 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D1 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D2 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D3 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D4 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D5 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D6 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A2 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A4 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A6 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B1 = CLBLM_R_X7Y104_SLICE_X8Y104_DO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B2 = CLBLM_L_X8Y103_SLICE_X10Y103_BO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B3 = CLBLM_L_X8Y105_SLICE_X10Y105_AO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B4 = CLBLM_R_X7Y104_SLICE_X8Y104_BO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B5 = CLBLM_R_X5Y105_SLICE_X6Y105_AO5;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B6 = CLBLM_R_X7Y106_SLICE_X8Y106_AO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C1 = CLBLM_R_X5Y105_SLICE_X6Y105_AO5;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C2 = CLBLM_L_X8Y103_SLICE_X10Y103_BO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C3 = CLBLM_R_X7Y104_SLICE_X8Y104_DO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C4 = CLBLM_R_X7Y106_SLICE_X8Y106_AO5;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C5 = CLBLM_L_X8Y105_SLICE_X10Y105_AO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C6 = CLBLM_R_X7Y104_SLICE_X8Y104_BO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D1 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D2 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D3 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D4 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D5 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C4 = CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C5 = CLBLM_R_X5Y113_SLICE_X7Y113_DO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C6 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A1 = CLBLM_L_X10Y112_SLICE_X12Y112_AO5;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A2 = CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A3 = CLBLM_L_X10Y111_SLICE_X13Y111_AO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A4 = CLBLM_L_X10Y112_SLICE_X12Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A5 = CLBLM_L_X10Y110_SLICE_X13Y110_CO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A6 = CLBLM_L_X8Y109_SLICE_X11Y109_CO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B1 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B2 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B3 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B4 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B5 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C1 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C2 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C3 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C4 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C5 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D1 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D2 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D3 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D4 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D5 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A1 = CLBLM_R_X5Y112_SLICE_X6Y112_AO5;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A2 = CLBLM_L_X8Y113_SLICE_X11Y113_BO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A3 = CLBLM_L_X8Y113_SLICE_X11Y113_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A4 = CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A5 = CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A6 = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B1 = CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B2 = CLBLM_L_X10Y110_SLICE_X12Y110_BO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B3 = CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B4 = CLBLM_R_X5Y111_SLICE_X6Y111_AO5;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B5 = CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B6 = CLBLM_L_X10Y112_SLICE_X12Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C1 = CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C2 = CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D1 = CLBLM_L_X10Y111_SLICE_X12Y111_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D5 = CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B3 = CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_D1 = CLBLL_L_X2Y111_SLICE_X0Y111_AO5;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_T1 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A4 = CLBLM_R_X7Y104_SLICE_X8Y104_CO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A5 = CLBLM_L_X8Y104_SLICE_X10Y104_CO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A6 = CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B1 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B2 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B3 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B4 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B5 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B6 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C1 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C2 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C3 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C4 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C5 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C6 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D1 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D2 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D3 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D4 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D5 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D6 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A1 = CLBLM_R_X5Y104_SLICE_X6Y104_DO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A3 = CLBLM_L_X8Y104_SLICE_X10Y104_CO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A4 = CLBLM_R_X7Y104_SLICE_X8Y104_CO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A6 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B1 = CLBLM_R_X5Y104_SLICE_X6Y104_DO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B2 = CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B3 = CLBLM_R_X7Y105_SLICE_X8Y105_CO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B4 = CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B5 = CLBLM_R_X7Y105_SLICE_X8Y105_BO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B6 = CLBLM_R_X5Y106_SLICE_X6Y106_AO5;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C2 = CLBLM_L_X8Y104_SLICE_X10Y104_CO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C3 = CLBLM_R_X5Y104_SLICE_X6Y104_DO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C4 = CLBLM_R_X7Y106_SLICE_X8Y106_AO5;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C6 = CLBLM_R_X7Y104_SLICE_X8Y104_CO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D2 = CLBLM_L_X8Y104_SLICE_X10Y104_CO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D4 = CLBLM_R_X7Y106_SLICE_X8Y106_AO5;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D5 = CLBLM_R_X5Y104_SLICE_X6Y104_DO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D6 = CLBLM_R_X7Y104_SLICE_X8Y104_CO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A1 = CLBLM_R_X5Y111_SLICE_X6Y111_AO5;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A2 = CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A3 = CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A4 = CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A5 = CLBLM_L_X8Y114_SLICE_X10Y114_AO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_A6 = CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B1 = CLBLM_R_X5Y111_SLICE_X6Y111_AO5;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B2 = CLBLM_L_X10Y113_SLICE_X12Y113_BO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B3 = CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B4 = CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B5 = CLBLM_L_X8Y114_SLICE_X10Y114_AO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_B6 = CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_D = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C1 = CLBLM_L_X10Y112_SLICE_X13Y112_BO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C2 = CLBLM_L_X10Y112_SLICE_X12Y112_CO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C3 = CLBLM_L_X10Y112_SLICE_X13Y112_CO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C4 = CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C5 = CLBLM_R_X5Y111_SLICE_X6Y111_AO5;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_C6 = CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D1 = CLBLM_L_X10Y112_SLICE_X13Y112_DO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D2 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D4 = CLBLM_L_X10Y113_SLICE_X12Y113_AO5;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_L_X8Y113_SLICE_X11Y113_D6 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_D = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_D = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A1 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A2 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A3 = CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_A6 = 1'b1;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B1 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B3 = CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B4 = CLBLM_L_X8Y113_SLICE_X11Y113_CO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_B6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C1 = CLBLM_L_X8Y114_SLICE_X10Y114_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C2 = CLBLM_L_X8Y113_SLICE_X11Y113_CO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C3 = CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C4 = CLBLM_L_X8Y113_SLICE_X10Y113_AO5;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C5 = CLBLM_L_X8Y113_SLICE_X10Y113_DO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_C6 = CLBLM_R_X7Y113_SLICE_X9Y113_AO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A2 = CLBLM_R_X3Y104_SLICE_X2Y104_BO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D1 = CLBLM_L_X10Y111_SLICE_X12Y111_AO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D3 = CLBLM_L_X10Y112_SLICE_X12Y112_DO6;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y113_SLICE_X10Y113_D6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A5 = CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A6 = CLBLL_L_X2Y106_SLICE_X0Y106_AO5;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B2 = CLBLM_R_X3Y107_SLICE_X2Y107_BO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B5 = CLBLL_L_X2Y105_SLICE_X0Y105_AO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C1 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C2 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C3 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C4 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C5 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C6 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D1 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D2 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D3 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D4 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D5 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D6 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B2 = CLBLM_L_X10Y113_SLICE_X12Y113_AO5;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A2 = CLBLM_R_X7Y106_SLICE_X8Y106_DO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A3 = CLBLM_R_X7Y105_SLICE_X9Y105_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A1 = CLBLL_L_X2Y106_SLICE_X0Y106_AO5;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B4 = CLBLM_L_X10Y112_SLICE_X13Y112_DO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A4 = CLBLL_L_X2Y105_SLICE_X1Y105_BO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A5 = CLBLM_R_X3Y104_SLICE_X2Y104_BO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A6 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B2 = CLBLM_R_X7Y106_SLICE_X8Y106_DO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C1 = CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B6 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C2 = CLBLM_R_X7Y106_SLICE_X8Y106_DO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C1 = CLBLL_L_X4Y104_SLICE_X4Y104_AO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C2 = CLBLL_L_X2Y106_SLICE_X0Y106_AO5;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C3 = CLBLM_R_X3Y104_SLICE_X2Y104_AO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C4 = CLBLM_R_X3Y109_SLICE_X3Y109_AO5;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C5 = CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C6 = CLBLM_R_X3Y104_SLICE_X2Y104_BO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D1 = CLBLM_R_X7Y104_SLICE_X8Y104_CO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D6 = CLBLM_L_X8Y104_SLICE_X10Y104_CO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D1 = CLBLM_R_X3Y104_SLICE_X2Y104_BO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D2 = CLBLL_L_X2Y106_SLICE_X0Y106_AO5;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D3 = CLBLM_R_X3Y104_SLICE_X2Y104_AO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D4 = CLBLM_R_X3Y109_SLICE_X3Y109_AO5;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D5 = CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D6 = CLBLL_L_X4Y104_SLICE_X4Y104_AO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A2 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A5 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A6 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B3 = CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B4 = CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C4 = CLBLM_L_X8Y114_SLICE_X10Y114_AO5;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C5 = CLBLM_R_X7Y113_SLICE_X9Y113_BO5;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C1 = CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C2 = CLBLM_R_X7Y107_SLICE_X9Y107_AO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C3 = CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C4 = CLBLM_R_X7Y107_SLICE_X8Y107_AO5;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C5 = CLBLM_R_X7Y107_SLICE_X8Y107_DO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C6 = CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C6 = CLBLM_L_X10Y112_SLICE_X13Y112_CO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D1 = CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D5 = CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D2 = CLBLM_L_X10Y112_SLICE_X13Y112_DO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D3 = CLBLM_L_X8Y110_SLICE_X11Y110_AO5;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A2 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A3 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A4 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A5 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_A6 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B2 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B3 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B4 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B5 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_B6 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C2 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C3 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C4 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C5 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_C6 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D2 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D3 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D4 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D5 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X11Y114_D6 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A4 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A5 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_A6 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B2 = CLBLM_L_X8Y114_SLICE_X10Y114_CO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B4 = CLBLM_L_X8Y113_SLICE_X11Y113_DO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_B6 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C4 = CLBLM_R_X5Y113_SLICE_X7Y113_AO5;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C1 = CLBLM_R_X7Y113_SLICE_X9Y113_BO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C5 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C3 = CLBLM_L_X10Y112_SLICE_X12Y112_CO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C4 = CLBLM_L_X10Y112_SLICE_X13Y112_CO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_C6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A6 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C6 = CLBLM_R_X5Y115_SLICE_X7Y115_BO6;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D1 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D2 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D3 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D4 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D5 = 1'b1;
  assign CLBLM_L_X8Y114_SLICE_X10Y114_D6 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B1 = CLBLL_L_X2Y107_SLICE_X0Y107_AO5;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B5 = CLBLL_L_X2Y105_SLICE_X1Y105_AO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C4 = CLBLL_L_X2Y105_SLICE_X0Y105_AO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C6 = CLBLM_R_X3Y107_SLICE_X2Y107_BO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D1 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D2 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D3 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D4 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D5 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D6 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A1 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A3 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A5 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A6 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A3 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C6 = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A6 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B3 = CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B5 = CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B1 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B3 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B6 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C3 = CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C5 = CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D2 = CLBLM_L_X8Y106_SLICE_X11Y106_AO5;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D3 = CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D1 = CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D2 = CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D3 = CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D4 = CLBLL_L_X2Y106_SLICE_X1Y106_AO5;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D5 = CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D6 = CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D1 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D2 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D3 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D4 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D6 = CLBLM_L_X10Y106_SLICE_X13Y106_BO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A1 = CLBLM_R_X7Y107_SLICE_X8Y107_AO5;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A2 = CLBLM_R_X5Y107_SLICE_X6Y107_AO5;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A3 = CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A4 = CLBLM_R_X7Y106_SLICE_X8Y106_BO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A5 = CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A6 = CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B1 = CLBLM_L_X8Y108_SLICE_X10Y108_CO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B4 = CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B5 = CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C1 = CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C2 = CLBLM_R_X7Y107_SLICE_X8Y107_AO5;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C3 = CLBLM_R_X7Y106_SLICE_X8Y106_BO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C4 = CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C5 = CLBLM_R_X5Y107_SLICE_X6Y107_AO5;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C6 = CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D1 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D2 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D3 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D4 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D5 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D6 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = CLBLL_L_X2Y110_SLICE_X0Y110_BO6;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B4 = CLBLM_L_X8Y105_SLICE_X10Y105_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C4 = CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C5 = CLBLM_R_X5Y116_SLICE_X6Y116_AO5;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C6 = CLBLM_R_X7Y115_SLICE_X8Y115_BO5;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A1 = CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A3 = CLBLL_L_X2Y107_SLICE_X1Y107_AO5;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A4 = CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A6 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B3 = CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B4 = CLBLL_L_X2Y108_SLICE_X0Y108_AO5;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B6 = CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C1 = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C5 = CLBLL_L_X2Y108_SLICE_X0Y108_BO5;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C6 = CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D2 = CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D4 = CLBLL_L_X2Y107_SLICE_X0Y107_CO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D6 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A6 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A2 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B1 = CLBLL_L_X2Y107_SLICE_X1Y107_DO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B4 = CLBLL_L_X2Y107_SLICE_X0Y107_DO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B1 = CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B2 = CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B3 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B4 = CLBLM_R_X7Y109_SLICE_X8Y109_BO5;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B5 = CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B6 = CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B6 = CLBLL_L_X2Y107_SLICE_X1Y107_CO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C2 = CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C3 = CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C1 = CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C2 = CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C3 = CLBLM_R_X7Y109_SLICE_X8Y109_BO5;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C4 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C5 = CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C6 = CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D1 = CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D2 = CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D3 = CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D1 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D3 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D5 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D6 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A1 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A5 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A6 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B1 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B5 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B6 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C1 = CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C2 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C3 = CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C4 = CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C5 = CLBLM_R_X7Y109_SLICE_X8Y109_BO5;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C6 = CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D1 = CLBLM_R_X7Y104_SLICE_X8Y104_AO5;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D3 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D6 = CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B2 = CLBLL_L_X2Y108_SLICE_X0Y108_AO5;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B3 = CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B4 = CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C5 = CLBLL_L_X2Y108_SLICE_X0Y108_DO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C6 = CLBLL_L_X2Y107_SLICE_X0Y107_BO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D1 = CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D2 = CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D3 = CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D4 = CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D5 = CLBLM_R_X3Y108_SLICE_X2Y108_AO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D6 = CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B2 = CLBLM_R_X3Y106_SLICE_X2Y106_AO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A4 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A5 = CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B6 = CLBLL_L_X2Y108_SLICE_X1Y108_CO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A2 = CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C3 = CLBLL_L_X2Y107_SLICE_X1Y107_DO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C5 = CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D1 = CLBLM_R_X3Y108_SLICE_X2Y108_BO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D2 = CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D3 = CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D4 = CLBLL_L_X2Y108_SLICE_X1Y108_AO5;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D5 = CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D6 = CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C6 = CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D4 = CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D6 = CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A1 = CLBLM_R_X7Y111_SLICE_X9Y111_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A2 = CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A6 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B1 = CLBLM_R_X7Y111_SLICE_X9Y111_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B2 = CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B6 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C1 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C2 = CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C6 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D3 = CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D4 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D5 = CLBLM_R_X7Y111_SLICE_X9Y111_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D6 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = CLBLL_L_X2Y110_SLICE_X0Y110_BO5;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = CLBLL_L_X2Y109_SLICE_X0Y109_DO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A2 = CLBLL_L_X2Y107_SLICE_X1Y107_BO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A4 = CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A6 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B3 = CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B4 = CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B6 = CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D2 = CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D6 = CLBLL_L_X2Y107_SLICE_X0Y107_CO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = CLBLL_L_X2Y110_SLICE_X0Y110_CO5;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A4 = CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A5 = CLBLM_R_X3Y108_SLICE_X2Y108_BO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A6 = CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A1 = CLBLM_L_X8Y111_SLICE_X11Y111_DO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A5 = CLBLM_L_X8Y111_SLICE_X11Y111_BO5;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B5 = CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B6 = CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B1 = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B2 = CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C1 = CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C2 = CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C3 = CLBLM_R_X11Y111_SLICE_X14Y111_DO6;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_A4 = CLBLM_R_X5Y102_SLICE_X7Y102_AO5;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_A5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_A6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C6 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D2 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_B1 = 1'b1;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_B2 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D6 = CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_B3 = 1'b1;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_B4 = 1'b1;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_B6 = 1'b1;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_C1 = 1'b1;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_C2 = 1'b1;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_C3 = 1'b1;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_C4 = 1'b1;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_C5 = 1'b1;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_C6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A2 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A5 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A6 = 1'b1;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_D1 = 1'b1;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_D2 = 1'b1;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_D3 = 1'b1;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_D4 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B6 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_D5 = 1'b1;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_D6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B1 = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C1 = CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C2 = CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C3 = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C4 = CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C5 = CLBLM_R_X7Y109_SLICE_X8Y109_BO5;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C6 = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_A1 = CLBLM_R_X5Y102_SLICE_X6Y102_AO5;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_A3 = CLBLM_R_X5Y102_SLICE_X7Y102_AO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_A5 = 1'b1;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_A6 = 1'b1;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_B1 = CLBLM_R_X5Y102_SLICE_X6Y102_AO5;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_B2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_B3 = CLBLM_R_X5Y102_SLICE_X7Y102_AO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_B4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_B5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_B6 = CLBLM_R_X5Y102_SLICE_X6Y102_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D1 = CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_C1 = CLBLM_R_X5Y101_SLICE_X6Y101_AO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_C2 = CLBLM_R_X5Y101_SLICE_X7Y101_AO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_C3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_C4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_C5 = CLBLM_R_X5Y102_SLICE_X7Y102_CO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_C6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_D1 = 1'b1;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_D2 = 1'b1;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_D3 = 1'b1;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_D4 = 1'b1;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_D5 = 1'b1;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_D6 = 1'b1;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_D = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_D = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D = LIOB33_X0Y107_IOB_X0Y107_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B1 = CLBLL_L_X2Y110_SLICE_X0Y110_DO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B4 = CLBLL_L_X2Y109_SLICE_X1Y109_AO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C1 = CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C2 = CLBLL_L_X2Y110_SLICE_X1Y110_AO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C5 = CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D3 = CLBLL_L_X2Y108_SLICE_X0Y108_BO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D4 = CLBLL_L_X2Y110_SLICE_X0Y110_CO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D6 = CLBLL_L_X2Y107_SLICE_X0Y107_BO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C6 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A1 = CLBLM_L_X8Y111_SLICE_X11Y111_DO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A4 = CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B3 = CLBLM_L_X8Y111_SLICE_X11Y111_DO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B4 = CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B6 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B1 = CLBLM_L_X8Y111_SLICE_X11Y111_BO5;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D1 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C2 = CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D6 = 1'b1;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_A2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_A4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_A5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_A6 = 1'b1;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_B1 = CLBLM_R_X7Y102_SLICE_X8Y102_BO5;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_B2 = CLBLL_L_X4Y104_SLICE_X4Y104_AO5;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_B3 = CLBLM_R_X5Y102_SLICE_X7Y102_AO5;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D6 = 1'b1;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_B4 = CLBLM_R_X7Y102_SLICE_X8Y102_DO6;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_B5 = CLBLM_R_X7Y102_SLICE_X9Y102_AO6;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_B6 = CLBLM_R_X7Y102_SLICE_X8Y102_CO5;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_C1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_C2 = CLBLM_R_X7Y102_SLICE_X8Y102_DO6;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_C3 = CLBLM_R_X7Y102_SLICE_X8Y102_BO5;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_C4 = CLBLM_R_X5Y102_SLICE_X7Y102_AO5;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_C5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_C6 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A4 = CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A6 = CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_D1 = CLBLM_R_X7Y102_SLICE_X9Y102_AO6;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_D2 = CLBLM_R_X7Y102_SLICE_X8Y102_BO5;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_D3 = CLBLM_R_X7Y102_SLICE_X8Y102_CO5;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_D4 = CLBLM_R_X5Y102_SLICE_X7Y102_AO5;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_D5 = CLBLM_R_X7Y102_SLICE_X8Y102_DO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B6 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_D6 = CLBLL_L_X4Y104_SLICE_X4Y104_AO5;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B2 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C4 = CLBLM_L_X10Y112_SLICE_X13Y112_CO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_A1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_A2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_A3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C6 = CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_A6 = 1'b1;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_B1 = CLBLM_R_X3Y104_SLICE_X3Y104_AO6;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_B2 = CLBLM_R_X5Y101_SLICE_X6Y101_AO5;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_B3 = CLBLM_R_X5Y102_SLICE_X7Y102_AO6;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_B4 = CLBLL_L_X4Y104_SLICE_X4Y104_AO5;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_B5 = CLBLM_R_X5Y102_SLICE_X6Y102_CO6;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_B6 = CLBLM_R_X5Y102_SLICE_X6Y102_AO5;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_C1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_C2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_C3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_C4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_C5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_C6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_D1 = CLBLM_R_X5Y102_SLICE_X6Y102_CO6;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_D2 = CLBLM_R_X5Y101_SLICE_X6Y101_AO5;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_D3 = CLBLM_R_X5Y102_SLICE_X7Y102_AO6;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_D4 = CLBLM_R_X5Y102_SLICE_X6Y102_AO5;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_D5 = CLBLM_R_X3Y104_SLICE_X3Y104_AO6;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_D6 = CLBLL_L_X4Y104_SLICE_X4Y104_AO5;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D5 = CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D6 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A6 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B4 = CLBLM_R_X3Y106_SLICE_X3Y106_AO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B5 = CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C1 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C6 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D6 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A1 = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A2 = CLBLM_R_X3Y109_SLICE_X2Y109_BO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A6 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B2 = CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B5 = CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C6 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A1 = CLBLM_L_X8Y113_SLICE_X10Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A2 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A4 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_A6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D1 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D2 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D4 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D6 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B1 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_A2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_A3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_A4 = CLBLM_R_X7Y102_SLICE_X9Y102_DO6;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_A5 = CLBLM_R_X7Y102_SLICE_X8Y102_AO6;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_A6 = CLBLM_R_X5Y101_SLICE_X7Y101_AO5;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C1 = CLBLM_R_X7Y114_SLICE_X9Y114_AO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C2 = CLBLM_L_X10Y113_SLICE_X12Y113_CO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_C3 = CLBLM_L_X10Y112_SLICE_X12Y112_CO6;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_B1 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_B2 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_B3 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_B4 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_B5 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_B6 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D2 = CLBLM_L_X10Y105_SLICE_X13Y105_DO6;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_C1 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_C2 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_C3 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_C4 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_C5 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_C6 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D6 = CLBLM_L_X10Y113_SLICE_X12Y113_AO5;
  assign CLBLM_R_X7Y113_SLICE_X9Y113_D4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A1 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A2 = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A4 = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_A6 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_D1 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_D2 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_D3 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_D4 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_D5 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_D6 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B4 = CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_B5 = CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_A1 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_A3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_A4 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_A5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_A6 = 1'b1;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C2 = CLBLM_L_X8Y113_SLICE_X10Y113_AO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_C3 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_B1 = CLBLM_R_X5Y102_SLICE_X6Y102_DO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_B2 = CLBLM_R_X5Y102_SLICE_X7Y102_BO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_B3 = CLBLM_R_X7Y102_SLICE_X9Y102_BO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_B4 = CLBLM_R_X5Y102_SLICE_X7Y102_DO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_B5 = CLBLM_R_X5Y103_SLICE_X6Y103_AO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_B6 = CLBLM_R_X5Y103_SLICE_X6Y103_AO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D2 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_C1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_C2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_C3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_C4 = CLBLM_R_X5Y102_SLICE_X7Y102_CO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_C5 = CLBLM_R_X5Y102_SLICE_X6Y102_DO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_C6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D4 = CLBLM_R_X7Y111_SLICE_X8Y111_AO5;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D5 = CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  assign CLBLM_R_X7Y113_SLICE_X8Y113_D6 = CLBLM_R_X7Y113_SLICE_X8Y113_BO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_D1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_D2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_D3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_D4 = CLBLM_R_X5Y102_SLICE_X7Y102_CO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_D5 = CLBLM_R_X5Y102_SLICE_X6Y102_DO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_D6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C1 = CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C3 = CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_D = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_D = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D4 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A2 = CLBLM_L_X10Y112_SLICE_X12Y112_CO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A3 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A5 = CLBLM_L_X10Y112_SLICE_X13Y112_CO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_A6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B1 = CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B5 = CLBLM_R_X7Y114_SLICE_X9Y114_CO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_B6 = CLBLM_R_X7Y114_SLICE_X9Y114_AO5;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A1 = CLBLM_R_X5Y103_SLICE_X6Y103_DO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A5 = CLBLM_R_X5Y103_SLICE_X7Y103_AO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C2 = CLBLM_L_X10Y112_SLICE_X12Y112_CO6;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_C3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B1 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B2 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B3 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B4 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B5 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D2 = CLBLM_R_X7Y113_SLICE_X9Y113_CO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C1 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C2 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C3 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C4 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C5 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y114_SLICE_X9Y114_D4 = CLBLM_R_X7Y114_SLICE_X9Y114_AO5;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A2 = CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_A6 = CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D1 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D2 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D3 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D4 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D5 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D6 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B4 = CLBLM_L_X8Y113_SLICE_X10Y113_CO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B2 = CLBLM_R_X7Y114_SLICE_X9Y114_BO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_B3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A1 = CLBLM_R_X5Y103_SLICE_X6Y103_DO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C1 = CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A2 = CLBLM_R_X7Y103_SLICE_X8Y103_AO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A3 = CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A4 = CLBLM_R_X5Y104_SLICE_X6Y104_BO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A5 = CLBLM_R_X5Y105_SLICE_X6Y105_AO5;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A6 = CLBLM_R_X7Y105_SLICE_X8Y105_AO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B5 = CLBLM_R_X7Y102_SLICE_X9Y102_DO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B6 = CLBLM_R_X5Y102_SLICE_X7Y102_DO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D1 = CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C2 = CLBLM_R_X7Y103_SLICE_X8Y103_AO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C3 = CLBLM_R_X5Y103_SLICE_X6Y103_DO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C6 = CLBLM_R_X5Y104_SLICE_X6Y104_BO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D5 = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_D6 = CLBLM_R_X7Y111_SLICE_X9Y111_AO5;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D1 = CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D2 = CLBLM_R_X7Y103_SLICE_X8Y103_AO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D3 = CLBLM_R_X5Y103_SLICE_X6Y103_DO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D4 = CLBLM_R_X7Y105_SLICE_X8Y105_AO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D5 = CLBLM_R_X5Y105_SLICE_X6Y105_AO5;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D6 = CLBLM_R_X5Y104_SLICE_X6Y104_BO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_D1 = CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A3 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B3 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B6 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A1 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A2 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A3 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A4 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A5 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C3 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B1 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B2 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B3 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B4 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B5 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D2 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C1 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C2 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C3 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C4 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C5 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D3 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A3 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A6 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D1 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D2 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D3 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D4 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D5 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B1 = CLBLM_L_X8Y114_SLICE_X10Y114_BO5;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B2 = CLBLM_L_X8Y114_SLICE_X10Y114_BO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B4 = CLBLM_L_X8Y114_SLICE_X10Y114_CO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A2 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A5 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C3 = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B1 = CLBLM_R_X5Y102_SLICE_X6Y102_DO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B2 = CLBLM_R_X5Y102_SLICE_X7Y102_BO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B3 = CLBLM_R_X5Y103_SLICE_X6Y103_AO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B4 = CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B5 = CLBLM_R_X5Y102_SLICE_X6Y102_BO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B6 = CLBLM_R_X3Y105_SLICE_X3Y105_AO5;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D1 = CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D2 = CLBLM_R_X7Y111_SLICE_X9Y111_AO5;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D3 = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C1 = CLBLM_R_X5Y104_SLICE_X7Y104_AO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C2 = CLBLM_R_X5Y104_SLICE_X6Y104_CO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C6 = CLBLM_R_X5Y105_SLICE_X6Y105_DO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D4 = CLBLM_R_X7Y115_SLICE_X8Y115_AO5;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D5 = CLBLM_L_X8Y114_SLICE_X10Y114_BO5;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D6 = CLBLM_L_X8Y114_SLICE_X10Y114_CO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D1 = CLBLL_L_X4Y104_SLICE_X5Y104_BO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D2 = CLBLM_R_X5Y101_SLICE_X6Y101_CO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_D1 = CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_D1 = CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_T1 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_D1 = CLBLL_L_X2Y111_SLICE_X0Y111_BO5;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1 = CLBLL_L_X2Y111_SLICE_X1Y111_AO5;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1 = CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A1 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A2 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A3 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A4 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A5 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A6 = 1'b1;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_D = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B1 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B2 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B3 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B4 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B5 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B6 = 1'b1;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_D = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_D = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C1 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C2 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C3 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C4 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C5 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C6 = 1'b1;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_D = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D1 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D2 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D3 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D4 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D5 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D6 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A2 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A4 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A6 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B4 = CLBLM_R_X5Y104_SLICE_X6Y104_CO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B6 = CLBLL_L_X4Y104_SLICE_X5Y104_DO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C1 = CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C2 = CLBLM_R_X5Y104_SLICE_X6Y104_AO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C3 = CLBLM_R_X5Y104_SLICE_X6Y104_DO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C4 = CLBLM_R_X5Y106_SLICE_X6Y106_AO5;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C5 = CLBLM_R_X7Y105_SLICE_X8Y105_BO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C6 = CLBLL_L_X4Y104_SLICE_X5Y104_DO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D4 = CLBLM_R_X5Y104_SLICE_X6Y104_CO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D6 = CLBLL_L_X4Y104_SLICE_X5Y104_DO6;
  assign LIOB33_X0Y117_IOB_X0Y118_O = CLBLL_L_X2Y111_SLICE_X0Y111_AO5;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A1 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A2 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A3 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A4 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A5 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A6 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B1 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B2 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B3 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B4 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B5 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B6 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C1 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C2 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C3 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C4 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C5 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C6 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D1 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D2 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D3 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D4 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D5 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D6 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A2 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A5 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A6 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B2 = CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B3 = CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B6 = CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C5 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C1 = CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C2 = CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C3 = CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C4 = CLBLM_R_X5Y107_SLICE_X6Y107_AO5;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C5 = CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C6 = CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C6 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D1 = CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D2 = CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D3 = CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D4 = CLBLM_R_X5Y107_SLICE_X6Y107_AO5;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D5 = CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D6 = CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D6 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_D1 = CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_D1 = CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1 = CLBLL_L_X4Y115_SLICE_X5Y115_AO5;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1 = CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C4 = CLBLM_R_X7Y111_SLICE_X9Y111_AO5;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A1 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A2 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A3 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A4 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A5 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C6 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B1 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B2 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B3 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B4 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B5 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B6 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C1 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C2 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C3 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C4 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C5 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C6 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D2 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D1 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D2 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D3 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D4 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D5 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D6 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D4 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A2 = CLBLM_R_X7Y108_SLICE_X8Y108_CO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A3 = CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A4 = CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A6 = CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B1 = CLBLM_R_X7Y108_SLICE_X8Y108_CO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B2 = CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B3 = CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B4 = CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C1 = CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C2 = CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C3 = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C4 = CLBLM_R_X5Y107_SLICE_X6Y107_CO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C5 = CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C6 = CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D4 = CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D5 = CLBLL_L_X2Y107_SLICE_X1Y107_DO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D6 = CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A6 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B2 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B6 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C2 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C6 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D1 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D2 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D3 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D4 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D5 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D6 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A3 = CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A4 = CLBLM_R_X7Y107_SLICE_X8Y107_CO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B1 = CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B2 = CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B3 = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B4 = CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B5 = CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B6 = CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C3 = CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C4 = CLBLM_R_X7Y107_SLICE_X8Y107_CO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D1 = CLBLM_R_X7Y108_SLICE_X8Y108_CO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D2 = CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D3 = CLBLM_R_X7Y107_SLICE_X9Y107_CO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D4 = CLBLM_R_X5Y107_SLICE_X6Y107_CO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D5 = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D6 = CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A3 = CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A4 = CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_D1 = 1'b0;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B3 = CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B5 = CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C1 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C2 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C3 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C4 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C5 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C6 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_T1 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_D1 = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D1 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D2 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D3 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D4 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D5 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D6 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_T1 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A1 = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A2 = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A3 = CLBLM_L_X8Y104_SLICE_X10Y104_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A4 = CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A5 = CLBLM_L_X10Y110_SLICE_X13Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A6 = CLBLM_R_X7Y104_SLICE_X8Y104_AO5;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B1 = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B3 = CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B4 = CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B6 = CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C1 = CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C2 = CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C3 = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C4 = CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C5 = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C6 = CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D1 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D2 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D3 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D4 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D5 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D6 = 1'b1;
  assign LIOB33_X0Y119_IOB_X0Y120_O = CLBLL_L_X2Y110_SLICE_X0Y110_CO5;
  assign LIOB33_X0Y119_IOB_X0Y119_O = CLBLL_L_X2Y110_SLICE_X0Y110_AO5;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A1 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A2 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A3 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A4 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A5 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A6 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B1 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B2 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B3 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B4 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B5 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B6 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C1 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C2 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C3 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C4 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C5 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C6 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D1 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D2 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D3 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D4 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D5 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D6 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A1 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A3 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A6 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B5 = CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B6 = CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C1 = CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C4 = CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D1 = CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D4 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D6 = CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A2 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A3 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A6 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B2 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B3 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B6 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C2 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C3 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D2 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D3 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D6 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A2 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A6 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B2 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B5 = CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B6 = CLBLM_R_X7Y113_SLICE_X8Y113_AO5;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C5 = CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D2 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_D1 = CLBLM_R_X3Y112_SLICE_X3Y112_BO5;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_T1 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A1 = CLBLM_R_X7Y110_SLICE_X8Y110_AO5;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A2 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A5 = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_A6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B1 = CLBLM_R_X7Y110_SLICE_X8Y110_AO5;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B2 = CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B3 = CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B4 = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B5 = CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_B6 = CLBLM_R_X5Y115_SLICE_X6Y115_CO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = CLBLL_L_X2Y110_SLICE_X0Y110_AO5;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C1 = CLBLM_R_X5Y113_SLICE_X6Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C2 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_C3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B1 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B2 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B3 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B4 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B5 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D1 = CLBLM_R_X5Y114_SLICE_X7Y114_AO5;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D2 = CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C1 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C2 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C3 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C4 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C5 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D3 = CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  assign CLBLM_R_X5Y113_SLICE_X7Y113_D4 = CLBLM_R_X5Y113_SLICE_X7Y113_AO5;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A1 = CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A2 = CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A3 = CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A4 = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A5 = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_A6 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D1 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D2 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D3 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D4 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D5 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B1 = CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B2 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_B5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A1 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A2 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A3 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A4 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A5 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C1 = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C2 = CLBLM_R_X5Y113_SLICE_X6Y113_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C3 = CLBLM_R_X5Y113_SLICE_X7Y113_BO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_C4 = CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B1 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B2 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B3 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B4 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B5 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C1 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C2 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C3 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C4 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C5 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C6 = 1'b1;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D5 = CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  assign CLBLM_R_X5Y113_SLICE_X6Y113_D6 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D1 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D2 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D3 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D4 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D5 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D6 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_C2 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_C3 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_C4 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_C5 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_C6 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A1 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A2 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A3 = CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A4 = CLBLM_R_X7Y114_SLICE_X8Y114_DO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A5 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_A6 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B1 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B2 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B3 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B4 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B5 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_B6 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A2 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A3 = CLBLM_R_X3Y103_SLICE_X3Y103_AO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A6 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C1 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C2 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C3 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D1 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D2 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C1 = CLBLM_R_X3Y103_SLICE_X3Y103_AO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C3 = CLBLM_R_X3Y104_SLICE_X2Y104_BO5;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C5 = CLBLM_R_X5Y102_SLICE_X6Y102_AO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C6 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D3 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_D4 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A2 = CLBLM_R_X7Y113_SLICE_X9Y113_AO5;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A4 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A5 = CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_A6 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D2 = CLBLM_R_X5Y101_SLICE_X6Y101_BO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D4 = CLBLM_R_X3Y104_SLICE_X3Y104_AO5;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D6 = CLBLM_R_X3Y104_SLICE_X2Y104_CO5;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B1 = CLBLL_L_X4Y114_SLICE_X5Y114_CO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B2 = CLBLM_R_X7Y113_SLICE_X9Y113_AO5;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B3 = CLBLM_R_X7Y114_SLICE_X8Y114_AO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B4 = CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_B5 = CLBLM_R_X7Y113_SLICE_X8Y113_CO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A1 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A5 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A6 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C1 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C2 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_C3 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B6 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D1 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D2 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D3 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C2 = CLBLM_R_X5Y102_SLICE_X6Y102_AO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C3 = CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C5 = CLBLM_R_X3Y104_SLICE_X2Y104_BO5;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C6 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D4 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D5 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X6Y114_D6 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D1 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D2 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D3 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D4 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D5 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D6 = 1'b1;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_O = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = CLBLL_L_X4Y114_SLICE_X5Y114_AO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = CLBLL_L_X4Y114_SLICE_X5Y114_AO5;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A4 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_A6 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B1 = CLBLM_R_X5Y115_SLICE_X6Y115_AO5;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B2 = CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B3 = CLBLM_R_X5Y113_SLICE_X7Y113_AO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B4 = CLBLM_R_X7Y115_SLICE_X8Y115_CO5;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B5 = CLBLM_R_X5Y115_SLICE_X7Y115_AO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_B6 = CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A1 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A3 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A6 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C2 = CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_C3 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B1 = CLBLL_L_X2Y105_SLICE_X1Y105_DO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B2 = CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B3 = CLBLM_R_X5Y102_SLICE_X6Y102_BO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B4 = CLBLL_L_X4Y104_SLICE_X4Y104_BO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B5 = CLBLM_R_X3Y105_SLICE_X3Y105_AO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B6 = CLBLM_R_X3Y105_SLICE_X3Y105_AO5;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D1 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D2 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C3 = CLBLM_R_X3Y104_SLICE_X3Y104_CO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C4 = CLBLL_L_X2Y105_SLICE_X1Y105_DO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D3 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X7Y115_D4 = 1'b1;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A1 = CLBLM_R_X7Y115_SLICE_X8Y115_DO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A2 = CLBLM_R_X7Y115_SLICE_X8Y115_CO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A3 = CLBLM_R_X7Y115_SLICE_X8Y115_BO5;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_A6 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D3 = CLBLM_R_X3Y104_SLICE_X3Y104_DO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D4 = CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B1 = CLBLM_L_X8Y114_SLICE_X10Y114_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B2 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B3 = CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_B5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A1 = CLBLM_R_X3Y107_SLICE_X3Y107_BO5;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A2 = CLBLL_L_X4Y104_SLICE_X4Y104_BO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A3 = CLBLM_R_X3Y105_SLICE_X3Y105_AO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A4 = CLBLM_R_X3Y107_SLICE_X2Y107_BO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A5 = CLBLL_L_X2Y105_SLICE_X1Y105_CO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A6 = CLBLL_L_X2Y105_SLICE_X1Y105_DO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C1 = CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C2 = CLBLM_R_X5Y115_SLICE_X7Y115_AO5;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_C3 = CLBLM_R_X7Y115_SLICE_X8Y115_CO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B1 = CLBLL_L_X2Y105_SLICE_X1Y105_AO5;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B3 = CLBLM_R_X3Y104_SLICE_X3Y104_CO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B6 = CLBLM_R_X3Y104_SLICE_X2Y104_CO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D1 = CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D2 = CLBLL_L_X4Y115_SLICE_X5Y115_BO6;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D3 = CLBLM_R_X5Y114_SLICE_X7Y114_AO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C2 = CLBLM_R_X3Y104_SLICE_X3Y104_CO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C4 = CLBLL_L_X2Y105_SLICE_X1Y105_DO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D4 = CLBLM_R_X5Y115_SLICE_X6Y115_AO5;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D5 = CLBLM_R_X5Y116_SLICE_X6Y116_AO5;
  assign CLBLM_R_X5Y115_SLICE_X6Y115_D6 = CLBLM_R_X7Y114_SLICE_X8Y114_CO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D2 = CLBLL_L_X2Y105_SLICE_X0Y105_BO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D5 = CLBLM_R_X3Y105_SLICE_X2Y105_BO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A1 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A2 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A3 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A4 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A5 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B1 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B2 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B3 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B4 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B5 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B6 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C3 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C4 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C5 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C6 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A4 = CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A6 = CLBLM_R_X3Y106_SLICE_X3Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B1 = CLBLM_R_X3Y105_SLICE_X2Y105_DO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B2 = CLBLM_R_X3Y105_SLICE_X3Y105_DO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B3 = CLBLL_L_X4Y105_SLICE_X4Y105_AO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D1 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D5 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D2 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C2 = CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C4 = CLBLL_L_X2Y106_SLICE_X1Y106_DO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A2 = CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A3 = CLBLM_R_X7Y115_SLICE_X8Y115_BO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A5 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A6 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D4 = CLBLM_R_X3Y106_SLICE_X3Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D6 = CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B6 = CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B1 = CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B2 = CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B3 = CLBLM_R_X7Y115_SLICE_X8Y115_BO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B4 = CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B5 = CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A2 = CLBLL_L_X2Y106_SLICE_X1Y106_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C4 = CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C5 = CLBLM_R_X7Y114_SLICE_X9Y114_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C6 = CLBLM_R_X7Y115_SLICE_X8Y115_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A4 = CLBLM_R_X3Y106_SLICE_X2Y106_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A6 = CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C2 = CLBLM_R_X5Y115_SLICE_X6Y115_AO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B2 = CLBLL_L_X2Y105_SLICE_X0Y105_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B5 = CLBLM_R_X3Y105_SLICE_X2Y105_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D1 = CLBLM_R_X5Y115_SLICE_X6Y115_BO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D2 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D3 = CLBLM_R_X7Y114_SLICE_X8Y114_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C2 = CLBLM_R_X3Y105_SLICE_X2Y105_CO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C3 = CLBLL_L_X2Y105_SLICE_X0Y105_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C4 = CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D5 = CLBLM_R_X5Y114_SLICE_X6Y114_BO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D6 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D1 = CLBLL_L_X4Y105_SLICE_X5Y105_AO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D2 = CLBLM_R_X3Y105_SLICE_X2Y105_CO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D3 = CLBLL_L_X2Y106_SLICE_X1Y106_AO5;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D4 = CLBLL_L_X2Y105_SLICE_X0Y105_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D5 = CLBLL_L_X2Y106_SLICE_X1Y106_BO5;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D6 = CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  assign LIOB33_X0Y121_IOB_X0Y122_O = CLBLL_L_X2Y110_SLICE_X0Y110_BO6;
  assign LIOB33_X0Y121_IOB_X0Y121_O = CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A1 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A5 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A6 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B1 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B4 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_D1 = CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_D = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C4 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_T1 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D1 = CLBLL_L_X4Y105_SLICE_X4Y105_AO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D3 = CLBLM_R_X3Y106_SLICE_X2Y106_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_D = LIOB33_X0Y103_IOB_X0Y103_I;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_D1 = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A1 = CLBLL_L_X2Y107_SLICE_X1Y107_AO5;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A2 = CLBLL_L_X2Y105_SLICE_X1Y105_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A6 = CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_T1 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B1 = CLBLM_R_X3Y107_SLICE_X3Y107_AO5;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B2 = CLBLL_L_X2Y107_SLICE_X1Y107_AO5;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B3 = CLBLM_R_X3Y109_SLICE_X3Y109_AO5;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B4 = CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B5 = CLBLL_L_X2Y105_SLICE_X1Y105_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B6 = CLBLM_R_X3Y108_SLICE_X2Y108_AO5;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C1 = CLBLM_R_X3Y108_SLICE_X2Y108_CO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C2 = CLBLL_L_X2Y105_SLICE_X1Y105_CO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C3 = CLBLM_R_X3Y107_SLICE_X3Y107_BO5;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C4 = CLBLM_R_X3Y107_SLICE_X3Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C5 = CLBLM_R_X3Y107_SLICE_X2Y107_DO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C6 = CLBLM_R_X3Y107_SLICE_X2Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D1 = CLBLL_L_X2Y105_SLICE_X1Y105_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D2 = CLBLM_R_X3Y107_SLICE_X3Y107_AO5;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D3 = CLBLL_L_X2Y107_SLICE_X1Y107_AO5;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D4 = CLBLM_R_X3Y109_SLICE_X3Y109_AO5;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D5 = CLBLM_R_X3Y108_SLICE_X2Y108_AO5;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D6 = CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  assign LIOB33_X0Y123_IOB_X0Y124_O = CLBLL_L_X2Y110_SLICE_X0Y110_BO5;
  assign LIOB33_X0Y123_IOB_X0Y123_O = CLBLL_L_X2Y109_SLICE_X0Y109_DO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A3 = CLBLM_R_X3Y106_SLICE_X2Y106_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A4 = CLBLL_L_X2Y108_SLICE_X1Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B3 = CLBLL_L_X4Y107_SLICE_X4Y107_DO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B5 = CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B6 = CLBLM_R_X3Y106_SLICE_X3Y106_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C1 = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C2 = CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C3 = CLBLM_R_X3Y106_SLICE_X3Y106_DO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D1 = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D4 = CLBLM_R_X3Y106_SLICE_X3Y106_DO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D5 = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A1 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A3 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A6 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B5 = CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B6 = CLBLM_R_X3Y108_SLICE_X2Y108_CO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C1 = CLBLM_R_X3Y108_SLICE_X2Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C2 = CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C3 = CLBLL_L_X2Y108_SLICE_X0Y108_AO5;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C4 = CLBLM_R_X3Y108_SLICE_X2Y108_AO5;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C5 = CLBLM_R_X3Y107_SLICE_X3Y107_AO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C6 = CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D1 = CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D4 = CLBLM_R_X3Y108_SLICE_X2Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C1 = CLBLM_R_X11Y105_SLICE_X15Y105_AO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D6 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B3 = CLBLM_R_X7Y105_SLICE_X9Y105_AO6;
  assign LIOB33_X0Y125_IOB_X0Y125_O = CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  assign LIOB33_X0Y125_IOB_X0Y126_O = CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C3 = CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C4 = CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C5 = CLBLM_R_X7Y107_SLICE_X9Y107_DO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C6 = CLBLM_L_X8Y107_SLICE_X10Y107_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A2 = CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B1 = CLBLL_L_X4Y109_SLICE_X4Y109_BO5;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B2 = CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C1 = CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C2 = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D1 = CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D2 = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D4 = CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B2 = CLBLL_L_X4Y106_SLICE_X4Y106_BO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B5 = CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B6 = CLBLM_R_X3Y106_SLICE_X3Y106_AO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_D1 = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_T1 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_D1 = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_T1 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_B3 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_B4 = 1'b1;
  assign LIOB33_X0Y127_IOB_X0Y127_O = CLBLL_L_X2Y111_SLICE_X0Y111_BO5;
  assign LIOB33_X0Y127_IOB_X0Y128_O = CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_B5 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_B6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D3 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D4 = 1'b1;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A1 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A3 = CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A4 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A6 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B1 = CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B5 = CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B6 = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C1 = CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C5 = CLBLL_L_X4Y110_SLICE_X5Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C6 = CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D1 = CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D3 = CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D4 = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D6 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A1 = CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A2 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A3 = CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A6 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B4 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B6 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C1 = CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C2 = CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C5 = CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C5 = CLBLM_R_X7Y113_SLICE_X9Y113_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D1 = CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D4 = CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D6 = CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  assign CLBLM_R_X7Y114_SLICE_X8Y114_C6 = CLBLM_R_X7Y111_SLICE_X9Y111_AO5;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C4 = 1'b1;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C5 = 1'b1;
  assign LIOB33_X0Y129_IOB_X0Y130_O = CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  assign LIOB33_X0Y129_IOB_X0Y129_O = CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  assign CLBLM_R_X5Y114_SLICE_X7Y114_C6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A2 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A3 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B1 = CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B2 = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B3 = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B4 = CLBLL_L_X4Y110_SLICE_X4Y110_BO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B5 = CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B6 = CLBLM_R_X3Y111_SLICE_X3Y111_AO5;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C1 = CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C2 = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C3 = CLBLM_R_X3Y111_SLICE_X2Y111_DO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C4 = CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C5 = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C6 = CLBLL_L_X4Y110_SLICE_X4Y110_BO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D1 = CLBLM_R_X3Y110_SLICE_X3Y110_AO5;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D2 = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D3 = CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D4 = CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D5 = CLBLL_L_X4Y110_SLICE_X4Y110_DO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D6 = CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A2 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A4 = CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A5 = CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B2 = CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B4 = CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C3 = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C4 = CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C6 = CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D1 = CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D2 = CLBLM_R_X3Y110_SLICE_X2Y110_AO5;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D3 = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D4 = CLBLM_R_X3Y109_SLICE_X2Y109_AO5;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D5 = CLBLM_R_X3Y110_SLICE_X2Y110_BO5;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D6 = CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  assign LIOB33_X0Y131_IOB_X0Y132_O = CLBLL_L_X2Y111_SLICE_X1Y111_AO5;
  assign LIOB33_X0Y131_IOB_X0Y131_O = CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_D1 = CLBLM_R_X5Y113_SLICE_X7Y113_CO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_T1 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_D1 = CLBLM_R_X5Y113_SLICE_X6Y113_AO5;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_T1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A3 = CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A4 = CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A6 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B1 = CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B3 = CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B5 = CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B6 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C1 = CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C3 = CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C5 = CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C6 = CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D1 = CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D2 = CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D3 = CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D4 = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D5 = CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D6 = CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A3 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A4 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A6 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B3 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B4 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B6 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C3 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C4 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C6 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D3 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D4 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D6 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A1 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A2 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A3 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A4 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A5 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_A6 = 1'b1;
  assign LIOB33_X0Y133_IOB_X0Y134_O = 1'b0;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B1 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B2 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B3 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B4 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B5 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_B6 = 1'b1;
  assign LIOB33_X0Y133_IOB_X0Y133_O = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C1 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C2 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C3 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C4 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C5 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_C6 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D1 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D2 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D3 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D4 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D5 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X17Y107_D6 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A4 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_A6 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B1 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B2 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B3 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B4 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B5 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_B6 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C1 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C2 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C3 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C4 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C5 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_C6 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D1 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D2 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D3 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D4 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D5 = 1'b1;
  assign CLBLM_L_X12Y107_SLICE_X16Y107_D6 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A4 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A6 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOB33_X0Y135_IOB_X0Y135_O = CLBLM_R_X3Y112_SLICE_X3Y112_BO5;
  assign LIOB33_X0Y135_IOB_X0Y136_O = CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A1 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A2 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A3 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A4 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A5 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_A6 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B1 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B2 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B3 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B4 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B5 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_B6 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C1 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C2 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C3 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C4 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C5 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_C6 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D4 = CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D1 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D3 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D2 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D5 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D6 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D5 = CLBLM_L_X10Y112_SLICE_X13Y112_AO5;
  assign CLBLM_L_X12Y108_SLICE_X17Y108_D4 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D6 = CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_A6 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B5 = CLBLM_L_X12Y108_SLICE_X16Y108_AO6;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_B6 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C1 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C2 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C3 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C4 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C5 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_C6 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D1 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D1 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D2 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D3 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D4 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D5 = 1'b1;
  assign CLBLM_L_X12Y108_SLICE_X16Y108_D6 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D2 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B2 = CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C2 = CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C3 = CLBLM_L_X8Y108_SLICE_X10Y108_CO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C4 = CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign LIOB33_X0Y137_IOB_X0Y138_O = CLBLL_L_X4Y114_SLICE_X4Y114_BO6;
  assign LIOB33_X0Y137_IOB_X0Y137_O = CLBLL_L_X4Y114_SLICE_X4Y114_AO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D5 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D6 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A1 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A2 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A3 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A4 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A5 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_A6 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B1 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B2 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B3 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B4 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B5 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_B6 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C1 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C2 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C3 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C4 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C5 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_C6 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D1 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D2 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D3 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D4 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D5 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X17Y109_D6 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A2 = CLBLM_L_X12Y108_SLICE_X16Y108_AO6;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_A6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B1 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B2 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B3 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B4 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B5 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_B6 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C1 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C2 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C3 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C4 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C5 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_C6 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D1 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D2 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D3 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D4 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D5 = 1'b1;
  assign CLBLM_L_X12Y109_SLICE_X16Y109_D6 = 1'b1;
  assign LIOB33_X0Y139_IOB_X0Y140_O = CLBLL_L_X4Y114_SLICE_X5Y114_AO6;
  assign LIOB33_X0Y139_IOB_X0Y139_O = CLBLL_L_X4Y114_SLICE_X5Y114_AO5;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_B1 = 1'b1;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_B2 = 1'b1;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_B3 = 1'b1;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_B4 = 1'b1;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_B5 = 1'b1;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_B6 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A3 = CLBLM_L_X12Y109_SLICE_X16Y109_AO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_A6 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B1 = CLBLM_L_X12Y110_SLICE_X17Y110_DO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B3 = CLBLM_R_X11Y108_SLICE_X15Y108_BO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B5 = CLBLM_R_X11Y110_SLICE_X15Y110_AO5;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_B6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_C1 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C1 = CLBLM_R_X11Y110_SLICE_X15Y110_AO5;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C4 = CLBLM_R_X11Y108_SLICE_X15Y108_BO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_C2 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C5 = CLBLM_L_X12Y110_SLICE_X17Y110_DO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_C6 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_C3 = 1'b1;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D1 = CLBLM_L_X12Y109_SLICE_X16Y109_AO6;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D2 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X12Y110_SLICE_X17Y110_D6 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A3 = CLBLM_L_X12Y110_SLICE_X17Y110_CO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A4 = CLBLM_L_X12Y110_SLICE_X16Y110_BO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_A6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B5 = CLBLM_L_X12Y109_SLICE_X16Y109_AO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_B6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C2 = CLBLM_L_X12Y110_SLICE_X17Y110_CO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_C6 = CLBLM_L_X12Y110_SLICE_X16Y110_BO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D1 = CLBLM_L_X12Y108_SLICE_X16Y108_AO6;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X12Y110_SLICE_X16Y110_D6 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign LIOB33_X0Y141_IOB_X0Y142_O = CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  assign LIOB33_X0Y141_IOB_X0Y141_O = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_D = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOB33_X0Y143_IOB_X0Y143_O = CLBLL_L_X4Y115_SLICE_X5Y115_AO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A6 = CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C1 = CLBLL_L_X4Y106_SLICE_X5Y106_AO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C2 = CLBLL_L_X4Y107_SLICE_X5Y107_AO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C3 = CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C4 = CLBLL_L_X4Y107_SLICE_X4Y107_AO5;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C5 = CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C6 = CLBLL_L_X4Y107_SLICE_X4Y107_BO5;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1 = CLBLM_R_X5Y113_SLICE_X6Y113_CO6;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B6 = CLBLL_L_X2Y105_SLICE_X0Y105_AO6;
  assign LIOB33_X0Y145_IOB_X0Y146_O = CLBLM_R_X5Y113_SLICE_X6Y113_AO6;
  assign LIOB33_X0Y145_IOB_X0Y145_O = CLBLM_R_X5Y115_SLICE_X7Y115_CO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B1 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A1 = CLBLM_R_X11Y104_SLICE_X14Y104_AO5;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A3 = CLBLM_L_X10Y103_SLICE_X12Y103_CO5;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A4 = CLBLM_L_X10Y103_SLICE_X13Y103_BO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A6 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C4 = CLBLM_L_X10Y107_SLICE_X12Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C5 = CLBLM_R_X11Y107_SLICE_X15Y107_BO5;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C1 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C2 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C3 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C4 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C5 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C6 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C6 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D1 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D2 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D3 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D4 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D5 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D6 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A3 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A5 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A6 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B3 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B5 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B6 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C4 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C5 = RIOB33_X105Y111_IOB_X1Y112_I;
endmodule
