module top(
  input LIOB33_SING_X0Y50_IOB_X0Y50_IPAD,
  input LIOB33_X0Y51_IOB_X0Y51_IPAD,
  input LIOB33_X0Y51_IOB_X0Y52_IPAD,
  input LIOB33_X0Y53_IOB_X0Y53_IPAD,
  input LIOB33_X0Y53_IOB_X0Y54_IPAD,
  input LIOB33_X0Y55_IOB_X0Y55_IPAD,
  input LIOB33_X0Y55_IOB_X0Y56_IPAD,
  input LIOB33_X0Y57_IOB_X0Y57_IPAD,
  input LIOB33_X0Y57_IOB_X0Y58_IPAD,
  input LIOB33_X0Y59_IOB_X0Y59_IPAD,
  input LIOB33_X0Y59_IOB_X0Y60_IPAD,
  input LIOB33_X0Y61_IOB_X0Y61_IPAD,
  input LIOB33_X0Y61_IOB_X0Y62_IPAD,
  input LIOB33_X0Y63_IOB_X0Y63_IPAD,
  input LIOB33_X0Y63_IOB_X0Y64_IPAD,
  input LIOB33_X0Y65_IOB_X0Y65_IPAD,
  input LIOB33_X0Y65_IOB_X0Y66_IPAD,
  input LIOB33_X0Y67_IOB_X0Y67_IPAD,
  input LIOB33_X0Y67_IOB_X0Y68_IPAD,
  input LIOB33_X0Y69_IOB_X0Y69_IPAD,
  input LIOB33_X0Y69_IOB_X0Y70_IPAD,
  input LIOB33_X0Y71_IOB_X0Y71_IPAD,
  input LIOB33_X0Y71_IOB_X0Y72_IPAD,
  input LIOB33_X0Y73_IOB_X0Y73_IPAD,
  input LIOB33_X0Y73_IOB_X0Y74_IPAD,
  input LIOB33_X0Y75_IOB_X0Y75_IPAD,
  input LIOB33_X0Y75_IOB_X0Y76_IPAD,
  input LIOB33_X0Y77_IOB_X0Y77_IPAD,
  input LIOB33_X0Y77_IOB_X0Y78_IPAD,
  input LIOB33_X0Y79_IOB_X0Y79_IPAD,
  input RIOB33_SING_X105Y100_IOB_X1Y100_IPAD,
  input RIOB33_SING_X105Y149_IOB_X1Y149_IPAD,
  input RIOB33_X105Y101_IOB_X1Y101_IPAD,
  input RIOB33_X105Y101_IOB_X1Y102_IPAD,
  input RIOB33_X105Y103_IOB_X1Y103_IPAD,
  input RIOB33_X105Y103_IOB_X1Y104_IPAD,
  input RIOB33_X105Y105_IOB_X1Y105_IPAD,
  input RIOB33_X105Y105_IOB_X1Y106_IPAD,
  input RIOB33_X105Y107_IOB_X1Y107_IPAD,
  input RIOB33_X105Y107_IOB_X1Y108_IPAD,
  input RIOB33_X105Y109_IOB_X1Y109_IPAD,
  input RIOB33_X105Y109_IOB_X1Y110_IPAD,
  input RIOB33_X105Y111_IOB_X1Y111_IPAD,
  input RIOB33_X105Y111_IOB_X1Y112_IPAD,
  input RIOB33_X105Y113_IOB_X1Y113_IPAD,
  input RIOB33_X105Y113_IOB_X1Y114_IPAD,
  input RIOB33_X105Y115_IOB_X1Y115_IPAD,
  input RIOB33_X105Y115_IOB_X1Y116_IPAD,
  input RIOB33_X105Y117_IOB_X1Y117_IPAD,
  input RIOB33_X105Y117_IOB_X1Y118_IPAD,
  input RIOB33_X105Y119_IOB_X1Y119_IPAD,
  input RIOB33_X105Y119_IOB_X1Y120_IPAD,
  input RIOB33_X105Y121_IOB_X1Y121_IPAD,
  input RIOB33_X105Y121_IOB_X1Y122_IPAD,
  input RIOB33_X105Y123_IOB_X1Y123_IPAD,
  input RIOB33_X105Y123_IOB_X1Y124_IPAD,
  input RIOB33_X105Y125_IOB_X1Y125_IPAD,
  input RIOB33_X105Y125_IOB_X1Y126_IPAD,
  input RIOB33_X105Y127_IOB_X1Y127_IPAD,
  input RIOB33_X105Y127_IOB_X1Y128_IPAD,
  input RIOB33_X105Y129_IOB_X1Y129_IPAD,
  input RIOB33_X105Y129_IOB_X1Y130_IPAD,
  input RIOB33_X105Y131_IOB_X1Y131_IPAD,
  input RIOB33_X105Y131_IOB_X1Y132_IPAD,
  input RIOB33_X105Y133_IOB_X1Y133_IPAD,
  input RIOB33_X105Y133_IOB_X1Y134_IPAD,
  input RIOB33_X105Y135_IOB_X1Y135_IPAD,
  input RIOB33_X105Y135_IOB_X1Y136_IPAD,
  input RIOB33_X105Y137_IOB_X1Y137_IPAD,
  input RIOB33_X105Y137_IOB_X1Y138_IPAD,
  input RIOB33_X105Y139_IOB_X1Y139_IPAD,
  input RIOB33_X105Y139_IOB_X1Y140_IPAD,
  input RIOB33_X105Y141_IOB_X1Y141_IPAD,
  input RIOB33_X105Y141_IOB_X1Y142_IPAD,
  input RIOB33_X105Y143_IOB_X1Y143_IPAD,
  input RIOB33_X105Y143_IOB_X1Y144_IPAD,
  input RIOB33_X105Y145_IOB_X1Y145_IPAD,
  input RIOB33_X105Y145_IOB_X1Y146_IPAD,
  input RIOB33_X105Y147_IOB_X1Y147_IPAD,
  input RIOB33_X105Y147_IOB_X1Y148_IPAD,
  output LIOB33_SING_X0Y100_IOB_X0Y100_OPAD,
  output LIOB33_SING_X0Y149_IOB_X0Y149_OPAD,
  output LIOB33_SING_X0Y150_IOB_X0Y150_OPAD,
  output LIOB33_SING_X0Y199_IOB_X0Y199_OPAD,
  output LIOB33_X0Y101_IOB_X0Y101_OPAD,
  output LIOB33_X0Y101_IOB_X0Y102_OPAD,
  output LIOB33_X0Y103_IOB_X0Y103_OPAD,
  output LIOB33_X0Y103_IOB_X0Y104_OPAD,
  output LIOB33_X0Y105_IOB_X0Y105_OPAD,
  output LIOB33_X0Y105_IOB_X0Y106_OPAD,
  output LIOB33_X0Y107_IOB_X0Y107_OPAD,
  output LIOB33_X0Y107_IOB_X0Y108_OPAD,
  output LIOB33_X0Y109_IOB_X0Y109_OPAD,
  output LIOB33_X0Y109_IOB_X0Y110_OPAD,
  output LIOB33_X0Y111_IOB_X0Y111_OPAD,
  output LIOB33_X0Y111_IOB_X0Y112_OPAD,
  output LIOB33_X0Y113_IOB_X0Y113_OPAD,
  output LIOB33_X0Y113_IOB_X0Y114_OPAD,
  output LIOB33_X0Y115_IOB_X0Y115_OPAD,
  output LIOB33_X0Y115_IOB_X0Y116_OPAD,
  output LIOB33_X0Y117_IOB_X0Y117_OPAD,
  output LIOB33_X0Y117_IOB_X0Y118_OPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD,
  output LIOB33_X0Y125_IOB_X0Y125_OPAD,
  output LIOB33_X0Y125_IOB_X0Y126_OPAD,
  output LIOB33_X0Y127_IOB_X0Y127_OPAD,
  output LIOB33_X0Y127_IOB_X0Y128_OPAD,
  output LIOB33_X0Y129_IOB_X0Y129_OPAD,
  output LIOB33_X0Y129_IOB_X0Y130_OPAD,
  output LIOB33_X0Y131_IOB_X0Y131_OPAD,
  output LIOB33_X0Y131_IOB_X0Y132_OPAD,
  output LIOB33_X0Y133_IOB_X0Y133_OPAD,
  output LIOB33_X0Y133_IOB_X0Y134_OPAD,
  output LIOB33_X0Y135_IOB_X0Y135_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output LIOB33_X0Y141_IOB_X0Y141_OPAD,
  output LIOB33_X0Y141_IOB_X0Y142_OPAD,
  output LIOB33_X0Y143_IOB_X0Y143_OPAD,
  output LIOB33_X0Y145_IOB_X0Y145_OPAD,
  output LIOB33_X0Y145_IOB_X0Y146_OPAD,
  output LIOB33_X0Y147_IOB_X0Y147_OPAD,
  output LIOB33_X0Y147_IOB_X0Y148_OPAD,
  output LIOB33_X0Y151_IOB_X0Y151_OPAD,
  output LIOB33_X0Y151_IOB_X0Y152_OPAD,
  output LIOB33_X0Y153_IOB_X0Y153_OPAD,
  output LIOB33_X0Y153_IOB_X0Y154_OPAD,
  output LIOB33_X0Y155_IOB_X0Y155_OPAD,
  output LIOB33_X0Y155_IOB_X0Y156_OPAD,
  output LIOB33_X0Y157_IOB_X0Y157_OPAD,
  output LIOB33_X0Y157_IOB_X0Y158_OPAD,
  output LIOB33_X0Y159_IOB_X0Y159_OPAD,
  output LIOB33_X0Y159_IOB_X0Y160_OPAD,
  output LIOB33_X0Y161_IOB_X0Y161_OPAD,
  output LIOB33_X0Y161_IOB_X0Y162_OPAD,
  output LIOB33_X0Y163_IOB_X0Y163_OPAD,
  output LIOB33_X0Y163_IOB_X0Y164_OPAD,
  output LIOB33_X0Y165_IOB_X0Y165_OPAD,
  output LIOB33_X0Y165_IOB_X0Y166_OPAD,
  output LIOB33_X0Y167_IOB_X0Y167_OPAD,
  output LIOB33_X0Y167_IOB_X0Y168_OPAD,
  output LIOB33_X0Y169_IOB_X0Y169_OPAD,
  output LIOB33_X0Y169_IOB_X0Y170_OPAD,
  output LIOB33_X0Y171_IOB_X0Y171_OPAD,
  output LIOB33_X0Y171_IOB_X0Y172_OPAD,
  output LIOB33_X0Y173_IOB_X0Y173_OPAD,
  output LIOB33_X0Y173_IOB_X0Y174_OPAD,
  output LIOB33_X0Y175_IOB_X0Y175_OPAD,
  output LIOB33_X0Y175_IOB_X0Y176_OPAD,
  output LIOB33_X0Y177_IOB_X0Y177_OPAD,
  output LIOB33_X0Y177_IOB_X0Y178_OPAD,
  output LIOB33_X0Y179_IOB_X0Y179_OPAD,
  output LIOB33_X0Y179_IOB_X0Y180_OPAD,
  output LIOB33_X0Y181_IOB_X0Y181_OPAD,
  output LIOB33_X0Y181_IOB_X0Y182_OPAD,
  output LIOB33_X0Y183_IOB_X0Y183_OPAD,
  output LIOB33_X0Y183_IOB_X0Y184_OPAD,
  output LIOB33_X0Y185_IOB_X0Y185_OPAD,
  output LIOB33_X0Y185_IOB_X0Y186_OPAD,
  output LIOB33_X0Y187_IOB_X0Y187_OPAD,
  output LIOB33_X0Y187_IOB_X0Y188_OPAD,
  output LIOB33_X0Y189_IOB_X0Y189_OPAD,
  output LIOB33_X0Y189_IOB_X0Y190_OPAD,
  output LIOB33_X0Y191_IOB_X0Y191_OPAD,
  output LIOB33_X0Y191_IOB_X0Y192_OPAD,
  output LIOB33_X0Y193_IOB_X0Y193_OPAD,
  output LIOB33_X0Y193_IOB_X0Y194_OPAD,
  output LIOB33_X0Y195_IOB_X0Y195_OPAD,
  output LIOB33_X0Y195_IOB_X0Y196_OPAD,
  output LIOB33_X0Y197_IOB_X0Y197_OPAD,
  output LIOB33_X0Y197_IOB_X0Y198_OPAD,
  output LIOB33_X0Y79_IOB_X0Y80_OPAD,
  output RIOB33_SING_X105Y150_IOB_X1Y150_OPAD,
  output RIOB33_SING_X105Y199_IOB_X1Y199_OPAD,
  output RIOB33_X105Y151_IOB_X1Y151_OPAD,
  output RIOB33_X105Y151_IOB_X1Y152_OPAD,
  output RIOB33_X105Y153_IOB_X1Y153_OPAD,
  output RIOB33_X105Y153_IOB_X1Y154_OPAD,
  output RIOB33_X105Y155_IOB_X1Y155_OPAD,
  output RIOB33_X105Y155_IOB_X1Y156_OPAD,
  output RIOB33_X105Y157_IOB_X1Y157_OPAD,
  output RIOB33_X105Y157_IOB_X1Y158_OPAD,
  output RIOB33_X105Y159_IOB_X1Y159_OPAD,
  output RIOB33_X105Y159_IOB_X1Y160_OPAD,
  output RIOB33_X105Y161_IOB_X1Y161_OPAD,
  output RIOB33_X105Y161_IOB_X1Y162_OPAD,
  output RIOB33_X105Y163_IOB_X1Y163_OPAD,
  output RIOB33_X105Y163_IOB_X1Y164_OPAD,
  output RIOB33_X105Y165_IOB_X1Y165_OPAD,
  output RIOB33_X105Y165_IOB_X1Y166_OPAD,
  output RIOB33_X105Y167_IOB_X1Y167_OPAD,
  output RIOB33_X105Y167_IOB_X1Y168_OPAD,
  output RIOB33_X105Y169_IOB_X1Y169_OPAD,
  output RIOB33_X105Y169_IOB_X1Y170_OPAD,
  output RIOB33_X105Y171_IOB_X1Y171_OPAD,
  output RIOB33_X105Y171_IOB_X1Y172_OPAD,
  output RIOB33_X105Y173_IOB_X1Y173_OPAD,
  output RIOB33_X105Y173_IOB_X1Y174_OPAD,
  output RIOB33_X105Y175_IOB_X1Y175_OPAD,
  output RIOB33_X105Y175_IOB_X1Y176_OPAD,
  output RIOB33_X105Y177_IOB_X1Y177_OPAD,
  output RIOB33_X105Y177_IOB_X1Y178_OPAD,
  output RIOB33_X105Y179_IOB_X1Y179_OPAD,
  output RIOB33_X105Y179_IOB_X1Y180_OPAD,
  output RIOB33_X105Y181_IOB_X1Y181_OPAD,
  output RIOB33_X105Y181_IOB_X1Y182_OPAD,
  output RIOB33_X105Y183_IOB_X1Y183_OPAD,
  output RIOB33_X105Y183_IOB_X1Y184_OPAD,
  output RIOB33_X105Y185_IOB_X1Y185_OPAD,
  output RIOB33_X105Y185_IOB_X1Y186_OPAD,
  output RIOB33_X105Y187_IOB_X1Y187_OPAD,
  output RIOB33_X105Y187_IOB_X1Y188_OPAD,
  output RIOB33_X105Y189_IOB_X1Y189_OPAD,
  output RIOB33_X105Y189_IOB_X1Y190_OPAD,
  output RIOB33_X105Y191_IOB_X1Y191_OPAD,
  output RIOB33_X105Y191_IOB_X1Y192_OPAD,
  output RIOB33_X105Y193_IOB_X1Y193_OPAD,
  output RIOB33_X105Y193_IOB_X1Y194_OPAD,
  output RIOB33_X105Y195_IOB_X1Y195_OPAD,
  output RIOB33_X105Y195_IOB_X1Y196_OPAD,
  output RIOB33_X105Y197_IOB_X1Y197_OPAD,
  output RIOB33_X105Y197_IOB_X1Y198_OPAD
  );
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_AMUX;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_AO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_A_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_BO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_BO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_B_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_CO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_CO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_C_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_DO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_DO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X0Y115_D_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_AO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_A_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_BO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_BO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_B_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_CO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_CO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_C_XOR;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D1;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D2;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D3;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D4;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_DO5;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_DO6;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D_CY;
  wire [0:0] CLBLL_L_X2Y115_SLICE_X1Y115_D_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_AMUX;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_AO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_A_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_BMUX;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_BO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_BO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_B_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_CMUX;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_CO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_C_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_DO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_DO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X0Y117_D_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_AO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_A_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_BO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_BO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_B_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_CO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_CO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_C_XOR;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D1;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D2;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D3;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D4;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_DO5;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_DO6;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D_CY;
  wire [0:0] CLBLL_L_X2Y117_SLICE_X1Y117_D_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_AMUX;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_AO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_A_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_BO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_BO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_B_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_CO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_CO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_C_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_DO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_DO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X0Y118_D_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A5Q;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_AMUX;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_AO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_AO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_AQ;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_A_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B5Q;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_BMUX;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_BO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_BQ;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_BX;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_B_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_CLK;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_CMUX;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_CO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_C_XOR;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D1;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D2;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D3;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D4;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_DO5;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_DO6;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D_CY;
  wire [0:0] CLBLL_L_X2Y118_SLICE_X1Y118_D_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_AO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_A_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_BO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_B_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_CO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_C_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_DMUX;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_DO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_DO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X0Y119_D_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_AO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_AQ;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_A_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_BO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_B_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_CLK;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_CO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_C_XOR;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D1;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D2;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D3;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D4;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_DO5;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_DO6;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D_CY;
  wire [0:0] CLBLL_L_X2Y119_SLICE_X1Y119_D_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_AO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_A_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_BO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_B_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_CO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_C_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_DO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X0Y120_D_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_AO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_AQ;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_A_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_BO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_B_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_CLK;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_CO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_C_XOR;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D1;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D2;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D3;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D4;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_DO5;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D_CY;
  wire [0:0] CLBLL_L_X2Y120_SLICE_X1Y120_D_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A5Q;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_AMUX;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_AO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_AQ;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_AX;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_A_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_BMUX;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_BO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_BQ;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_BX;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_B_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_CLK;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_CO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_CO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_C_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_DO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_DO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X0Y121_D_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_AMUX;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_AO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_A_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B5Q;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_BMUX;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_BO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_BQ;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_B_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_CLK;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_CMUX;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_CO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_C_XOR;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D1;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D2;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D3;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D4;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_DO5;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D_CY;
  wire [0:0] CLBLL_L_X2Y121_SLICE_X1Y121_D_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_AO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_AO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_A_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_BO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_BO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_B_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_CO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_CO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_C_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_DO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_DO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X0Y122_D_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A5Q;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_AMUX;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_AO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_AO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_AQ;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_A_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_BO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_BO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_BQ;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_B_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_CLK;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_CO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_CO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_C_XOR;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D1;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D2;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D3;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D4;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_DO5;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_DO6;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D_CY;
  wire [0:0] CLBLL_L_X2Y122_SLICE_X1Y122_D_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_AO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_AO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_A_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_BO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_BO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_B_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_CO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_CO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_C_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_DO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_DO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X0Y125_D_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_AO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_AO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_AQ;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_A_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_BO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_BO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_BQ;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_B_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_CLK;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_CMUX;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_CO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_CO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_C_XOR;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D1;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D2;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D3;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D4;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_DO5;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_DO6;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D_CY;
  wire [0:0] CLBLL_L_X2Y125_SLICE_X1Y125_D_XOR;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_A;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_A1;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_A2;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_A3;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_A4;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_A5;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_A6;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_AMUX;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_AO5;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_AO6;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_A_CY;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_A_XOR;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_B;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_B1;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_B2;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_B3;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_B4;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_B5;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_B6;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_BO5;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_BO6;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_B_CY;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_B_XOR;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_C;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_C1;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_C2;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_C3;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_C4;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_C5;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_C6;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_CO5;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_CO6;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_C_CY;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_C_XOR;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_D;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_D1;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_D2;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_D3;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_D4;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_D5;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_D6;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_DO5;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_DO6;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_D_CY;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X0Y126_D_XOR;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_A;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_A1;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_A2;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_A3;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_A4;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_A5;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_A6;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_AO5;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_AO6;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_AQ;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_A_CY;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_A_XOR;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_B;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_B1;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_B2;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_B3;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_B4;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_B5;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_B6;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_BO5;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_BO6;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_B_CY;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_B_XOR;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_C;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_C1;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_C2;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_C3;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_C4;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_C5;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_C6;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_CLK;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_CO5;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_CO6;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_C_CY;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_C_XOR;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_D;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_D1;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_D2;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_D3;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_D4;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_D5;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_D6;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_DO5;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_DO6;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_D_CY;
  wire [0:0] CLBLL_L_X2Y126_SLICE_X1Y126_D_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_AO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_AO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_A_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_BMUX;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_BO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_BO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_B_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_CO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_CO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_C_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_DO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_DO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X0Y127_D_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_AO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_AO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_A_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_BO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_BO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_B_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_CO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_CO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_C_XOR;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D1;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D2;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D3;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D4;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_DO5;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_DO6;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D_CY;
  wire [0:0] CLBLL_L_X2Y127_SLICE_X1Y127_D_XOR;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A1;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A2;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A3;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A4;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_AMUX;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_AO5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_AO6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A_CY;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_A_XOR;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B1;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B2;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B3;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B4;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_BMUX;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_BO5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_BO6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B_CY;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_B_XOR;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C1;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C2;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C3;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C4;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_CMUX;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_CO5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_CO6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C_CY;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_C_XOR;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D1;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D2;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D3;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D4;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_DO5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_DO6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D_CY;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X0Y128_D_XOR;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A1;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A2;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A3;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A4;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_AMUX;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_AO5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_AO6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A_CY;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_A_XOR;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B1;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B2;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B3;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B4;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_BMUX;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_BO5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_BO6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B_CY;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_B_XOR;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C1;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C2;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C3;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C4;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_CO5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_CO6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C_CY;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_C_XOR;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D1;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D2;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D3;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D4;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_DO5;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_DO6;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D_CY;
  wire [0:0] CLBLL_L_X2Y128_SLICE_X1Y128_D_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_AMUX;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_AO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_AO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_A_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_BO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_BO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_B_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_CMUX;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_CO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_CO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_C_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_DO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_DO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X0Y129_D_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_AO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_AO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_A_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_BO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_BO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_B_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_CO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_CO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_C_XOR;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D1;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D2;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D3;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D4;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_DO5;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_DO6;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D_CY;
  wire [0:0] CLBLL_L_X2Y129_SLICE_X1Y129_D_XOR;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_A;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_A1;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_A2;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_A3;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_A4;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_A5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_A6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_AMUX;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_AO5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_AO6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_A_CY;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_A_XOR;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_B;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_B1;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_B2;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_B3;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_B4;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_B5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_B6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_BMUX;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_BO5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_BO6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_B_CY;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_B_XOR;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_C;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_C1;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_C2;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_C3;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_C4;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_C5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_C6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_CMUX;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_CO5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_CO6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_C_CY;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_C_XOR;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_D;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_D1;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_D2;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_D3;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_D4;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_D5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_D6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_DMUX;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_DO5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_DO6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_D_CY;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X0Y130_D_XOR;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_A;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_A1;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_A2;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_A3;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_A4;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_A5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_A6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_AMUX;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_AO5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_AO6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_A_CY;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_A_XOR;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_B;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_B1;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_B2;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_B3;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_B4;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_B5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_B6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_BMUX;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_BO5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_BO6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_B_CY;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_B_XOR;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_C;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_C1;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_C2;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_C3;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_C4;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_C5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_C6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_CO5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_CO6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_C_CY;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_C_XOR;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_D;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_D1;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_D2;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_D3;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_D4;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_D5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_D6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_DO5;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_DO6;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_D_CY;
  wire [0:0] CLBLL_L_X2Y130_SLICE_X1Y130_D_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_AO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_AO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_A_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_BO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_BO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_B_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_CO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_CO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_C_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_DO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_DO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X0Y131_D_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_AO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_AO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_A_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_BO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_BO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_B_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_CO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_CO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_C_XOR;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D1;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D2;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D3;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D4;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_DO5;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_DO6;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D_CY;
  wire [0:0] CLBLL_L_X2Y131_SLICE_X1Y131_D_XOR;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A1;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A2;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A3;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A4;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_AO5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_AO6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A_CY;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_A_XOR;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B1;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B2;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B3;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B4;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_BO5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_BO6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B_CY;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_B_XOR;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C1;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C2;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C3;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C4;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_CO5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_CO6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C_CY;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_C_XOR;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D1;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D2;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D3;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D4;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_DO5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_DO6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D_CY;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X0Y132_D_XOR;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A1;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A2;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A3;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A4;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_AO5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_AO6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A_CY;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_A_XOR;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B1;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B2;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B3;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B4;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_BO5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_BO6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B_CY;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_B_XOR;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C1;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C2;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C3;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C4;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_CO5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_CO6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C_CY;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_C_XOR;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D1;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D2;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D3;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D4;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_DO5;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_DO6;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D_CY;
  wire [0:0] CLBLL_L_X2Y132_SLICE_X1Y132_D_XOR;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_A;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_A1;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_A2;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_A3;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_A4;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_A5;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_A6;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_AO5;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_AO6;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_A_CY;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_A_XOR;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_B;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_B1;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_B2;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_B3;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_B4;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_B5;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_B6;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_BO5;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_BO6;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_B_CY;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_B_XOR;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_C;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_C1;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_C2;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_C3;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_C4;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_C5;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_C6;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_CO5;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_CO6;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_C_CY;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_C_XOR;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_D;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_D1;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_D2;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_D3;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_D4;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_D5;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_D6;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_DO5;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_DO6;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_D_CY;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X54Y124_D_XOR;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_A;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_A1;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_A2;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_A3;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_A4;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_A5;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_A6;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_AO5;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_AO6;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_A_CY;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_A_XOR;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_B;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_B1;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_B2;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_B3;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_B4;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_B5;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_B6;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_BO5;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_BO6;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_B_CY;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_B_XOR;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_C;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_C1;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_C2;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_C3;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_C4;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_C5;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_C6;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_CO5;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_CO6;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_C_CY;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_C_XOR;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_D;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_D1;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_D2;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_D3;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_D4;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_D5;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_D6;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_DO5;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_DO6;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_D_CY;
  wire [0:0] CLBLL_L_X36Y124_SLICE_X55Y124_D_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AMUX;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_A_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_BO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_B_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CLK;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_C_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_DO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X4Y117_D_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_AO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_AQ;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_A_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_BO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_BQ;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_B_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CLK;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CMUX;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_C_XOR;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D1;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D2;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D3;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D4;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_DO5;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D_CY;
  wire [0:0] CLBLL_L_X4Y117_SLICE_X5Y117_D_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_AO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_AO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_AQ;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_A_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_BO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_BO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_B_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_CLK;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_CO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_CO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_C_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_DO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_DO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X4Y118_D_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_AO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_AO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_A_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_BO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_BO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_BQ;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_B_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C5Q;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_CLK;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_CMUX;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_CO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_CO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_CQ;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_C_XOR;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D1;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D2;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D3;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D4;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_DO5;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_DO6;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D_CY;
  wire [0:0] CLBLL_L_X4Y118_SLICE_X5Y118_D_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_A_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_BO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_B_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CLK;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_CQ;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_C_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_DO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_DO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_DQ;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X4Y119_D_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_AO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_A_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_BO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_BQ;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_B_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_CLK;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_CO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_CQ;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_C_XOR;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D1;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D2;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D3;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D4;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_DMUX;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_DO5;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_DO6;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D_CY;
  wire [0:0] CLBLL_L_X4Y119_SLICE_X5Y119_D_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A5Q;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AMUX;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AQ;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_AX;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_A_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_BO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_BQ;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_B_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C5Q;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_CLK;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_CMUX;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_CO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_CQ;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_C_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_DO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_DO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_DQ;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X4Y120_D_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A5Q;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AMUX;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AQ;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_AX;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_A_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_BO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_BO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_BQ;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_B_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_CLK;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_CO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_CO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_CQ;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_C_XOR;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D1;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D2;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D3;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D4;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_DO5;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D_CY;
  wire [0:0] CLBLL_L_X4Y120_SLICE_X5Y120_D_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_AO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_AO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_AQ;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_A_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_BO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_BO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_BQ;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_B_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_CLK;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_CO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_CQ;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_C_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_DO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_DO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_DQ;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X4Y121_D_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_AO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_AO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_AQ;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_A_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_BO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_BO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_BQ;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_B_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_CLK;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_CO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_CO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_CQ;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_C_XOR;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D1;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D2;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D3;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D4;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_DO5;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_DO6;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D_CY;
  wire [0:0] CLBLL_L_X4Y121_SLICE_X5Y121_D_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A5Q;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_AMUX;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_AO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_AO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_AQ;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_AX;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_A_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_BO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_BO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_BQ;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_B_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_CLK;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_CMUX;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_CO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_CO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_C_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_DO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_DO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_DQ;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X4Y122_D_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_AO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_AO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_AQ;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_A_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_BO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_BO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_BQ;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_B_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C5Q;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_CLK;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_CMUX;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_CO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_CO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_CQ;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_C_XOR;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D1;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D2;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D3;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D4;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_DO5;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_DO6;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_DQ;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D_CY;
  wire [0:0] CLBLL_L_X4Y122_SLICE_X5Y122_D_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_AO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_AO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_AQ;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_A_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_BO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_BO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_BQ;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_B_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_CLK;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_CO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_CO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_C_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_DO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_DO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X4Y123_D_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_AO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_AO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_AQ;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_A_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B5Q;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_BMUX;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_BO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_BO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_BQ;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_B_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_CLK;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_CMUX;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_CO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_CO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_C_XOR;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D1;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D2;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D3;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D4;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_DO5;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_DO6;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D_CY;
  wire [0:0] CLBLL_L_X4Y123_SLICE_X5Y123_D_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A5Q;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_AMUX;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_AO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_AO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_AQ;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_AX;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_A_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_BO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_BO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_BQ;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_B_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_CLK;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_CO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_CO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_CQ;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_C_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_DO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_DO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_DQ;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X4Y124_D_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_AO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_AO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_A_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_BO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_BO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_BQ;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_B_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_CLK;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_CO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_CO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_CQ;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_C_XOR;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D1;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D2;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D3;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D4;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_DO5;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_DO6;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_DQ;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D_CY;
  wire [0:0] CLBLL_L_X4Y124_SLICE_X5Y124_D_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_AO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_AO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_AQ;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_A_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_BO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_BO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_BQ;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_B_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C5Q;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_CLK;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_CMUX;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_CO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_CO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_CQ;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_C_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_DO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_DO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X4Y125_D_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_AO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_AO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_AQ;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_A_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_BO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_BO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_BQ;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_B_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_CLK;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_CO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_CO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_C_XOR;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D1;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D2;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D3;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D4;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_DO5;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_DO6;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D_CY;
  wire [0:0] CLBLL_L_X4Y125_SLICE_X5Y125_D_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_AO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_AO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_AQ;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_A_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_BMUX;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_BO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_BO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_B_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_CLK;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_CMUX;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_CO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_CO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_C_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_DO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X4Y126_D_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_AO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_AO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_A_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_BO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_BO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_B_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_CO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_CO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_C_XOR;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D1;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D2;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D3;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D4;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_DO5;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_DO6;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D_CY;
  wire [0:0] CLBLL_L_X4Y126_SLICE_X5Y126_D_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_AMUX;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_AO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_AO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_A_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_BO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_BO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_B_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_CMUX;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_CO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_CO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_C_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_DO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_DO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X4Y127_D_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_AO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_AO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_A_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_BO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_BO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_B_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_CMUX;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_CO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_CO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_C_XOR;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D1;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D2;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D3;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D4;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_DO5;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_DO6;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D_CY;
  wire [0:0] CLBLL_L_X4Y127_SLICE_X5Y127_D_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_AO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_AO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_A_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_BO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_BO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_B_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_CO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_CO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_C_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_DO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_DO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X4Y128_D_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_AO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_AO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_A_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_BO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_BO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_B_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_CMUX;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_CO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_CO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_C_XOR;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D1;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D2;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D3;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D4;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_DO5;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_DO6;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D_CY;
  wire [0:0] CLBLL_L_X4Y128_SLICE_X5Y128_D_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_AO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_AO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_AQ;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_BMUX;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_BO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_BO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_CLK;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_CO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_CO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_DO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_DO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_AO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_AO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_AQ;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_BO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_BO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_CLK;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_CO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_CO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_DO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_DO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_AMUX;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_AO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_AO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_BO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_BO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_CO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_CO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_DO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_DO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_AO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_AO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_BO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_BO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_CO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_CO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_DO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_DO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_AO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_AO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_BO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_CO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_CO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_DO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_DO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_AO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_AO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_BO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_BO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_CO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_CO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_DO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_DO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_AO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_BO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_BO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_CO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_CO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_DO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_DO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_AO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_AO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_BO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_BO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_CO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_CO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_DO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_DO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_AO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_AO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_A_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_BO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_BO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_B_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_CLK;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_CO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_CO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_C_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_DO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_DO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X12Y117_D_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_AO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_AO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_A_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_BO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_B_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_CO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_C_XOR;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D1;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D2;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D3;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D4;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_DO5;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D_CY;
  wire [0:0] CLBLM_L_X10Y117_SLICE_X13Y117_D_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_AO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_AO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_A_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_BO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_BO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_B_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_CLK;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_CO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_CO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_C_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_DO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_DO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X12Y118_D_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_AO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_AO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_AQ;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_A_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_BO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_BO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_B_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_CLK;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_CO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_C_XOR;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D1;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D2;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D3;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D4;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_DO5;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_DO6;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D_CY;
  wire [0:0] CLBLM_L_X10Y118_SLICE_X13Y118_D_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_AO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_AO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_A_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_BO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_BQ;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_B_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_CLK;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_CO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_CO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_CQ;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_C_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_DO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_DO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_DQ;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X12Y119_D_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_AO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_AO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_A_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_BO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_BO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_BQ;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_B_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_CLK;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_CO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_CO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_C_XOR;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D1;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D2;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D3;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D4;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_DO5;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_DO6;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D_CY;
  wire [0:0] CLBLM_L_X10Y119_SLICE_X13Y119_D_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_AO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_AQ;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_A_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_BO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_BQ;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_B_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_CLK;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_CO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_CQ;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_C_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_DO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X12Y120_D_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A5Q;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_AMUX;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_AO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_AO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_AQ;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_A_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_BMUX;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_BO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_BO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_BQ;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_B_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_CLK;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_CO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_CO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_CQ;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_C_XOR;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D1;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D2;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D3;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D4;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_DO5;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_DO6;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D_CY;
  wire [0:0] CLBLM_L_X10Y120_SLICE_X13Y120_D_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_AO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_AO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_A_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_BO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_BO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_BQ;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_B_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C5Q;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_CLK;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_CMUX;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_CO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_CO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_CQ;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_C_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_DO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_DO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_DQ;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X12Y121_D_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_AO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_AO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_AQ;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_A_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B5Q;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_BMUX;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_BO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_BO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_BQ;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_B_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_CLK;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_CO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_CO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_CQ;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_C_XOR;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D1;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D2;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D3;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D4;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_DO5;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_DO6;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D_CY;
  wire [0:0] CLBLM_L_X10Y121_SLICE_X13Y121_D_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_AO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_AO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_AQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_A_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_BO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_BO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_BQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_B_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_CLK;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_CO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_CO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_C_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_DO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_DO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X12Y122_D_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_AO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_AO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_AQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_A_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_BMUX;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_BO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_BO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_B_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C5Q;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_CLK;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_CMUX;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_CO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_CO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_CQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_C_XOR;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D1;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D2;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D3;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D4;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_DO5;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_DO6;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_DQ;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D_CY;
  wire [0:0] CLBLM_L_X10Y122_SLICE_X13Y122_D_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_AO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_AQ;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_A_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_BO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_BO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_BQ;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_B_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_CLK;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_CO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_CQ;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_C_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_DMUX;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_DO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X12Y123_D_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_AO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_AO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_A_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_BO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_BO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_BQ;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_B_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CLK;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_CQ;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_C_XOR;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D1;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D2;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D3;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D4;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_DMUX;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_DO5;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D_CY;
  wire [0:0] CLBLM_L_X10Y123_SLICE_X13Y123_D_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_AMUX;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_AO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_AO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_AX;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_A_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_BMUX;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_BO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_BO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_B_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_CE;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_CLK;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_CMUX;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_CO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_CO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_C_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_DO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_DO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_D_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X12Y124_SR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A5Q;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_AMUX;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_AO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_AO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_AQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_AX;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_A_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B5Q;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_BMUX;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_BO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_BO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_BQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_BX;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_B_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C5Q;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_CLK;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_CMUX;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_CO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_CO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_CQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_CX;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_C_XOR;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D1;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D2;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D3;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D4;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D5Q;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_DMUX;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_DO5;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_DO6;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_DQ;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_DX;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D_CY;
  wire [0:0] CLBLM_L_X10Y124_SLICE_X13Y124_D_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_AO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_AO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_A_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_BO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_BO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_BQ;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_B_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_CLK;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_CO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_CO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_CQ;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_C_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_DO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_DO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_DQ;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X12Y125_D_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_AO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_AO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_AQ;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_A_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_BO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_BO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_BQ;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_B_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_CLK;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_CO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_CO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_CQ;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_C_XOR;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D1;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D2;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D3;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D4;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_DMUX;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_DO5;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_DO6;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D_CY;
  wire [0:0] CLBLM_L_X10Y125_SLICE_X13Y125_D_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A5Q;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_AMUX;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_AO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_AO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_AX;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_A_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_BMUX;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_BO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_BO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_B_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_CLK;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_CO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_CO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_CQ;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_C_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_DMUX;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_DO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_DO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X12Y126_D_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_AO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_AO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_AQ;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_A_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_BO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_BO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_BQ;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_B_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_CLK;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_CO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_CO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_CQ;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_C_XOR;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D1;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D2;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D3;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D4;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_DO5;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_DO6;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_DQ;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D_CY;
  wire [0:0] CLBLM_L_X10Y126_SLICE_X13Y126_D_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_AO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_AO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_A_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_BO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_BO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_B_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_CLK;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_CO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_CO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_CQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_C_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_DO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_DO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_DQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X12Y127_D_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_AO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_AO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_AQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_A_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_BO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_BO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_BQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_B_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_CLK;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_CO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_CO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_CQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_C_XOR;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D1;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D2;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D3;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D4;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_DO5;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_DO6;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_DQ;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D_CY;
  wire [0:0] CLBLM_L_X10Y127_SLICE_X13Y127_D_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_AO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_AO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_A_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_BO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_BO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_BQ;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_B_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_CLK;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_CO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_CO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_CQ;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_C_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_DO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_DO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_DQ;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X12Y128_D_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_AO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_AO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_AQ;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_A_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_BO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_BO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_BQ;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_B_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_CLK;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_CMUX;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_CO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_C_XOR;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D1;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D2;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D3;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D4;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_DO5;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_DO6;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D_CY;
  wire [0:0] CLBLM_L_X10Y128_SLICE_X13Y128_D_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A5Q;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_AMUX;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_AO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_AO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_AX;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_A_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_BO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_BO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_BQ;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_B_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_CLK;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_CO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_CO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_C_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_DO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_DO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X12Y129_D_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_AO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_AO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_AQ;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_A_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_BMUX;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_BO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_BO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_B_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_CLK;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_CO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_CO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_C_XOR;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D1;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D2;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D3;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D4;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_DO5;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D_CY;
  wire [0:0] CLBLM_L_X10Y129_SLICE_X13Y129_D_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_AO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_AO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_AX;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_BO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_BO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CE;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CLK;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_DO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_DO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_SR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_AO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_AO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_BO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_BO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_CO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_CO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_DO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_DO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_AO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_AO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_AX;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_BO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_BO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_BX;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_CLK;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_CO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_CO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_DO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_AO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_AO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_BO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_BO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_CO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_CO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_DO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_AMUX;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_AO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_AO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_BMUX;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_BO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_BO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_CO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_CO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_DO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_DO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_AO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_AO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_BO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_BO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_CO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_CO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_DO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_DO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_AO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_AO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_AQ;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_A_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_BO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_BO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_BQ;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_B_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_CLK;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_CO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_CO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_C_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_DO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_DO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X16Y121_D_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_AO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_AO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_A_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_BO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_BO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_B_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_CO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_CO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_C_XOR;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D1;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D2;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D3;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D4;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_DO5;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_DO6;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D_CY;
  wire [0:0] CLBLM_L_X12Y121_SLICE_X17Y121_D_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_AO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_AO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_AQ;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_A_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_BO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_BO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_BQ;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_B_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_CLK;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_CO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_CO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_C_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_DO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_DO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X16Y126_D_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_AO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_AO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_A_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_BO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_BO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_B_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_CO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_CO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_C_XOR;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D1;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D2;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D3;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D4;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_DO5;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_DO6;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D_CY;
  wire [0:0] CLBLM_L_X12Y126_SLICE_X17Y126_D_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_AO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_AO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_AQ;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_A_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_BO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_BO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_B_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_CLK;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_CO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_CO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_C_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_DO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_DO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X16Y127_D_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_AO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_AO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_A_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_BO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_BO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_B_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_CO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_CO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_C_XOR;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D1;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D2;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D3;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D4;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_DO5;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D_CY;
  wire [0:0] CLBLM_L_X12Y127_SLICE_X17Y127_D_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_AMUX;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_AO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_AO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_A_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_BO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_BO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_BQ;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_B_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_CLK;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_CMUX;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_CO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_CO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_C_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_DO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_DO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X10Y116_D_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_AO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_AO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_A_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_BO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_B_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_CO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_C_XOR;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D1;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D2;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D3;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D4;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_DO5;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D_CY;
  wire [0:0] CLBLM_L_X8Y116_SLICE_X11Y116_D_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_AO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_AO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_A_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_BO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_BO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_B_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_CLK;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_CMUX;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_CO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_CO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_C_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_DMUX;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_DO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_DO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X10Y117_D_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_AMUX;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_AO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_AO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_A_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_BO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_BO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_B_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_CO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_C_XOR;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D1;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D2;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D3;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D4;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_DO5;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_DO6;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D_CY;
  wire [0:0] CLBLM_L_X8Y117_SLICE_X11Y117_D_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_AMUX;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_AO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_AO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_A_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_BO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_BO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_BQ;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_B_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_CLK;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_CO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_CO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_CQ;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_C_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_DO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_DO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X10Y118_D_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_AO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_AO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_AQ;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_A_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_BO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_BO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_BQ;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_B_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_CLK;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_CMUX;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_CO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_CO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_C_XOR;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D1;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D2;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D3;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D4;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_DO5;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_DO6;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D_CY;
  wire [0:0] CLBLM_L_X8Y118_SLICE_X11Y118_D_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_AO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_AO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_A_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_BO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_BO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_BQ;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_B_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_CLK;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_CO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_CO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_C_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_DO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_DO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X10Y119_D_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_AO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_AO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_A_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_BO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_BO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_BQ;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_B_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_CLK;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_CO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_CO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_CQ;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_C_XOR;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D1;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D2;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D3;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D4;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_DO5;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_DO6;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D_CY;
  wire [0:0] CLBLM_L_X8Y119_SLICE_X11Y119_D_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_AO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_AO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_A_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_BO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_BO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_BQ;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_B_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_CLK;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_CO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_CO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_C_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_DO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_DO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X10Y120_D_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_AO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_AO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_A_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_BO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_B_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_CO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_CO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_C_XOR;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D1;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D2;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D3;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D4;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_DO5;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_DO6;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D_CY;
  wire [0:0] CLBLM_L_X8Y120_SLICE_X11Y120_D_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_AMUX;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_AO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_AO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_A_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_BO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_BO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_BQ;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_B_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_CLK;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_CO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_CO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_CQ;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_C_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_DMUX;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_DO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X10Y121_D_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_AO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_AO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_A_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_BO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_BO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_B_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_CLK;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_CO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_CO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_CQ;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_C_XOR;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D1;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D2;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D3;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D4;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_DMUX;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_DO5;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_DO6;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D_CY;
  wire [0:0] CLBLM_L_X8Y121_SLICE_X11Y121_D_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A5Q;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_AMUX;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_AO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_AO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_A_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_BO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_BO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_BQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_BX;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_B_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_CLK;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_CO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_CO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_C_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_DO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_DO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X10Y122_D_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A5Q;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_AMUX;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_AO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_AO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_AQ;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_A_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_BO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_BO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_B_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_CLK;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_CO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_CO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_C_XOR;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D1;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D2;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D3;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D4;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_DO5;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_DO6;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D_CY;
  wire [0:0] CLBLM_L_X8Y122_SLICE_X11Y122_D_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_AO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_AO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_A_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_BO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_BO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_BQ;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_B_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C5Q;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_CLK;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_CMUX;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_CO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_CO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_CQ;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_C_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_DO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X10Y123_D_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_AO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_AO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_AQ;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_A_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_BO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_BO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_BQ;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_B_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C5Q;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_CLK;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_CMUX;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_CO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_CO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_CQ;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_C_XOR;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D1;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D2;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D3;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D4;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_DMUX;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_DO5;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_DO6;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D_CY;
  wire [0:0] CLBLM_L_X8Y123_SLICE_X11Y123_D_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_AO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_AO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_AQ;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_A_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B5Q;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_BMUX;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_BO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_BO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_BQ;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_B_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_CLK;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_CO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_CO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_C_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_DO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_DO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X10Y124_D_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_AO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_AO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_A_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_BO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_BO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_BQ;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_B_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_CLK;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_CMUX;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_CO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_CO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_C_XOR;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D1;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D2;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D3;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D4;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_DO5;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_DO6;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D_CY;
  wire [0:0] CLBLM_L_X8Y124_SLICE_X11Y124_D_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_AO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_AO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_A_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_BMUX;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_BO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_BO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_B_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_CLK;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_CO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_CO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_CQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_C_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_DO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_DO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_DQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X10Y125_D_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_AO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_AO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_A_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_BO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_BO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_B_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_CLK;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_CO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_CO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_C_XOR;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D1;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D2;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D3;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D4;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_DO5;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_DO6;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D_CY;
  wire [0:0] CLBLM_L_X8Y125_SLICE_X11Y125_D_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_AMUX;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_AO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_AO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_AX;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_A_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_BO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_BO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_B_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_CE;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_CLK;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_CO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_CO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_C_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_DO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_DO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_D_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X10Y126_SR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_AO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_AO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_AQ;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_A_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B5Q;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_BMUX;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_BO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_BO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_BQ;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_B_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_CLK;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_CO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_CO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_CQ;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_C_XOR;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D1;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D2;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D3;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D4;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_DO5;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_DO6;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_DQ;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D_CY;
  wire [0:0] CLBLM_L_X8Y126_SLICE_X11Y126_D_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_AO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_AO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_AQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_A_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_BO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_BO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_BQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_B_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_CLK;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_CO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_CO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_CQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_C_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_DMUX;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_DO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_DO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X10Y127_D_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_AO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_AO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_A_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_BO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_BO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_BQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_B_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_CLK;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_CO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_CO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_CQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_C_XOR;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D1;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D2;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D3;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D4;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_DO5;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_DO6;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_DQ;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D_CY;
  wire [0:0] CLBLM_L_X8Y127_SLICE_X11Y127_D_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_AO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_AO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_AQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_A_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_BO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_BO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_BQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_B_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_CLK;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_CO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_CO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_CQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_C_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_DO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_DO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X10Y128_D_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_AO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_AO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_AQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_A_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_BO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_BO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_BQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_B_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_CLK;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_CO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_CO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_CQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_C_XOR;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D1;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D2;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D3;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D4;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_DO5;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_DO6;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_DQ;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D_CY;
  wire [0:0] CLBLM_L_X8Y128_SLICE_X11Y128_D_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_AMUX;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_AO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_AO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_AX;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_A_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_BMUX;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_BO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_BO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_B_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_CE;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_CLK;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_CO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_CO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_C_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_DO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_DO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_D_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X10Y129_SR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_AO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_AO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_AQ;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_A_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B5Q;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_BMUX;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_BO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_BO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_BQ;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_B_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_CLK;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_CO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_CO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_C_XOR;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D1;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D2;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D3;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D4;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_DO5;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_DO6;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D_CY;
  wire [0:0] CLBLM_L_X8Y129_SLICE_X11Y129_D_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_AO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_AO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_BO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_BO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_BQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_CLK;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_CO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_CO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_CQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_DO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_DO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_AMUX;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_AO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_AO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_BO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_BO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_CO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_CO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_DO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_DO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AMUX;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AX;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_BMUX;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_BO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_BO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CE;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CLK;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_DO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_DO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_SR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_BO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_BO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CLK;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_DO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D_XOR;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_A;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_A1;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_A2;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_A3;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_A4;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_A5;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_A6;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_AO5;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_AO6;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_A_CY;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_A_XOR;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_B;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_B1;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_B2;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_B3;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_B4;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_B5;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_B6;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_BO5;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_BO6;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_B_CY;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_B_XOR;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_C;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_C1;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_C2;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_C3;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_C4;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_C5;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_C6;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_CO5;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_CO6;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_C_CY;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_C_XOR;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_D;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_D1;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_D2;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_D3;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_D4;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_D5;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_D6;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_DO5;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_DO6;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_D_CY;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X162Y140_D_XOR;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_A;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_A1;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_A2;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_A3;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_A4;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_A5;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_A6;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_AMUX;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_AO5;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_AO6;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_A_CY;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_A_XOR;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_B;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_B1;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_B2;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_B3;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_B4;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_B5;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_B6;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_BO5;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_BO6;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_B_CY;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_B_XOR;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_C;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_C1;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_C2;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_C3;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_C4;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_C5;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_C6;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_CO5;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_CO6;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_C_CY;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_C_XOR;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_D;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_D1;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_D2;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_D3;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_D4;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_D5;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_D6;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_DO5;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_DO6;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_D_CY;
  wire [0:0] CLBLM_R_X103Y140_SLICE_X163Y140_D_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_AO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_AO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_BO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_BO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_CO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_CO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_DO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_DO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_BO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_BO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_CO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_CO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_DO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_DO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D_XOR;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_A;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_A1;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_A2;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_A3;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_A4;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_A5;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_A6;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_AO5;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_AO6;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_A_CY;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_A_XOR;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_B;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_B1;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_B2;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_B3;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_B4;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_B5;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_B6;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_BO5;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_BO6;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_B_CY;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_B_XOR;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_C;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_C1;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_C2;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_C3;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_C4;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_C5;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_C6;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_CO5;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_CO6;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_C_CY;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_C_XOR;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_D;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_D1;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_D2;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_D3;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_D4;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_D5;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_D6;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_DO5;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_DO6;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_D_CY;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X162Y171_D_XOR;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_A;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_A1;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_A2;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_A3;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_A4;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_A5;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_A6;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_AMUX;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_AO5;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_AO6;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_A_CY;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_A_XOR;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_B;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_B1;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_B2;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_B3;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_B4;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_B5;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_B6;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_BMUX;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_BO5;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_BO6;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_B_CY;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_B_XOR;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_C;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_C1;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_C2;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_C3;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_C4;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_C5;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_C6;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_CO5;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_CO6;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_C_CY;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_C_XOR;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_D;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_D1;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_D2;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_D3;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_D4;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_D5;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_D6;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_DO5;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_DO6;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_D_CY;
  wire [0:0] CLBLM_R_X103Y171_SLICE_X163Y171_D_XOR;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A1;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A2;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A3;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A4;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_AO5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_AO6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A_CY;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_A_XOR;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B1;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B2;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B3;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B4;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_BO5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_BO6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B_CY;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_B_XOR;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C1;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C2;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C3;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C4;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_CO5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_CO6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C_CY;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_C_XOR;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D1;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D2;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D3;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D4;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_DO5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_DO6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D_CY;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X162Y173_D_XOR;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A1;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A2;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A3;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A4;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_AMUX;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_AO5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_AO6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A_CY;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_A_XOR;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B1;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B2;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B3;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B4;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_BO5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_BO6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B_CY;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_B_XOR;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C1;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C2;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C3;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C4;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_CO5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_CO6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C_CY;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_C_XOR;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D1;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D2;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D3;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D4;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_DO5;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_DO6;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D_CY;
  wire [0:0] CLBLM_R_X103Y173_SLICE_X163Y173_D_XOR;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_A;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_A1;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_A2;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_A3;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_A4;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_A5;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_A6;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_AO5;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_AO6;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_A_CY;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_A_XOR;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_B;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_B1;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_B2;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_B3;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_B4;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_B5;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_B6;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_BO5;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_BO6;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_B_CY;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_B_XOR;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_C;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_C1;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_C2;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_C3;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_C4;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_C5;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_C6;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_CO5;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_CO6;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_C_CY;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_C_XOR;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_D;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_D1;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_D2;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_D3;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_D4;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_D5;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_D6;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_DO5;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_DO6;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_D_CY;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X162Y175_D_XOR;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_A;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_A1;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_A2;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_A3;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_A4;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_A5;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_A6;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_AO5;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_AO6;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_A_CY;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_A_XOR;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_B;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_B1;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_B2;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_B3;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_B4;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_B5;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_B6;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_BO5;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_BO6;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_B_CY;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_B_XOR;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_C;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_C1;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_C2;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_C3;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_C4;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_C5;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_C6;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_CO5;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_CO6;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_C_CY;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_C_XOR;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_D;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_D1;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_D2;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_D3;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_D4;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_D5;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_D6;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_DO5;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_DO6;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_D_CY;
  wire [0:0] CLBLM_R_X103Y175_SLICE_X163Y175_D_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_AO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_AO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_BO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_BO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_CO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_CO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_DO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_DO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AMUX;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_BO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_BO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_CO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_CO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_DO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_DO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_AO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_A_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_BO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_BO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_BQ;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_B_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_CLK;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_CO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_CO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_C_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_DO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X14Y119_D_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_AMUX;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_AO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_AO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_A_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_BO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_BO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_B_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_CO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_C_XOR;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D1;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D2;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D3;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D4;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_DO5;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_DO6;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D_CY;
  wire [0:0] CLBLM_R_X11Y119_SLICE_X15Y119_D_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_AO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_AO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_A_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_BO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_BO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_BQ;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_B_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_CLK;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_CO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_CO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_CQ;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_C_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_DO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X14Y120_D_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_AO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_AO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_AQ;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_A_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_BMUX;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_BO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_BO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_B_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_CLK;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_CMUX;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_CO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_CO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_C_XOR;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D1;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D2;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D3;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D4;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_DO5;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_DO6;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D_CY;
  wire [0:0] CLBLM_R_X11Y120_SLICE_X15Y120_D_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_AO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_AO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_AQ;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_A_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_BO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_BO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_BQ;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_B_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_CLK;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_CO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_CQ;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_C_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_DO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X14Y121_D_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_AO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_AO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_AQ;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_A_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_BO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_BO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_B_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_CLK;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_CO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_CO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_C_XOR;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D1;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D2;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D3;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D4;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_DO5;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D_CY;
  wire [0:0] CLBLM_R_X11Y121_SLICE_X15Y121_D_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_AO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_AO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_A_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_BO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_BO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_BQ;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_B_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_CLK;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_CO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_CO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_CQ;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_C_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_DO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_DO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_DQ;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X14Y122_D_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_AO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_AO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_AQ;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_A_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_BO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_BO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_BQ;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_B_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_CLK;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_CO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_CO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_C_XOR;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D1;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D2;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D3;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D4;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_DO5;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_DO6;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D_CY;
  wire [0:0] CLBLM_R_X11Y122_SLICE_X15Y122_D_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_AO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_AO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_AQ;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_A_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_BO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_BO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_BQ;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_B_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_CLK;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_CO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_CO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_CQ;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_C_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_DO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_DO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_DQ;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X14Y123_D_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_AO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_AO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_AQ;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_A_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_BO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_BO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_B_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_CLK;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_CO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_CO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_C_XOR;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D1;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D2;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D3;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D4;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_DO5;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_DO6;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D_CY;
  wire [0:0] CLBLM_R_X11Y123_SLICE_X15Y123_D_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A5Q;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_AMUX;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_AO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_AO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_AQ;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_A_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_BO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_BO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_BQ;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_B_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_CLK;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_CO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_CO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_CQ;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_C_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_DMUX;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_DO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_DO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X14Y124_D_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_AO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_AO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_A_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_BO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_BO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_B_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_CO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_CO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_C_XOR;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D1;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D2;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D3;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D4;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_DO5;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D_CY;
  wire [0:0] CLBLM_R_X11Y124_SLICE_X15Y124_D_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_AO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_AO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_A_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_BO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_BO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_BQ;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_B_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_CLK;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_CO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_CO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_CQ;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_C_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_DO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_DO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X14Y125_D_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_AO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_AO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_A_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_BO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_BO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_B_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_CO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_CO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_C_XOR;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D1;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D2;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D3;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D4;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_DO5;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_DO6;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D_CY;
  wire [0:0] CLBLM_R_X11Y125_SLICE_X15Y125_D_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_AMUX;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_AO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_AO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_AQ;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_A_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_BO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_BO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_BQ;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_B_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_CLK;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_CO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_CO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_CQ;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_C_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_DO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_DO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_DQ;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X14Y126_D_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_AO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_AO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_AQ;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_A_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_BO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_BO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_BQ;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_B_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_CLK;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_CO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_CO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_CQ;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_C_XOR;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D1;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D2;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D3;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D4;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_DMUX;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_DO5;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_DO6;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D_CY;
  wire [0:0] CLBLM_R_X11Y126_SLICE_X15Y126_D_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_AO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_AO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_AQ;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_A_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_BMUX;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_BO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_BO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_B_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_CLK;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_CO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_CO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_C_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_DO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_DO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X14Y127_D_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_AO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_AO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_AQ;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_A_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_BMUX;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_BO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_BO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_B_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_CLK;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_CMUX;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_CO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_CO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_C_XOR;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D1;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D2;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D3;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D4;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_DMUX;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_DO5;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_DO6;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D_CY;
  wire [0:0] CLBLM_R_X11Y127_SLICE_X15Y127_D_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_AMUX;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_AO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_AO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_AX;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_A_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_BO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_BO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_B_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_CE;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_CLK;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_CO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_CO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_C_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_DO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_DO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_D_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X14Y128_SR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_AO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_AO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_A_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_BO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_BO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_B_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_CLK;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_CO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_CO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_C_XOR;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D1;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D2;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D3;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D4;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_DO5;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_DO6;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D_CY;
  wire [0:0] CLBLM_R_X11Y128_SLICE_X15Y128_D_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_AO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_AO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_A_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_BO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_BO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_BQ;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_B_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_CLK;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_CO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_CO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_C_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_DMUX;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_DO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_DO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X14Y129_D_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_AMUX;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_AO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_AO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_A_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_BO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_BO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_B_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_CO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_CO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_C_XOR;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D1;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D2;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D3;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D4;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_DO5;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_DO6;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D_CY;
  wire [0:0] CLBLM_R_X11Y129_SLICE_X15Y129_D_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_AO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_AO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_AQ;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_A_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_BMUX;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_BO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_BO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_B_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_CLK;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_CO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_CO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_C_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_DO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_DO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X14Y130_D_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_AO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_AO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_A_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_BO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_BO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_B_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_CO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_CO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_C_XOR;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D1;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D2;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D3;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D4;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_DO5;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_DO6;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D_CY;
  wire [0:0] CLBLM_R_X11Y130_SLICE_X15Y130_D_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_AO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_AO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_BO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_BO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_CO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_DO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_DO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_AO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_AO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_AQ;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_BO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_BO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_CLK;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_CO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_CO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_DO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_DO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_AO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_AO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_BO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_BO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_CO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_CO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_DO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_DO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_AO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_AO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_BO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_BO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_CO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_CO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_DO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_DO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_AO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_AO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_A_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_BO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_BO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_B_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_CLK;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_CO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_C_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_DO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X18Y127_D_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_AO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_AO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_A_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_BO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_BO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_B_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_CO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_C_XOR;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D1;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D2;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D3;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D4;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_DO5;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_DO6;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D_CY;
  wire [0:0] CLBLM_R_X13Y127_SLICE_X19Y127_D_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_AO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_A_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_BMUX;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_BO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_B_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_CLK;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_CMUX;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_CO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_C_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_DO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X2Y118_D_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_AO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_AQ;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_A_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_BO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_BQ;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_B_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_CLK;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_CMUX;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_CO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_C_XOR;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D1;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D2;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D3;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D4;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_DO5;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D_CY;
  wire [0:0] CLBLM_R_X3Y118_SLICE_X3Y118_D_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_AO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_AQ;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_A_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_BO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_BQ;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_B_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_CLK;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_CMUX;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_CO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_C_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_DO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_DO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X2Y119_D_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_AO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_AQ;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_A_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_BMUX;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_BO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_B_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_CLK;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_CO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_C_XOR;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D1;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D2;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D3;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D4;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_DO5;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D_CY;
  wire [0:0] CLBLM_R_X3Y119_SLICE_X3Y119_D_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_AQ;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_A_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_BO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_BQ;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_B_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_CLK;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_CO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_CQ;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_C_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_DO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X2Y120_D_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_AO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_AO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_AQ;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_A_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_BO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_BQ;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_B_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_CLK;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_CO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_C_XOR;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D1;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D2;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D3;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D4;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_DO5;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D_CY;
  wire [0:0] CLBLM_R_X3Y120_SLICE_X3Y120_D_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_AO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_AQ;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_A_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_BO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_BQ;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_B_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C5Q;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_CLK;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_CMUX;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_CO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_CQ;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_C_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_DO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_DO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X2Y121_D_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_AO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_AO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_AQ;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_A_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_BO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_BQ;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_B_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_CLK;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_CMUX;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_CO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_C_XOR;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D1;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D2;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D3;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D4;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_DO5;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_DO6;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D_CY;
  wire [0:0] CLBLM_R_X3Y121_SLICE_X3Y121_D_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A5Q;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_AMUX;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_AO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_AQ;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_AX;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_A_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_BMUX;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_BO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_BO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_B_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_CLK;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_CO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_CQ;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_C_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_DO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_DO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_DQ;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X2Y122_D_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_AO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_AQ;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_A_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_BO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_BQ;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_B_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_CLK;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_CMUX;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_CO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_CO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_C_XOR;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D1;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D2;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D3;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D4;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_DO5;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_DO6;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D_CY;
  wire [0:0] CLBLM_R_X3Y122_SLICE_X3Y122_D_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_AO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_AO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_AQ;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_A_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_BO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_BO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_BQ;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_B_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_CLK;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_CO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_CO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_CQ;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_C_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_DO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_DO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_DQ;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X2Y123_D_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_AO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_AO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_AQ;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_A_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_BO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_BO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_BQ;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_B_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_CLK;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_CO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_CQ;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_C_XOR;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D1;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D2;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D3;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D4;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_DO5;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_DO6;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D_CY;
  wire [0:0] CLBLM_R_X3Y123_SLICE_X3Y123_D_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A5Q;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_AMUX;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_AO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_AQ;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_A_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B5Q;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_BMUX;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_BO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_BO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_BQ;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_B_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_CLK;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_CO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_CO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_CQ;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_C_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_DO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_DO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_DQ;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X2Y124_D_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_AO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_AO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_AQ;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_A_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_BO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_BO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_BQ;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_B_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C5Q;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_CLK;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_CMUX;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_CO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_CO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_CQ;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_C_XOR;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D1;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D2;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D3;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D4;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_DO5;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_DO6;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D_CY;
  wire [0:0] CLBLM_R_X3Y124_SLICE_X3Y124_D_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_AO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_AO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_AQ;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_A_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_BO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_B_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_CLK;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_CO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_CO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_C_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_DO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_DO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X2Y125_D_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_AO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_AQ;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_A_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_BO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_BO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_BQ;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_B_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_CLK;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_CMUX;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_CO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_CO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_C_XOR;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D1;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D2;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D3;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D4;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_DO5;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_DO6;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D_CY;
  wire [0:0] CLBLM_R_X3Y125_SLICE_X3Y125_D_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A5Q;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_AMUX;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_AO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_AO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_AQ;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_AX;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_A_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_BO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_BO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_B_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_CLK;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_CO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_CO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_C_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_DMUX;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_DO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_DO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X2Y126_D_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_AO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_AO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_A_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_BMUX;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_BO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_B_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_CO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_CO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_C_XOR;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D1;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D2;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D3;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D4;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_DO5;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_DO6;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D_CY;
  wire [0:0] CLBLM_R_X3Y126_SLICE_X3Y126_D_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_AO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_A_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_BO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_BO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_B_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_CMUX;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_CO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_CO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_C_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_DMUX;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_DO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_DO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X2Y127_D_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_AMUX;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_AO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_AO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_A_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_BO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_BO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_B_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_CMUX;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_CO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_CO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_C_XOR;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D1;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D2;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D3;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D4;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_DO5;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_DO6;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D_CY;
  wire [0:0] CLBLM_R_X3Y127_SLICE_X3Y127_D_XOR;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A1;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A2;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A3;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A4;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_AO5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_AO6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A_CY;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_A_XOR;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B1;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B2;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B3;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B4;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_BO5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_BO6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B_CY;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_B_XOR;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C1;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C2;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C3;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C4;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_CO5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_CO6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C_CY;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_C_XOR;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D1;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D2;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D3;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D4;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_DO5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_DO6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D_CY;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X2Y128_D_XOR;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A1;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A2;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A3;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A4;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_AMUX;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_AO5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_AO6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A_CY;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_A_XOR;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B1;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B2;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B3;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B4;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_BO5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_BO6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B_CY;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_B_XOR;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C1;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C2;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C3;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C4;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_CO5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_CO6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C_CY;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_C_XOR;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D1;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D2;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D3;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D4;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_DO5;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_DO6;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D_CY;
  wire [0:0] CLBLM_R_X3Y128_SLICE_X3Y128_D_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_AO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_AO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_AQ;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_A_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_BO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_BO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_B_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_CLK;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_CO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_CO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_C_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_DO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_DO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X2Y129_D_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_AMUX;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_AO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_AO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_A_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_BO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_BO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_B_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_CMUX;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_CO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_CO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_C_XOR;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D1;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D2;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D3;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D4;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_DMUX;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_DO5;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D_CY;
  wire [0:0] CLBLM_R_X3Y129_SLICE_X3Y129_D_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_AMUX;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_AO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_AO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_BMUX;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_BO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_BO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_CO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_CO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_DMUX;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_DO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_DO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_AMUX;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_AO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_AO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_BO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_BO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_CO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_CO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_DO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_DO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_AO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_AO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_AQ;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_BO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_BO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_BQ;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_CLK;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_CMUX;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_CO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_CO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_DO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_DO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_AO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_AO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_BO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_BO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_CO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_CO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_DO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_DO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A5Q;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_AMUX;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_AO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_AO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_AX;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_BO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_BO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_BQ;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_CLK;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_CMUX;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_CO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_CO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_DO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_DO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_AO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_AO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_BO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_BO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_CO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_CO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_DO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_DO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_AQ;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_A_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_BO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_B_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CLK;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_C_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_DO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X6Y116_D_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_A_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_BO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_BO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_BQ;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_B_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CLK;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_CQ;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_C_XOR;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D1;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D2;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D3;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D4;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_DMUX;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_DO5;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D_CY;
  wire [0:0] CLBLM_R_X5Y116_SLICE_X7Y116_D_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A5Q;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_AMUX;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_AO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_AO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_AQ;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_AX;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_A_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_BO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_BO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_BQ;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_B_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_CLK;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_CO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_CO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_CQ;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_C_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_DMUX;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_DO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_DO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X6Y117_D_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_AO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_AO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_A_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_BMUX;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_BO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_BO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_B_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_CLK;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_CO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_CO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_C_XOR;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D1;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D2;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D3;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D4;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_DO5;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_DO6;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D_CY;
  wire [0:0] CLBLM_R_X5Y117_SLICE_X7Y117_D_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_AMUX;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_AO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_AO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_A_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B5Q;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_BMUX;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_BO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_BX;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_B_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_CLK;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_CMUX;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_CO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_CO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_C_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_DO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_DQ;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X6Y118_D_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A5Q;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_AMUX;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_AO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_AO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_AQ;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_AX;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_A_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_BMUX;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_BO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_BO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_B_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_CLK;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_CO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_C_XOR;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D1;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D2;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D3;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D4;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_DO5;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D_CY;
  wire [0:0] CLBLM_R_X5Y118_SLICE_X7Y118_D_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_AO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_AO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_AQ;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_A_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_BMUX;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_BO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_BO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_B_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CLK;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_CQ;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_C_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_DO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_DO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_DQ;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X6Y119_D_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_AO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_AO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_A_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_BO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_BQ;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_B_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_CLK;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_CO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_CO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_CQ;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_C_XOR;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D1;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D2;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D3;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D4;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_DO5;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_DO6;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D_CY;
  wire [0:0] CLBLM_R_X5Y119_SLICE_X7Y119_D_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_AO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_AO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_A_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_BO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_BO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_BQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_B_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CLK;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_CQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_C_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_DO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_DQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X6Y120_D_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A5Q;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_AMUX;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_AO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_AO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_A_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_BO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_BO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_BQ;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_B_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_CLK;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_CO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_CO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_C_XOR;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D1;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D2;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D3;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D4;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_DO5;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_DO6;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D_CY;
  wire [0:0] CLBLM_R_X5Y120_SLICE_X7Y120_D_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_AO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_AO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_A_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_BO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_BO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_B_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_CLK;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_CMUX;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_CO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_CO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_C_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_DO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_DO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X6Y121_D_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_AO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_AO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_AQ;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_A_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_BMUX;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_BO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_BO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_B_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_CLK;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_CO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_CO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_C_XOR;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D1;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D2;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D3;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D4;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_DO5;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_DO6;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D_CY;
  wire [0:0] CLBLM_R_X5Y121_SLICE_X7Y121_D_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_AO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_AO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_AQ;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_A_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_BO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_BO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_B_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_CLK;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_CO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_CO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_CQ;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_C_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_DMUX;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_DO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X6Y122_D_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_AO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_AO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_AQ;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_A_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_BO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_BO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_BQ;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_B_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_CLK;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_CO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_CO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_C_XOR;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D1;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D2;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D3;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D4;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_DO5;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_DO6;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D_CY;
  wire [0:0] CLBLM_R_X5Y122_SLICE_X7Y122_D_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_AO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_AO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_AQ;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_A_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B5Q;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_BMUX;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_BO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_BO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_BQ;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_B_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_CLK;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_CO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_CO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_CQ;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_C_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_DO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_DO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X6Y123_D_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_AO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_AO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_AQ;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_A_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_BO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_BO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_BQ;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_B_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C5Q;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_CLK;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_CMUX;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_CO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_CO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_CQ;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_C_XOR;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D1;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D2;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D3;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D4;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_DO5;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_DO6;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D_CY;
  wire [0:0] CLBLM_R_X5Y123_SLICE_X7Y123_D_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A5Q;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_AMUX;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_AO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_AO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_AX;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_A_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_BO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_BO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_B_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_CLK;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_CO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_CO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_CQ;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_C_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_DMUX;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_DO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_DO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X6Y124_D_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_AO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_AO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_A_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_BO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_BO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_BQ;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_B_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C5Q;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_CLK;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_CMUX;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_CO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_CO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_CQ;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_C_XOR;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D1;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D2;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D3;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D4;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_DO5;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_DO6;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D_CY;
  wire [0:0] CLBLM_R_X5Y124_SLICE_X7Y124_D_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A5Q;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_AMUX;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_AO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_AO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_AX;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_A_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_BO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_BO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_BQ;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_B_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_CLK;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_CMUX;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_CO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_CO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_C_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_DO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X6Y125_D_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_AO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_AO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_AQ;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_A_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_BO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_BO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_BQ;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_B_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_CLK;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_CO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_CO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_C_XOR;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D1;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D2;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D3;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D4;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_DO5;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_DO6;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D_CY;
  wire [0:0] CLBLM_R_X5Y125_SLICE_X7Y125_D_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_BO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_BO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_BQ;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_CLK;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_CO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_CO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_CQ;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_DO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_DO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_DQ;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A5Q;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_AMUX;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_AO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_AO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_AQ;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_BO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_BO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_BQ;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_CLK;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_CMUX;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_CO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_DO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_DO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_AO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_AO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_BO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_BO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CLK;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_DO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_DO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_AO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_AO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B5Q;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_BMUX;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_BO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_BO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_BQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_CLK;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_CO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_CO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_CQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_DO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_DO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A5Q;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_AMUX;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_AO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_AO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_AX;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_BO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_BO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_CLK;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_CMUX;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_CO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_CO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_DO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_DO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_DQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A5Q;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_AMUX;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_AO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_AO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_AQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B5Q;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_BMUX;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_BO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_BO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_BQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_CLK;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_CO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_CO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_DO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_DO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_AO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_AO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_AQ;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_BO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_BO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_BQ;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_CLK;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_CO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_CO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_CQ;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_DO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_DO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_AO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_AO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_BO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_BO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_CLK;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_CO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_CO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_DO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_DO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_AO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_AO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_BO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_BO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_CLK;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_CO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_CO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_DO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_DO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_AO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_AO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_AQ;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_BO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_BO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_BQ;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_CLK;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_CMUX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_CO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_CO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_DO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_DO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_AMUX;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_AO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_A_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_BO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_BO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_B_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_CO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_CO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_C_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_DO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_DO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X8Y115_D_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_AMUX;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_AO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_AO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_A_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_BO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_BO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_B_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_CO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_CO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_C_XOR;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D1;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D2;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D3;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D4;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_DO5;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D_CY;
  wire [0:0] CLBLM_R_X7Y115_SLICE_X9Y115_D_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_AO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_AO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_AQ;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_A_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_BMUX;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_BO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_B_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_CLK;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_CO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_C_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_DO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X8Y116_D_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_AO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_AO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_AQ;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_A_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_BO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_BO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_BQ;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_B_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_CLK;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_CO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_C_XOR;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D1;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D2;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D3;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D4;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_DO5;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_DO6;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D_CY;
  wire [0:0] CLBLM_R_X7Y116_SLICE_X9Y116_D_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_AO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_AO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_A_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_BO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_BO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_B_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_CLK;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_CO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_CO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_CQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_C_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_DO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_DO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_DQ;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X8Y117_D_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_AMUX;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_AO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_AO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_A_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_BMUX;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_BO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_BO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_B_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_CO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_CO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_C_XOR;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D1;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D2;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D3;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D4;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_DO5;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_DO6;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D_CY;
  wire [0:0] CLBLM_R_X7Y117_SLICE_X9Y117_D_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_AO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_AO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_AQ;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_A_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_BO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_BO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_B_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C5Q;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_CLK;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_CMUX;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_CO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_CO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_C_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_DO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_DO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_DQ;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X8Y118_D_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_AO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_AO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_AQ;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_A_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_BMUX;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_BO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_BO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_B_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_CLK;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_CO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_CO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_C_XOR;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D1;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D2;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D3;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D4;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_DO5;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_DO6;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D_CY;
  wire [0:0] CLBLM_R_X7Y118_SLICE_X9Y118_D_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_A_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_BO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_BQ;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_B_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CLK;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_CQ;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_C_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_DO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_DO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_DQ;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X8Y119_D_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_AO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_AO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_AQ;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_A_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_BO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_BO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_BQ;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_B_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_CLK;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_CO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_CO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_C_XOR;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D1;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D2;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D3;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D4;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_DO5;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_DO6;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D_CY;
  wire [0:0] CLBLM_R_X7Y119_SLICE_X9Y119_D_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_AO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_AO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_AQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_A_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_BO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_BO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_BQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_B_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CLK;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_CQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_C_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_DO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_DQ;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X8Y120_D_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_AO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_A_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_BO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_BO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_B_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_CO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_C_XOR;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D1;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D2;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D3;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D4;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_DO5;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_DO6;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D_CY;
  wire [0:0] CLBLM_R_X7Y120_SLICE_X9Y120_D_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A5Q;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AMUX;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_AX;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_A_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_BO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_BO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_B_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CLK;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_C_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_DMUX;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_DO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X8Y121_D_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_A_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B5Q;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_BMUX;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_BO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_BO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_B_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CLK;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_C_XOR;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D1;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D2;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D3;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D4;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_DO5;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D_CY;
  wire [0:0] CLBLM_R_X7Y121_SLICE_X9Y121_D_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_AO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_AO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_A_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_BO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_BO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_B_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_CLK;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_CO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_CO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_C_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_DMUX;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_DO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X8Y122_D_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_AO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_AO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_AQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_A_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_BO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_BO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_B_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_CLK;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_CO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_CO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_CQ;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_C_XOR;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D1;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D2;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D3;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D4;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_DO5;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_DO6;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D_CY;
  wire [0:0] CLBLM_R_X7Y122_SLICE_X9Y122_D_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_AO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_AO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_A_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B5Q;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_BMUX;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_BO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_BO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_B_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_CLK;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_CMUX;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_CO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_CO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_C_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_DO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_DO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X8Y123_D_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A5Q;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_AMUX;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_AO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_AO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_AQ;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_A_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_BO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_BO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_BQ;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_B_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_CLK;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_CO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_CO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_CQ;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_C_XOR;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D1;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D2;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D3;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D4;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_DMUX;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_DO5;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_DO6;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D_CY;
  wire [0:0] CLBLM_R_X7Y123_SLICE_X9Y123_D_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_AO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_AO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_A_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B5Q;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_BMUX;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_BO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_BO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_B_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_CLK;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_CMUX;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_CO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_CO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_C_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_DO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X8Y124_D_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_AO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_AO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_AQ;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_A_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_BMUX;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_BO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_BO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_B_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_CLK;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_CO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_CO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_C_XOR;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D1;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D2;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D3;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D4;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_DO5;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_DO6;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D_CY;
  wire [0:0] CLBLM_R_X7Y124_SLICE_X9Y124_D_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_AO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_AO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_AQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_A_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_BO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_BO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_BQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_B_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_CLK;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_CO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_CO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_C_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_DO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_DO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_DQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X8Y125_D_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A5Q;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_AMUX;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_AO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_AQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_AX;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_A_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B5Q;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_BMUX;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_BO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_BX;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_B_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_CLK;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_CO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_CQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_C_XOR;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D1;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D2;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D3;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D4;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_DO5;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_DO6;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_DQ;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D_CY;
  wire [0:0] CLBLM_R_X7Y125_SLICE_X9Y125_D_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_AO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_AO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_AQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_A_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_BO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_BO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_B_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_CLK;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_CO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_CO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_CQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_C_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_DO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_DO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X8Y126_D_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_AO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_AO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_A_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B5Q;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_BMUX;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_BO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_BO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_BQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_B_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C5Q;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_CLK;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_CMUX;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_CO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_CO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_CQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_C_XOR;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D1;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D2;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D3;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D4;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D5Q;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_DMUX;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_DO5;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_DO6;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_DQ;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D_CY;
  wire [0:0] CLBLM_R_X7Y126_SLICE_X9Y126_D_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_AO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_AO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_A_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_BO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_BO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_BQ;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_B_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_CLK;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_CO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_CO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_CQ;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_C_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_DO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_DO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_DQ;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X8Y127_D_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_AO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_AO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_AQ;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_A_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_BO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_BO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_BQ;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_B_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_CLK;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_CO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_CO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_CQ;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_C_XOR;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D1;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D2;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D3;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D4;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_DMUX;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_DO5;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_DO6;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D_CY;
  wire [0:0] CLBLM_R_X7Y127_SLICE_X9Y127_D_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_AO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_AO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_A_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_BO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_BO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_BQ;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_B_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_CLK;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_CO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_CO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_CQ;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_C_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_DO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_DO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_DQ;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X8Y128_D_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_AO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_AO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_AQ;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_A_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_BMUX;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_BO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_BO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_B_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_CLK;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_CO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_CO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_C_XOR;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D1;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D2;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D3;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D4;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_DO5;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_DO6;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D_CY;
  wire [0:0] CLBLM_R_X7Y128_SLICE_X9Y128_D_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A5Q;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_AMUX;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_AO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_AO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_BO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_BO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_BQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_CLK;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_CO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_CO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_CQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_DO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_DO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_DQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_AO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_AO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_AQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_BO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_BO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_BQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_CLK;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_CO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_CO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_CQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_DO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_DO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_DQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_AO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_AO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_BO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_BO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_CLK;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_CMUX;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_CO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_DO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_DO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_AO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_AO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_AQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_BMUX;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_BO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_BO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_CLK;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_CMUX;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_CO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_CO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_DMUX;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_DO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_DO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_AO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_AO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_BMUX;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_BO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_BO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CLK;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CMUX;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_DO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_DO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_AO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_AO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_BMUX;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_BO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_BO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_CLK;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_CO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_CO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_DO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_DO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D_XOR;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_O;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_O;
  wire [0:0] LIOB33_SING_X0Y150_IOB_X0Y150_O;
  wire [0:0] LIOB33_SING_X0Y199_IOB_X0Y199_O;
  wire [0:0] LIOB33_SING_X0Y50_IOB_X0Y50_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_O;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y151_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y152_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y153_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y154_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y155_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y156_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y157_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y158_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y159_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y160_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y161_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y162_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y163_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y164_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y165_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y166_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y167_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y168_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y169_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y170_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y171_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y172_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y173_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y174_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y175_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y176_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y177_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y178_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y179_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y180_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y181_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y182_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y183_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y184_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y185_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y186_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y187_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y188_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y189_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y190_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y191_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y192_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y193_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y194_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y195_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y196_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y197_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y198_O;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y51_I;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y52_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y53_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y54_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y55_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y56_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y57_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y58_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y59_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y60_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y61_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y62_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y63_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y64_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y65_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y66_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y67_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y68_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y69_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y70_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y71_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y72_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y73_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y74_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y75_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y76_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y77_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y78_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y79_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y80_O;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_D;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_O;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_TQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_TQ;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_O;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_O;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y73_D;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y73_O;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_D;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_O;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_D;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_O;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_D1;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_OQ;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_T1;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_TQ;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_I;
  wire [0:0] RIOB33_SING_X105Y149_IOB_X1Y149_I;
  wire [0:0] RIOB33_SING_X105Y150_IOB_X1Y150_O;
  wire [0:0] RIOB33_SING_X105Y199_IOB_X1Y199_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y114_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y115_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y116_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y117_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y118_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y119_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y120_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y121_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y122_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y123_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y124_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y125_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y126_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y127_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y128_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y129_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y130_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y131_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y132_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y133_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y134_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y135_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y136_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y137_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y138_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y139_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y140_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y141_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y142_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y143_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y144_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y145_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y146_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y147_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y148_I;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y151_O;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y152_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y153_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y154_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y155_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y156_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y157_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y158_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y159_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y160_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y161_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y162_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y163_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y164_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y165_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y166_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y167_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y168_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y169_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y170_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y171_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y172_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y173_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y174_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y175_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y176_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y177_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y178_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y179_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y180_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y181_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y182_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y183_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y184_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y185_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y186_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y187_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y188_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y189_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y190_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y191_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y192_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y193_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y194_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y195_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y196_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y197_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y198_O;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_D;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_O;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_D;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_O;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_O;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_TQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_TQ;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_DO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_CO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_BO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a0a0a0f0f0f0f)
  ) CLBLL_L_X2Y115_SLICE_X0Y115_ALUT (
.I0(CLBLM_R_X3Y120_SLICE_X3Y120_CO6),
.I1(1'b1),
.I2(CLBLL_L_X2Y119_SLICE_X0Y119_AO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X0Y115_AO5),
.O6(CLBLL_L_X2Y115_SLICE_X0Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_DO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_CO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_BO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y115_SLICE_X1Y115_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y115_SLICE_X1Y115_AO5),
.O6(CLBLL_L_X2Y115_SLICE_X1Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_DO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeefffffffaff)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_CLUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(CLBLM_R_X3Y128_SLICE_X3Y128_BO6),
.I2(CLBLL_L_X2Y127_SLICE_X0Y127_CO6),
.I3(RIOB33_X105Y137_IOB_X1Y137_I),
.I4(RIOB33_X105Y127_IOB_X1Y128_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_CO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefefffffffaffff)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_BLUT (
.I0(RIOB33_X105Y127_IOB_X1Y128_I),
.I1(CLBLL_L_X4Y128_SLICE_X4Y128_AO6),
.I2(RIOB33_X105Y129_IOB_X1Y129_I),
.I3(CLBLL_L_X2Y119_SLICE_X0Y119_CO6),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_BO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeefffffefeffff)
  ) CLBLL_L_X2Y117_SLICE_X0Y117_ALUT (
.I0(RIOB33_X105Y127_IOB_X1Y128_I),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(CLBLM_R_X3Y126_SLICE_X3Y126_AO6),
.I3(CLBLM_R_X3Y127_SLICE_X2Y127_DO6),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X0Y117_AO5),
.O6(CLBLL_L_X2Y117_SLICE_X0Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_DO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_CO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_BO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y117_SLICE_X1Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y117_SLICE_X1Y117_AO5),
.O6(CLBLL_L_X2Y117_SLICE_X1Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_DO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_CO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_BO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeefffffffaffff)
  ) CLBLL_L_X2Y118_SLICE_X0Y118_ALUT (
.I0(RIOB33_X105Y127_IOB_X1Y128_I),
.I1(CLBLM_R_X3Y130_SLICE_X3Y130_BO6),
.I2(CLBLM_R_X3Y128_SLICE_X2Y128_AO6),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X0Y118_AO5),
.O6(CLBLL_L_X2Y118_SLICE_X0Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y118_SLICE_X1Y118_AO5),
.Q(CLBLL_L_X2Y118_SLICE_X1Y118_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y118_SLICE_X2Y118_BO5),
.Q(CLBLL_L_X2Y118_SLICE_X1Y118_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y118_SLICE_X1Y118_AO6),
.Q(CLBLL_L_X2Y118_SLICE_X1Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y118_SLICE_X1Y118_BO6),
.Q(CLBLL_L_X2Y118_SLICE_X1Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_DO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff55553cc336c9)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_CLUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(CLBLL_L_X2Y119_SLICE_X0Y119_CO6),
.I2(CLBLL_L_X2Y118_SLICE_X1Y118_BQ),
.I3(CLBLM_R_X3Y120_SLICE_X3Y120_CO6),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_CO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heefe4454bbab1101)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X2Y118_SLICE_X1Y118_BQ),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.I5(CLBLL_L_X2Y119_SLICE_X0Y119_CO6),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_BO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00ccaaccaa)
  ) CLBLL_L_X2Y118_SLICE_X1Y118_ALUT (
.I0(CLBLL_L_X2Y118_SLICE_X1Y118_B5Q),
.I1(CLBLL_L_X2Y118_SLICE_X1Y118_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y118_SLICE_X1Y118_AO5),
.O6(CLBLL_L_X2Y118_SLICE_X1Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9966669999666699)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_DLUT (
.I0(CLBLM_R_X3Y130_SLICE_X3Y130_BO6),
.I1(CLBLM_R_X3Y127_SLICE_X2Y127_DO6),
.I2(1'b1),
.I3(CLBLL_L_X2Y127_SLICE_X0Y127_CO6),
.I4(CLBLM_R_X3Y128_SLICE_X2Y128_AO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_DO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9696696969699696)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_CLUT (
.I0(CLBLM_R_X3Y128_SLICE_X3Y128_BO6),
.I1(CLBLM_R_X3Y126_SLICE_X3Y126_AO6),
.I2(CLBLL_L_X4Y128_SLICE_X4Y128_AO6),
.I3(1'b1),
.I4(CLBLL_L_X4Y126_SLICE_X4Y126_DO6),
.I5(CLBLL_L_X2Y119_SLICE_X0Y119_DO6),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_CO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdcff50dcdc5050)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_BLUT (
.I0(CLBLL_L_X2Y121_SLICE_X0Y121_BO5),
.I1(CLBLM_R_X3Y119_SLICE_X2Y119_CO5),
.I2(CLBLL_L_X4Y126_SLICE_X4Y126_DO6),
.I3(CLBLM_R_X3Y128_SLICE_X2Y128_AO6),
.I4(CLBLM_R_X3Y128_SLICE_X3Y128_BO6),
.I5(LIOB33_X0Y51_IOB_X0Y51_I),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_BO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffec0000ffa00000)
  ) CLBLL_L_X2Y119_SLICE_X0Y119_ALUT (
.I0(LIOB33_X0Y53_IOB_X0Y53_I),
.I1(CLBLM_R_X3Y126_SLICE_X3Y126_AO6),
.I2(CLBLL_L_X4Y128_SLICE_X4Y128_AO6),
.I3(CLBLL_L_X2Y119_SLICE_X0Y119_BO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X5Y120_SLICE_X7Y120_A5Q),
.O5(CLBLL_L_X2Y119_SLICE_X0Y119_AO5),
.O6(CLBLL_L_X2Y119_SLICE_X0Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y119_SLICE_X1Y119_AO6),
.Q(CLBLL_L_X2Y119_SLICE_X1Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_DO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_CO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000202020202)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_BLUT (
.I0(CLBLM_R_X3Y119_SLICE_X3Y119_BO5),
.I1(CLBLM_R_X7Y117_SLICE_X9Y117_DO6),
.I2(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I3(CLBLM_R_X5Y120_SLICE_X7Y120_A5Q),
.I4(CLBLM_R_X3Y119_SLICE_X2Y119_CO5),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_BO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf088f088f044f044)
  ) CLBLL_L_X2Y119_SLICE_X1Y119_ALUT (
.I0(CLBLM_R_X3Y119_SLICE_X3Y119_CO6),
.I1(CLBLM_R_X3Y119_SLICE_X2Y119_CO6),
.I2(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLL_L_X2Y119_SLICE_X1Y119_AQ),
.O5(CLBLL_L_X2Y119_SLICE_X1Y119_AO5),
.O6(CLBLL_L_X2Y119_SLICE_X1Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_DO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_CO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_BO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X0Y120_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X0Y120_AO5),
.O6(CLBLL_L_X2Y120_SLICE_X0Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y120_SLICE_X1Y120_AO6),
.Q(CLBLL_L_X2Y120_SLICE_X1Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_DO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_CO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33ff77ff33ff37)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_BLUT (
.I0(LIOB33_X0Y53_IOB_X0Y53_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLL_L_X4Y126_SLICE_X4Y126_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X2Y121_SLICE_X1Y121_B5Q),
.I5(CLBLL_L_X2Y121_SLICE_X0Y121_A5Q),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_BO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ddf0ddf011f0dd)
  ) CLBLL_L_X2Y120_SLICE_X1Y120_ALUT (
.I0(LIOB33_X0Y53_IOB_X0Y53_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X10Y118_SLICE_X13Y118_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y126_SLICE_X4Y126_AQ),
.I5(CLBLL_L_X2Y121_SLICE_X0Y121_A5Q),
.O5(CLBLL_L_X2Y120_SLICE_X1Y120_AO5),
.O6(CLBLL_L_X2Y120_SLICE_X1Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y121_SLICE_X0Y121_BO6),
.Q(CLBLL_L_X2Y121_SLICE_X0Y121_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y121_SLICE_X0Y121_AO6),
.Q(CLBLL_L_X2Y121_SLICE_X0Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y121_SLICE_X1Y121_AO6),
.Q(CLBLL_L_X2Y121_SLICE_X0Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_DO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_CO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30fc30ffff5f5f)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y126_SLICE_X4Y126_AQ),
.I3(CLBLL_L_X4Y121_SLICE_X5Y121_BQ),
.I4(CLBLL_L_X2Y121_SLICE_X0Y121_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_BO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaafcfcfcfc)
  ) CLBLL_L_X2Y121_SLICE_X0Y121_ALUT (
.I0(LIOB33_X0Y79_IOB_X0Y79_I),
.I1(CLBLM_R_X5Y127_SLICE_X7Y127_BQ),
.I2(CLBLL_L_X2Y121_SLICE_X0Y121_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X2Y121_SLICE_X0Y121_AO5),
.O6(CLBLL_L_X2Y121_SLICE_X0Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y121_SLICE_X1Y121_BO5),
.Q(CLBLL_L_X2Y121_SLICE_X1Y121_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y121_SLICE_X1Y121_BO6),
.Q(CLBLL_L_X2Y121_SLICE_X1Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f050d050d0)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_DLUT (
.I0(CLBLM_R_X5Y127_SLICE_X7Y127_BQ),
.I1(CLBLM_R_X3Y123_SLICE_X3Y123_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLL_L_X4Y120_SLICE_X4Y120_CQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y121_SLICE_X2Y121_CQ),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_DO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccffffeceeffff)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_CLUT (
.I0(CLBLM_R_X5Y127_SLICE_X7Y127_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y120_SLICE_X4Y120_CQ),
.I3(CLBLM_R_X3Y123_SLICE_X3Y123_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X3Y121_SLICE_X2Y121_CQ),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_CO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33cc00b8b8b8b8)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_BLUT (
.I0(CLBLM_R_X3Y122_SLICE_X2Y122_A5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X2Y120_SLICE_X1Y120_AQ),
.I3(CLBLL_L_X2Y122_SLICE_X1Y122_BQ),
.I4(CLBLL_L_X4Y123_SLICE_X5Y123_AQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_BO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0ead5aaffaaff)
  ) CLBLL_L_X2Y121_SLICE_X1Y121_ALUT (
.I0(CLBLM_R_X11Y120_SLICE_X14Y120_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y123_SLICE_X5Y123_B5Q),
.I3(CLBLL_L_X2Y121_SLICE_X0Y121_BQ),
.I4(CLBLL_L_X2Y121_SLICE_X1Y121_CO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y121_SLICE_X1Y121_AO5),
.O6(CLBLL_L_X2Y121_SLICE_X1Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X0Y122_DO5),
.O6(CLBLL_L_X2Y122_SLICE_X0Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X0Y122_CO5),
.O6(CLBLL_L_X2Y122_SLICE_X0Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X0Y122_BO5),
.O6(CLBLL_L_X2Y122_SLICE_X0Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y122_SLICE_X0Y122_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X0Y122_AO5),
.O6(CLBLL_L_X2Y122_SLICE_X0Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y122_SLICE_X1Y122_AO5),
.Q(CLBLL_L_X2Y122_SLICE_X1Y122_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y122_SLICE_X1Y122_AO6),
.Q(CLBLL_L_X2Y122_SLICE_X1Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y122_SLICE_X1Y122_BO6),
.Q(CLBLL_L_X2Y122_SLICE_X1Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X1Y122_DO5),
.O6(CLBLL_L_X2Y122_SLICE_X1Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffa)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_CLUT (
.I0(CLBLL_L_X2Y122_SLICE_X1Y122_A5Q),
.I1(1'b1),
.I2(CLBLL_L_X4Y123_SLICE_X5Y123_B5Q),
.I3(CLBLM_R_X3Y125_SLICE_X2Y125_CO6),
.I4(CLBLM_R_X3Y126_SLICE_X2Y126_A5Q),
.I5(CLBLM_R_X5Y125_SLICE_X6Y125_A5Q),
.O5(CLBLL_L_X2Y122_SLICE_X1Y122_CO5),
.O6(CLBLL_L_X2Y122_SLICE_X1Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeaa5400fefe5454)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X2Y122_SLICE_X1Y122_BQ),
.I2(CLBLM_R_X3Y121_SLICE_X3Y121_AQ),
.I3(CLBLM_R_X11Y120_SLICE_X14Y120_DO6),
.I4(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.I5(CLBLM_R_X7Y123_SLICE_X9Y123_A5Q),
.O5(CLBLL_L_X2Y122_SLICE_X1Y122_BO5),
.O6(CLBLL_L_X2Y122_SLICE_X1Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00f0aaf0aa)
  ) CLBLL_L_X2Y122_SLICE_X1Y122_ALUT (
.I0(CLBLL_L_X4Y123_SLICE_X4Y123_BQ),
.I1(CLBLM_R_X3Y120_SLICE_X2Y120_AQ),
.I2(CLBLL_L_X2Y122_SLICE_X1Y122_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y127_IOB_X1Y127_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y122_SLICE_X1Y122_AO5),
.O6(CLBLL_L_X2Y122_SLICE_X1Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y125_SLICE_X0Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X0Y125_DO5),
.O6(CLBLL_L_X2Y125_SLICE_X0Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y125_SLICE_X0Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X0Y125_CO5),
.O6(CLBLL_L_X2Y125_SLICE_X0Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y125_SLICE_X0Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X0Y125_BO5),
.O6(CLBLL_L_X2Y125_SLICE_X0Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y125_SLICE_X0Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X0Y125_AO5),
.O6(CLBLL_L_X2Y125_SLICE_X0Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y125_SLICE_X1Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y125_SLICE_X1Y125_AO6),
.Q(CLBLL_L_X2Y125_SLICE_X1Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y125_SLICE_X1Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y125_SLICE_X1Y125_BO6),
.Q(CLBLL_L_X2Y125_SLICE_X1Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffefffe)
  ) CLBLL_L_X2Y125_SLICE_X1Y125_DLUT (
.I0(CLBLL_L_X2Y121_SLICE_X1Y121_BQ),
.I1(CLBLM_R_X3Y126_SLICE_X2Y126_A5Q),
.I2(CLBLM_R_X5Y125_SLICE_X6Y125_A5Q),
.I3(CLBLL_L_X4Y123_SLICE_X5Y123_B5Q),
.I4(1'b1),
.I5(CLBLL_L_X2Y122_SLICE_X1Y122_A5Q),
.O5(CLBLL_L_X2Y125_SLICE_X1Y125_DO5),
.O6(CLBLL_L_X2Y125_SLICE_X1Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffbfbff003300)
  ) CLBLL_L_X2Y125_SLICE_X1Y125_CLUT (
.I0(RIOB33_X105Y127_IOB_X1Y128_I),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(CLBLL_L_X4Y126_SLICE_X4Y126_DO6),
.I3(CLBLL_L_X4Y125_SLICE_X4Y125_CQ),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X1Y125_CO5),
.O6(CLBLL_L_X2Y125_SLICE_X1Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdf80d08fdf80d08)
  ) CLBLL_L_X2Y125_SLICE_X1Y125_BLUT (
.I0(CLBLL_L_X2Y119_SLICE_X1Y119_BO6),
.I1(CLBLL_L_X2Y125_SLICE_X1Y125_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X2Y121_SLICE_X1Y121_BQ),
.I4(CLBLM_R_X3Y123_SLICE_X2Y123_CQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y125_SLICE_X1Y125_BO5),
.O6(CLBLL_L_X2Y125_SLICE_X1Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000caaaa00c0)
  ) CLBLL_L_X2Y125_SLICE_X1Y125_ALUT (
.I0(CLBLM_R_X5Y120_SLICE_X7Y120_A5Q),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLL_L_X2Y125_SLICE_X1Y125_AQ),
.I3(CLBLL_L_X2Y118_SLICE_X1Y118_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X3Y130_SLICE_X2Y130_AO5),
.O5(CLBLL_L_X2Y125_SLICE_X1Y125_AO5),
.O6(CLBLL_L_X2Y125_SLICE_X1Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y126_SLICE_X0Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y126_SLICE_X0Y126_DO5),
.O6(CLBLL_L_X2Y126_SLICE_X0Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccfc444444f4)
  ) CLBLL_L_X2Y126_SLICE_X0Y126_CLUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(CLBLM_R_X3Y124_SLICE_X2Y124_A5Q),
.I2(LIOB33_X0Y65_IOB_X0Y65_I),
.I3(CLBLL_L_X2Y130_SLICE_X0Y130_BO6),
.I4(CLBLL_L_X2Y130_SLICE_X0Y130_CO6),
.I5(RIOB33_X105Y129_IOB_X1Y129_I),
.O5(CLBLL_L_X2Y126_SLICE_X0Y126_CO5),
.O6(CLBLL_L_X2Y126_SLICE_X0Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5050dcdcff50ffdc)
  ) CLBLL_L_X2Y126_SLICE_X0Y126_BLUT (
.I0(CLBLL_L_X2Y128_SLICE_X0Y128_BO5),
.I1(CLBLL_L_X2Y125_SLICE_X1Y125_BQ),
.I2(LIOB33_X0Y57_IOB_X0Y57_I),
.I3(CLBLM_R_X5Y128_SLICE_X6Y128_A5Q),
.I4(CLBLL_L_X2Y126_SLICE_X0Y126_AO6),
.I5(CLBLL_L_X2Y126_SLICE_X0Y126_AO5),
.O5(CLBLL_L_X2Y126_SLICE_X0Y126_BO5),
.O6(CLBLL_L_X2Y126_SLICE_X0Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffbffbfffff)
  ) CLBLL_L_X2Y126_SLICE_X0Y126_ALUT (
.I0(CLBLL_L_X2Y130_SLICE_X0Y130_CO6),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y126_SLICE_X0Y126_AO5),
.O6(CLBLL_L_X2Y126_SLICE_X0Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y126_SLICE_X1Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y126_SLICE_X1Y126_AO6),
.Q(CLBLL_L_X2Y126_SLICE_X1Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff0f00afaa)
  ) CLBLL_L_X2Y126_SLICE_X1Y126_DLUT (
.I0(RIOB33_X105Y117_IOB_X1Y117_I),
.I1(1'b1),
.I2(CLBLL_L_X2Y128_SLICE_X0Y128_BO5),
.I3(LIOB33_X0Y57_IOB_X0Y58_I),
.I4(CLBLM_R_X3Y129_SLICE_X3Y129_AO5),
.I5(CLBLL_L_X2Y126_SLICE_X1Y126_BO6),
.O5(CLBLL_L_X2Y126_SLICE_X1Y126_DO5),
.O6(CLBLL_L_X2Y126_SLICE_X1Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000ac00000000)
  ) CLBLL_L_X2Y126_SLICE_X1Y126_CLUT (
.I0(CLBLM_R_X3Y123_SLICE_X2Y123_BQ),
.I1(CLBLM_R_X3Y122_SLICE_X2Y122_AQ),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.I4(CLBLL_L_X2Y128_SLICE_X1Y128_BO5),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLL_L_X2Y126_SLICE_X1Y126_CO5),
.O6(CLBLL_L_X2Y126_SLICE_X1Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccdcffff00500050)
  ) CLBLL_L_X2Y126_SLICE_X1Y126_BLUT (
.I0(CLBLL_L_X2Y130_SLICE_X0Y130_CO6),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I3(CLBLL_L_X2Y130_SLICE_X0Y130_AO6),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(CLBLM_R_X3Y124_SLICE_X2Y124_BQ),
.O5(CLBLL_L_X2Y126_SLICE_X1Y126_BO5),
.O6(CLBLL_L_X2Y126_SLICE_X1Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd5c0eac0eac0eac0)
  ) CLBLL_L_X2Y126_SLICE_X1Y126_ALUT (
.I0(CLBLL_L_X2Y126_SLICE_X1Y126_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X2Y121_SLICE_X1Y121_BQ),
.I3(CLBLM_R_X3Y132_SLICE_X2Y132_CO5),
.I4(CLBLL_L_X2Y125_SLICE_X1Y125_AQ),
.I5(CLBLM_R_X3Y130_SLICE_X2Y130_AO5),
.O5(CLBLL_L_X2Y126_SLICE_X1Y126_AO5),
.O6(CLBLL_L_X2Y126_SLICE_X1Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdcdcdcdcffdcffdc)
  ) CLBLL_L_X2Y127_SLICE_X0Y127_DLUT (
.I0(CLBLL_L_X2Y128_SLICE_X0Y128_AO6),
.I1(CLBLL_L_X2Y126_SLICE_X1Y126_CO6),
.I2(CLBLM_R_X3Y124_SLICE_X2Y124_DQ),
.I3(CLBLL_L_X2Y122_SLICE_X1Y122_BQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y129_SLICE_X4Y129_BO6),
.O5(CLBLL_L_X2Y127_SLICE_X0Y127_DO5),
.O6(CLBLL_L_X2Y127_SLICE_X0Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbbfbffffaafa)
  ) CLBLL_L_X2Y127_SLICE_X0Y127_CLUT (
.I0(CLBLM_R_X3Y126_SLICE_X3Y126_BO6),
.I1(CLBLL_L_X2Y128_SLICE_X0Y128_AO5),
.I2(CLBLL_L_X2Y129_SLICE_X1Y129_DO6),
.I3(CLBLL_L_X2Y129_SLICE_X0Y129_CO6),
.I4(CLBLL_L_X2Y127_SLICE_X0Y127_DO6),
.I5(CLBLM_R_X5Y126_SLICE_X6Y126_BQ),
.O5(CLBLL_L_X2Y127_SLICE_X0Y127_CO5),
.O6(CLBLL_L_X2Y127_SLICE_X0Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000200000000)
  ) CLBLL_L_X2Y127_SLICE_X0Y127_BLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_R_X5Y126_SLICE_X6Y126_BQ),
.O5(CLBLL_L_X2Y127_SLICE_X0Y127_BO5),
.O6(CLBLL_L_X2Y127_SLICE_X0Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffafefaaee)
  ) CLBLL_L_X2Y127_SLICE_X0Y127_ALUT (
.I0(CLBLL_L_X2Y127_SLICE_X0Y127_BO6),
.I1(CLBLL_L_X2Y122_SLICE_X1Y122_BQ),
.I2(CLBLL_L_X2Y128_SLICE_X0Y128_AO6),
.I3(CLBLL_L_X4Y129_SLICE_X4Y129_BO6),
.I4(CLBLM_R_X3Y124_SLICE_X2Y124_DQ),
.I5(CLBLL_L_X2Y126_SLICE_X1Y126_CO6),
.O5(CLBLL_L_X2Y127_SLICE_X0Y127_AO5),
.O6(CLBLL_L_X2Y127_SLICE_X0Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h030300000f030f00)
  ) CLBLL_L_X2Y127_SLICE_X1Y127_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y130_SLICE_X0Y130_BO6),
.I2(CLBLL_L_X2Y130_SLICE_X0Y130_CO6),
.I3(CLBLM_R_X7Y127_SLICE_X8Y127_DQ),
.I4(LIOB33_X0Y67_IOB_X0Y67_I),
.I5(CLBLL_L_X2Y130_SLICE_X0Y130_AO6),
.O5(CLBLL_L_X2Y127_SLICE_X1Y127_DO5),
.O6(CLBLL_L_X2Y127_SLICE_X1Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffb)
  ) CLBLL_L_X2Y127_SLICE_X1Y127_CLUT (
.I0(CLBLL_L_X2Y127_SLICE_X1Y127_AO6),
.I1(CLBLL_L_X2Y129_SLICE_X1Y129_BO6),
.I2(CLBLL_L_X4Y125_SLICE_X5Y125_CO6),
.I3(CLBLL_L_X2Y129_SLICE_X1Y129_AO6),
.I4(CLBLL_L_X2Y127_SLICE_X0Y127_AO6),
.I5(CLBLM_R_X3Y126_SLICE_X3Y126_BO6),
.O5(CLBLL_L_X2Y127_SLICE_X1Y127_CO5),
.O6(CLBLL_L_X2Y127_SLICE_X1Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000550030307530)
  ) CLBLL_L_X2Y127_SLICE_X1Y127_BLUT (
.I0(CLBLL_L_X2Y128_SLICE_X1Y128_AO6),
.I1(CLBLL_L_X2Y130_SLICE_X0Y130_BO6),
.I2(CLBLM_R_X3Y125_SLICE_X3Y125_BQ),
.I3(CLBLM_R_X3Y122_SLICE_X3Y122_BQ),
.I4(CLBLL_L_X2Y130_SLICE_X0Y130_CO5),
.I5(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.O5(CLBLL_L_X2Y127_SLICE_X1Y127_BO5),
.O6(CLBLL_L_X2Y127_SLICE_X1Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffefffffffee)
  ) CLBLL_L_X2Y127_SLICE_X1Y127_ALUT (
.I0(CLBLL_L_X2Y127_SLICE_X1Y127_DO6),
.I1(CLBLM_R_X3Y127_SLICE_X2Y127_AO6),
.I2(CLBLM_R_X3Y129_SLICE_X3Y129_AO6),
.I3(CLBLL_L_X2Y127_SLICE_X1Y127_BO6),
.I4(CLBLM_R_X3Y126_SLICE_X2Y126_CO6),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLL_L_X2Y127_SLICE_X1Y127_AO5),
.O6(CLBLL_L_X2Y127_SLICE_X1Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0030003000ba00ba)
  ) CLBLL_L_X2Y128_SLICE_X0Y128_DLUT (
.I0(CLBLL_L_X2Y119_SLICE_X1Y119_AQ),
.I1(CLBLL_L_X2Y130_SLICE_X0Y130_BO6),
.I2(LIOB33_X0Y59_IOB_X0Y59_I),
.I3(CLBLL_L_X2Y130_SLICE_X0Y130_CO6),
.I4(1'b1),
.I5(CLBLL_L_X2Y130_SLICE_X0Y130_AO6),
.O5(CLBLL_L_X2Y128_SLICE_X0Y128_DO5),
.O6(CLBLL_L_X2Y128_SLICE_X0Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff05007777)
  ) CLBLL_L_X2Y128_SLICE_X0Y128_CLUT (
.I0(CLBLL_L_X2Y130_SLICE_X1Y130_AO6),
.I1(CLBLL_L_X2Y128_SLICE_X1Y128_AO5),
.I2(CLBLL_L_X2Y130_SLICE_X0Y130_CO6),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.I5(CLBLL_L_X2Y118_SLICE_X1Y118_CO6),
.O5(CLBLL_L_X2Y128_SLICE_X0Y128_CO5),
.O6(CLBLL_L_X2Y128_SLICE_X0Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffbfffffbfff)
  ) CLBLL_L_X2Y128_SLICE_X0Y128_BLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(CLBLL_L_X2Y130_SLICE_X0Y130_CO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y128_SLICE_X0Y128_BO5),
.O6(CLBLL_L_X2Y128_SLICE_X0Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffdfffffffffffb)
  ) CLBLL_L_X2Y128_SLICE_X0Y128_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y128_SLICE_X0Y128_AO5),
.O6(CLBLL_L_X2Y128_SLICE_X0Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0400000004030003)
  ) CLBLL_L_X2Y128_SLICE_X1Y128_DLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(CLBLL_L_X4Y130_SLICE_X4Y130_AO5),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(CLBLL_L_X2Y130_SLICE_X1Y130_AO5),
.I5(CLBLL_L_X2Y128_SLICE_X1Y128_BO6),
.O5(CLBLL_L_X2Y128_SLICE_X1Y128_DO5),
.O6(CLBLL_L_X2Y128_SLICE_X1Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h111f1111000f0000)
  ) CLBLL_L_X2Y128_SLICE_X1Y128_CLUT (
.I0(CLBLL_L_X2Y128_SLICE_X1Y128_AO6),
.I1(CLBLL_L_X2Y130_SLICE_X0Y130_CO6),
.I2(CLBLL_L_X2Y130_SLICE_X0Y130_CO5),
.I3(CLBLL_L_X2Y128_SLICE_X1Y128_AO5),
.I4(RIOB33_X105Y113_IOB_X1Y114_I),
.I5(CLBLM_R_X5Y127_SLICE_X7Y127_CQ),
.O5(CLBLL_L_X2Y128_SLICE_X1Y128_CO5),
.O6(CLBLL_L_X2Y128_SLICE_X1Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff33ffff00ff)
  ) CLBLL_L_X2Y128_SLICE_X1Y128_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(1'b1),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y128_SLICE_X1Y128_BO5),
.O6(CLBLL_L_X2Y128_SLICE_X1Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcfffffffff3ff)
  ) CLBLL_L_X2Y128_SLICE_X1Y128_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y128_SLICE_X1Y128_AO5),
.O6(CLBLL_L_X2Y128_SLICE_X1Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000003300f3f0)
  ) CLBLL_L_X2Y129_SLICE_X0Y129_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y128_SLICE_X1Y128_AO5),
.I2(LIOB33_X0Y53_IOB_X0Y54_I),
.I3(LIOB33_X0Y69_IOB_X0Y70_I),
.I4(CLBLL_L_X2Y130_SLICE_X1Y130_BO5),
.I5(CLBLL_L_X2Y130_SLICE_X0Y130_CO6),
.O5(CLBLL_L_X2Y129_SLICE_X0Y129_DO5),
.O6(CLBLL_L_X2Y129_SLICE_X0Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000004000000)
  ) CLBLL_L_X2Y129_SLICE_X0Y129_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(RIOB33_X105Y129_IOB_X1Y130_I),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(CLBLL_L_X2Y130_SLICE_X1Y130_AO5),
.I5(CLBLL_L_X2Y118_SLICE_X1Y118_CO6),
.O5(CLBLL_L_X2Y129_SLICE_X0Y129_CO5),
.O6(CLBLL_L_X2Y129_SLICE_X0Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0a000c0c0800)
  ) CLBLL_L_X2Y129_SLICE_X0Y129_BLUT (
.I0(CLBLL_L_X2Y130_SLICE_X0Y130_BO5),
.I1(CLBLL_L_X2Y130_SLICE_X0Y130_AO6),
.I2(CLBLL_L_X2Y118_SLICE_X1Y118_CO6),
.I3(CLBLL_L_X2Y130_SLICE_X0Y130_BO6),
.I4(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.I5(CLBLL_L_X2Y130_SLICE_X0Y130_CO6),
.O5(CLBLL_L_X2Y129_SLICE_X0Y129_BO5),
.O6(CLBLL_L_X2Y129_SLICE_X0Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdffffff02010000)
  ) CLBLL_L_X2Y129_SLICE_X0Y129_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLL_L_X2Y130_SLICE_X0Y130_CO5),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y129_SLICE_X0Y129_AO5),
.O6(CLBLL_L_X2Y129_SLICE_X0Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0004000000000000)
  ) CLBLL_L_X2Y129_SLICE_X1Y129_DLUT (
.I0(CLBLL_L_X2Y128_SLICE_X0Y128_CO6),
.I1(CLBLL_L_X4Y129_SLICE_X4Y129_BO6),
.I2(CLBLL_L_X2Y130_SLICE_X1Y130_CO6),
.I3(CLBLL_L_X2Y130_SLICE_X0Y130_AO5),
.I4(CLBLL_L_X2Y129_SLICE_X0Y129_AO6),
.I5(CLBLM_R_X3Y130_SLICE_X2Y130_BO6),
.O5(CLBLL_L_X2Y129_SLICE_X1Y129_DO5),
.O6(CLBLL_L_X2Y129_SLICE_X1Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000020)
  ) CLBLL_L_X2Y129_SLICE_X1Y129_CLUT (
.I0(CLBLL_L_X2Y129_SLICE_X0Y129_BO6),
.I1(CLBLL_L_X2Y129_SLICE_X0Y129_AO5),
.I2(CLBLM_R_X3Y129_SLICE_X3Y129_AO5),
.I3(CLBLM_R_X3Y130_SLICE_X3Y130_AO5),
.I4(CLBLL_L_X2Y128_SLICE_X1Y128_DO6),
.I5(CLBLL_L_X2Y130_SLICE_X1Y130_CO6),
.O5(CLBLL_L_X2Y129_SLICE_X1Y129_CO5),
.O6(CLBLL_L_X2Y129_SLICE_X1Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffbffffffffff)
  ) CLBLL_L_X2Y129_SLICE_X1Y129_BLUT (
.I0(CLBLM_R_X3Y130_SLICE_X3Y130_AO5),
.I1(CLBLL_L_X4Y129_SLICE_X4Y129_BO6),
.I2(CLBLL_L_X2Y128_SLICE_X0Y128_CO6),
.I3(CLBLM_R_X3Y130_SLICE_X2Y130_BO6),
.I4(CLBLL_L_X2Y130_SLICE_X1Y130_CO6),
.I5(CLBLL_L_X2Y129_SLICE_X0Y129_AO6),
.O5(CLBLL_L_X2Y129_SLICE_X1Y129_BO5),
.O6(CLBLL_L_X2Y129_SLICE_X1Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000004)
  ) CLBLL_L_X2Y129_SLICE_X1Y129_ALUT (
.I0(CLBLL_L_X2Y129_SLICE_X0Y129_AO5),
.I1(CLBLM_R_X3Y130_SLICE_X2Y130_BO6),
.I2(CLBLL_L_X2Y129_SLICE_X0Y129_CO6),
.I3(CLBLL_L_X2Y130_SLICE_X1Y130_CO6),
.I4(CLBLL_L_X2Y128_SLICE_X0Y128_CO6),
.I5(CLBLL_L_X2Y130_SLICE_X0Y130_AO5),
.O5(CLBLL_L_X2Y129_SLICE_X1Y129_AO5),
.O6(CLBLL_L_X2Y129_SLICE_X1Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000004400500000)
  ) CLBLL_L_X2Y130_SLICE_X0Y130_DLUT (
.I0(CLBLL_L_X2Y131_SLICE_X1Y131_AO6),
.I1(LIOB33_X0Y55_IOB_X0Y55_I),
.I2(LIOB33_X0Y61_IOB_X0Y61_I),
.I3(CLBLL_L_X2Y130_SLICE_X0Y130_CO6),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(RIOB33_X105Y133_IOB_X1Y134_I),
.O5(CLBLL_L_X2Y130_SLICE_X0Y130_DO5),
.O6(CLBLL_L_X2Y130_SLICE_X0Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffefffffffffffbf)
  ) CLBLL_L_X2Y130_SLICE_X0Y130_CLUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(RIOB33_X105Y135_IOB_X1Y136_I),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(RIOB33_X105Y129_IOB_X1Y130_I),
.I4(RIOB33_X105Y135_IOB_X1Y135_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y130_SLICE_X0Y130_CO5),
.O6(CLBLL_L_X2Y130_SLICE_X0Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfffbffffbddfbdd)
  ) CLBLL_L_X2Y130_SLICE_X0Y130_BLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y130_SLICE_X0Y130_BO5),
.O6(CLBLL_L_X2Y130_SLICE_X0Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdfffdf0000c000)
  ) CLBLL_L_X2Y130_SLICE_X0Y130_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(CLBLL_L_X2Y130_SLICE_X0Y130_CO5),
.I5(1'b1),
.O5(CLBLL_L_X2Y130_SLICE_X0Y130_AO5),
.O6(CLBLL_L_X2Y130_SLICE_X0Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y130_SLICE_X1Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y130_SLICE_X1Y130_DO5),
.O6(CLBLL_L_X2Y130_SLICE_X1Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000010103c03d0d0)
  ) CLBLL_L_X2Y130_SLICE_X1Y130_CLUT (
.I0(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(CLBLL_L_X2Y130_SLICE_X0Y130_CO6),
.O5(CLBLL_L_X2Y130_SLICE_X1Y130_CO5),
.O6(CLBLL_L_X2Y130_SLICE_X1Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbffffffff77ffff)
  ) CLBLL_L_X2Y130_SLICE_X1Y130_BLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(CLBLL_L_X2Y130_SLICE_X0Y130_CO6),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y130_SLICE_X1Y130_BO5),
.O6(CLBLL_L_X2Y130_SLICE_X1Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffddffdd44004400)
  ) CLBLL_L_X2Y130_SLICE_X1Y130_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(1'b1),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y130_SLICE_X1Y130_AO5),
.O6(CLBLL_L_X2Y130_SLICE_X1Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X0Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X0Y131_DO5),
.O6(CLBLL_L_X2Y131_SLICE_X0Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X0Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X0Y131_CO5),
.O6(CLBLL_L_X2Y131_SLICE_X0Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X0Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X0Y131_BO5),
.O6(CLBLL_L_X2Y131_SLICE_X0Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X0Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X0Y131_AO5),
.O6(CLBLL_L_X2Y131_SLICE_X0Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X1Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X1Y131_DO5),
.O6(CLBLL_L_X2Y131_SLICE_X1Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X1Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X1Y131_CO5),
.O6(CLBLL_L_X2Y131_SLICE_X1Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y131_SLICE_X1Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X1Y131_BO5),
.O6(CLBLL_L_X2Y131_SLICE_X1Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffffff00ffffff)
  ) CLBLL_L_X2Y131_SLICE_X1Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y131_SLICE_X1Y131_AO5),
.O6(CLBLL_L_X2Y131_SLICE_X1Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y132_SLICE_X0Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y132_SLICE_X0Y132_DO5),
.O6(CLBLL_L_X2Y132_SLICE_X0Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y132_SLICE_X0Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y132_SLICE_X0Y132_CO5),
.O6(CLBLL_L_X2Y132_SLICE_X0Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y132_SLICE_X0Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y132_SLICE_X0Y132_BO5),
.O6(CLBLL_L_X2Y132_SLICE_X0Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y132_SLICE_X0Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y132_SLICE_X0Y132_AO5),
.O6(CLBLL_L_X2Y132_SLICE_X0Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y132_SLICE_X1Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y132_SLICE_X1Y132_DO5),
.O6(CLBLL_L_X2Y132_SLICE_X1Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y132_SLICE_X1Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y132_SLICE_X1Y132_CO5),
.O6(CLBLL_L_X2Y132_SLICE_X1Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y132_SLICE_X1Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y132_SLICE_X1Y132_BO5),
.O6(CLBLL_L_X2Y132_SLICE_X1Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLL_L_X2Y132_SLICE_X1Y132_ALUT (
.I0(CLBLM_R_X3Y132_SLICE_X2Y132_A5Q),
.I1(CLBLM_R_X3Y123_SLICE_X2Y123_CQ),
.I2(CLBLM_R_X3Y129_SLICE_X2Y129_AQ),
.I3(CLBLM_R_X3Y132_SLICE_X2Y132_BQ),
.I4(CLBLM_R_X3Y131_SLICE_X2Y131_BQ),
.I5(CLBLM_R_X3Y131_SLICE_X2Y131_AQ),
.O5(CLBLL_L_X2Y132_SLICE_X1Y132_AO5),
.O6(CLBLL_L_X2Y132_SLICE_X1Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y117_SLICE_X4Y117_AO6),
.Q(CLBLL_L_X4Y117_SLICE_X4Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_DO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_CO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_BO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888b88ff000000)
  ) CLBLL_L_X4Y117_SLICE_X4Y117_ALUT (
.I0(CLBLL_L_X4Y122_SLICE_X4Y122_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y117_SLICE_X5Y117_CO6),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y117_SLICE_X4Y117_AO5),
.O6(CLBLL_L_X4Y117_SLICE_X4Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y117_SLICE_X5Y117_AO6),
.Q(CLBLL_L_X4Y117_SLICE_X5Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y117_SLICE_X5Y117_BO6),
.Q(CLBLL_L_X4Y117_SLICE_X5Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_DO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055005500500055)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_CLUT (
.I0(CLBLL_L_X4Y117_SLICE_X4Y117_AQ),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X3Y123_SLICE_X2Y123_DQ),
.I4(CLBLL_L_X4Y126_SLICE_X4Y126_DO6),
.I5(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_CO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000faaaf888)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_BLUT (
.I0(CLBLL_L_X4Y119_SLICE_X5Y119_DO6),
.I1(CLBLL_L_X4Y117_SLICE_X5Y117_BQ),
.I2(CLBLM_R_X3Y124_SLICE_X2Y124_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y116_SLICE_X7Y116_DO5),
.I5(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_BO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fffc000000fc)
  ) CLBLL_L_X4Y117_SLICE_X5Y117_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y117_SLICE_X6Y117_AQ),
.I2(CLBLL_L_X4Y117_SLICE_X5Y117_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y118_SLICE_X7Y118_DO6),
.I5(CLBLL_L_X4Y118_SLICE_X5Y118_CQ),
.O5(CLBLL_L_X4Y117_SLICE_X5Y117_AO5),
.O6(CLBLL_L_X4Y117_SLICE_X5Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y118_SLICE_X4Y118_AO6),
.Q(CLBLL_L_X4Y118_SLICE_X4Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_DO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_CO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_BO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff44ff4000440040)
  ) CLBLL_L_X4Y118_SLICE_X4Y118_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I2(CLBLL_L_X4Y118_SLICE_X4Y118_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y118_SLICE_X13Y118_AQ),
.I5(CLBLL_L_X2Y118_SLICE_X1Y118_A5Q),
.O5(CLBLL_L_X4Y118_SLICE_X4Y118_AO5),
.O6(CLBLL_L_X4Y118_SLICE_X4Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y118_SLICE_X5Y118_CO5),
.Q(CLBLL_L_X4Y118_SLICE_X5Y118_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y118_SLICE_X5Y118_AO6),
.Q(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y118_SLICE_X5Y118_BO6),
.Q(CLBLL_L_X4Y118_SLICE_X5Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y118_SLICE_X5Y118_CO6),
.Q(CLBLL_L_X4Y118_SLICE_X5Y118_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_DO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0dddd8888)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_DQ),
.I3(1'b1),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_CO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fbfc0000bbcc)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_BLUT (
.I0(CLBLM_R_X3Y119_SLICE_X3Y119_BO5),
.I1(CLBLL_L_X4Y118_SLICE_X5Y118_BQ),
.I2(CLBLM_R_X5Y130_SLICE_X7Y130_AQ),
.I3(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I4(CLBLM_R_X5Y118_SLICE_X6Y118_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_BO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88bb88bb88b8b8)
  ) CLBLL_L_X4Y118_SLICE_X5Y118_ALUT (
.I0(CLBLL_L_X4Y120_SLICE_X5Y120_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I3(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I4(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLL_L_X4Y118_SLICE_X5Y118_AO5),
.O6(CLBLL_L_X4Y118_SLICE_X5Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X4Y119_AO6),
.Q(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X4Y119_BO6),
.Q(CLBLL_L_X4Y119_SLICE_X4Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X4Y119_CO6),
.Q(CLBLL_L_X4Y119_SLICE_X4Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X4Y119_DO6),
.Q(CLBLL_L_X4Y119_SLICE_X4Y119_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff303030ff303030)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y120_SLICE_X1Y120_BO6),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_DQ),
.I3(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_DO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0afafa0a0a0a0)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_CLUT (
.I0(CLBLL_L_X4Y122_SLICE_X4Y122_AQ),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_CO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff410041ff000000)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_BLUT (
.I0(CLBLM_L_X8Y123_SLICE_X11Y123_CQ),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_BQ),
.I2(CLBLM_R_X3Y119_SLICE_X3Y119_BO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y120_SLICE_X12Y120_BQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_BO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbba1110bbba1110)
  ) CLBLL_L_X4Y119_SLICE_X4Y119_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y126_SLICE_X7Y126_CO5),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.I3(CLBLM_R_X3Y120_SLICE_X3Y120_BQ),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X4Y119_AO5),
.O6(CLBLL_L_X4Y119_SLICE_X4Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X5Y119_AO6),
.Q(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X5Y119_BO6),
.Q(CLBLL_L_X4Y119_SLICE_X5Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X5Y119_CO6),
.Q(CLBLL_L_X4Y119_SLICE_X5Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00500050aeae0404)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_BQ),
.I4(CLBLM_R_X3Y119_SLICE_X3Y119_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_DO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fc000cfafc0a0c)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_CLUT (
.I0(CLBLL_L_X4Y128_SLICE_X4Y128_AO6),
.I1(CLBLL_L_X4Y119_SLICE_X5Y119_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y117_SLICE_X4Y117_AO5),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_DQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_CO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff008888ff00cccc)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_BLUT (
.I0(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I1(CLBLL_L_X4Y119_SLICE_X5Y119_BQ),
.I2(1'b1),
.I3(CLBLM_R_X3Y121_SLICE_X2Y121_C5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_BO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccffccf0cc00)
  ) CLBLL_L_X4Y119_SLICE_X5Y119_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y117_SLICE_X5Y117_BQ),
.I2(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y126_SLICE_X7Y126_CO5),
.I5(CLBLL_L_X4Y119_SLICE_X4Y119_CQ),
.O5(CLBLL_L_X4Y119_SLICE_X5Y119_AO5),
.O6(CLBLL_L_X4Y119_SLICE_X5Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X8Y123_CO6),
.Q(CLBLL_L_X4Y120_SLICE_X4Y120_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y120_SLICE_X4Y120_CO5),
.Q(CLBLL_L_X4Y120_SLICE_X4Y120_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y120_SLICE_X4Y120_AO6),
.Q(CLBLL_L_X4Y120_SLICE_X4Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y120_SLICE_X4Y120_BO6),
.Q(CLBLL_L_X4Y120_SLICE_X4Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y120_SLICE_X4Y120_CO6),
.Q(CLBLL_L_X4Y120_SLICE_X4Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y120_SLICE_X4Y120_DO6),
.Q(CLBLL_L_X4Y120_SLICE_X4Y120_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hddd88888ddd8ddd8)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y120_SLICE_X4Y120_CQ),
.I2(CLBLL_L_X4Y120_SLICE_X4Y120_DQ),
.I3(CLBLM_R_X3Y121_SLICE_X3Y121_BQ),
.I4(CLBLM_R_X11Y120_SLICE_X14Y120_DO6),
.I5(CLBLM_R_X7Y123_SLICE_X9Y123_A5Q),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_DO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0afa0acfc0cfc0)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_CLUT (
.I0(CLBLM_R_X3Y123_SLICE_X3Y123_CQ),
.I1(CLBLL_L_X4Y120_SLICE_X4Y120_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y120_SLICE_X4Y120_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_CO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccf0003cfcc0300)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X5Y121_SLICE_X7Y121_BO6),
.I4(CLBLL_L_X4Y118_SLICE_X4Y118_AQ),
.I5(CLBLM_R_X5Y122_SLICE_X6Y122_CQ),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_BO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa8ffa8a8a8a8a8)
  ) CLBLL_L_X4Y120_SLICE_X4Y120_ALUT (
.I0(CLBLM_R_X5Y126_SLICE_X7Y126_CO6),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_BQ),
.I2(CLBLL_L_X4Y120_SLICE_X4Y120_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y121_SLICE_X5Y121_CQ),
.O5(CLBLL_L_X4Y120_SLICE_X4Y120_AO5),
.O6(CLBLL_L_X4Y120_SLICE_X4Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y119_SLICE_X5Y119_DO5),
.Q(CLBLL_L_X4Y120_SLICE_X5Y120_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y120_SLICE_X5Y120_AO6),
.Q(CLBLL_L_X4Y120_SLICE_X5Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y120_SLICE_X5Y120_BO6),
.Q(CLBLL_L_X4Y120_SLICE_X5Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y120_SLICE_X5Y120_CO6),
.Q(CLBLL_L_X4Y120_SLICE_X5Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000c0c00000)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_DLUT (
.I0(1'b1),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X5Y123_SLICE_X7Y123_BQ),
.I3(1'b1),
.I4(CLBLM_R_X3Y122_SLICE_X2Y122_CQ),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_DO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe54ae04ff55aa00)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y120_SLICE_X5Y120_CQ),
.I2(CLBLM_R_X11Y120_SLICE_X14Y120_DO6),
.I3(CLBLM_L_X12Y121_SLICE_X16Y121_AQ),
.I4(CLBLM_R_X3Y122_SLICE_X2Y122_CQ),
.I5(CLBLM_R_X7Y123_SLICE_X9Y123_A5Q),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_CO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff006c0000006c)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_BLUT (
.I0(CLBLL_L_X4Y120_SLICE_X5Y120_DO6),
.I1(CLBLL_L_X4Y120_SLICE_X5Y120_BQ),
.I2(CLBLL_L_X4Y120_SLICE_X5Y120_AQ),
.I3(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_CQ),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_BO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff5a005a)
  ) CLBLL_L_X4Y120_SLICE_X5Y120_ALUT (
.I0(CLBLL_L_X4Y120_SLICE_X5Y120_DO6),
.I1(1'b1),
.I2(CLBLL_L_X4Y120_SLICE_X5Y120_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y122_SLICE_X13Y122_AQ),
.I5(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.O5(CLBLL_L_X4Y120_SLICE_X5Y120_AO5),
.O6(CLBLL_L_X4Y120_SLICE_X5Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y121_SLICE_X4Y121_AO6),
.Q(CLBLL_L_X4Y121_SLICE_X4Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y121_SLICE_X4Y121_BO6),
.Q(CLBLL_L_X4Y121_SLICE_X4Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y121_SLICE_X4Y121_CO6),
.Q(CLBLL_L_X4Y121_SLICE_X4Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y121_SLICE_X4Y121_DO6),
.Q(CLBLL_L_X4Y121_SLICE_X4Y121_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8d888d888d888d88)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y121_SLICE_X4Y121_AQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X3Y120_SLICE_X3Y120_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y121_SLICE_X4Y121_DO5),
.O6(CLBLL_L_X4Y121_SLICE_X4Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe54fe54fe54aa00)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y121_SLICE_X4Y121_CQ),
.I2(CLBLM_R_X5Y122_SLICE_X7Y122_CO6),
.I3(CLBLM_R_X3Y121_SLICE_X2Y121_BQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.O5(CLBLL_L_X4Y121_SLICE_X4Y121_CO5),
.O6(CLBLL_L_X4Y121_SLICE_X4Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaaaaaff888888)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_BLUT (
.I0(CLBLM_R_X5Y126_SLICE_X7Y126_CO6),
.I1(CLBLL_L_X4Y121_SLICE_X4Y121_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y118_SLICE_X5Y118_BQ),
.I5(CLBLM_R_X3Y124_SLICE_X3Y124_CQ),
.O5(CLBLL_L_X4Y121_SLICE_X4Y121_BO5),
.O6(CLBLL_L_X4Y121_SLICE_X4Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00e2e2ff00aaaa)
  ) CLBLL_L_X4Y121_SLICE_X4Y121_ALUT (
.I0(CLBLM_R_X5Y122_SLICE_X7Y122_AQ),
.I1(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.I2(CLBLL_L_X4Y121_SLICE_X4Y121_AQ),
.I3(CLBLL_L_X4Y121_SLICE_X4Y121_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y125_SLICE_X4Y125_BQ),
.O5(CLBLL_L_X4Y121_SLICE_X4Y121_AO5),
.O6(CLBLL_L_X4Y121_SLICE_X4Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y121_SLICE_X5Y121_AO6),
.Q(CLBLL_L_X4Y121_SLICE_X5Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y121_SLICE_X5Y121_BO6),
.Q(CLBLL_L_X4Y121_SLICE_X5Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y121_SLICE_X5Y121_CO6),
.Q(CLBLL_L_X4Y121_SLICE_X5Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffeeffee)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_DLUT (
.I0(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.I1(CLBLM_R_X5Y122_SLICE_X6Y122_CQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y119_SLICE_X4Y119_CQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y120_SLICE_X4Y120_BQ),
.O5(CLBLL_L_X4Y121_SLICE_X5Y121_DO5),
.O6(CLBLL_L_X4Y121_SLICE_X5Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffccf0f0aa88)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_CLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLL_L_X4Y121_SLICE_X5Y121_CQ),
.I2(CLBLL_L_X4Y118_SLICE_X5Y118_C5Q),
.I3(CLBLM_R_X5Y121_SLICE_X7Y121_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.O5(CLBLL_L_X4Y121_SLICE_X5Y121_CO5),
.O6(CLBLL_L_X4Y121_SLICE_X5Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf505f000fc0cfc0c)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLL_L_X4Y121_SLICE_X5Y121_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y121_SLICE_X15Y121_AQ),
.I4(CLBLM_R_X3Y128_SLICE_X2Y128_AO6),
.I5(CLBLL_L_X4Y117_SLICE_X4Y117_AO5),
.O5(CLBLL_L_X4Y121_SLICE_X5Y121_BO5),
.O6(CLBLL_L_X4Y121_SLICE_X5Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf088f0bbf0ccf0ff)
  ) CLBLL_L_X4Y121_SLICE_X5Y121_ALUT (
.I0(CLBLL_L_X4Y120_SLICE_X4Y120_CQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y121_SLICE_X2Y121_CQ),
.I5(CLBLM_R_X3Y123_SLICE_X3Y123_CQ),
.O5(CLBLL_L_X4Y121_SLICE_X5Y121_AO5),
.O6(CLBLL_L_X4Y121_SLICE_X5Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y122_SLICE_X4Y122_CO6),
.Q(CLBLL_L_X4Y122_SLICE_X4Y122_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y122_SLICE_X4Y122_AO6),
.Q(CLBLL_L_X4Y122_SLICE_X4Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y122_SLICE_X4Y122_BO6),
.Q(CLBLL_L_X4Y122_SLICE_X4Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y122_SLICE_X4Y122_DO6),
.Q(CLBLL_L_X4Y122_SLICE_X4Y122_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccc0000)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y121_SLICE_X12Y121_DQ),
.I2(CLBLM_R_X3Y123_SLICE_X2Y123_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y122_SLICE_X4Y122_DO5),
.O6(CLBLL_L_X4Y122_SLICE_X4Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8bb8bbbbf000f000)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_CLUT (
.I0(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y123_SLICE_X6Y123_AQ),
.I3(CLBLL_L_X4Y122_SLICE_X4Y122_A5Q),
.I4(CLBLM_R_X5Y124_SLICE_X6Y124_DO5),
.I5(1'b1),
.O5(CLBLL_L_X4Y122_SLICE_X4Y122_CO5),
.O6(CLBLL_L_X4Y122_SLICE_X4Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0d1c0d1d1c0d1c0)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y122_SLICE_X5Y122_C5Q),
.I3(CLBLM_R_X5Y122_SLICE_X7Y122_BQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y122_SLICE_X7Y122_CO6),
.O5(CLBLL_L_X4Y122_SLICE_X4Y122_BO5),
.O6(CLBLL_L_X4Y122_SLICE_X4Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfacc50ccfacc50)
  ) CLBLL_L_X4Y122_SLICE_X4Y122_ALUT (
.I0(CLBLM_R_X5Y126_SLICE_X7Y126_CO5),
.I1(CLBLM_L_X10Y121_SLICE_X12Y121_DQ),
.I2(CLBLL_L_X4Y122_SLICE_X4Y122_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y121_SLICE_X7Y121_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y122_SLICE_X4Y122_AO5),
.O6(CLBLL_L_X4Y122_SLICE_X4Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y122_SLICE_X5Y122_CO5),
.Q(CLBLL_L_X4Y122_SLICE_X5Y122_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y122_SLICE_X5Y122_AO6),
.Q(CLBLL_L_X4Y122_SLICE_X5Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y122_SLICE_X5Y122_BO6),
.Q(CLBLL_L_X4Y122_SLICE_X5Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y122_SLICE_X5Y122_CO6),
.Q(CLBLL_L_X4Y122_SLICE_X5Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y122_SLICE_X5Y122_DO6),
.Q(CLBLL_L_X4Y122_SLICE_X5Y122_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f0f00000)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X8Y123_SLICE_X11Y123_BQ),
.I3(CLBLM_R_X3Y121_SLICE_X3Y121_AQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y122_SLICE_X5Y122_DO5),
.O6(CLBLL_L_X4Y122_SLICE_X5Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00f0fff000)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.I2(CLBLM_R_X5Y122_SLICE_X6Y122_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y122_SLICE_X5Y122_CO5),
.O6(CLBLL_L_X4Y122_SLICE_X5Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbe14aa00ee44aa00)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y122_SLICE_X5Y122_BQ),
.I2(CLBLL_L_X4Y123_SLICE_X5Y123_AQ),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.I4(CLBLM_R_X5Y124_SLICE_X6Y124_DO5),
.I5(CLBLL_L_X4Y123_SLICE_X5Y123_CO5),
.O5(CLBLL_L_X4Y122_SLICE_X5Y122_BO5),
.O6(CLBLL_L_X4Y122_SLICE_X5Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcff00fcfc0000)
  ) CLBLL_L_X4Y122_SLICE_X5Y122_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y122_SLICE_X7Y122_BQ),
.I2(CLBLL_L_X4Y122_SLICE_X5Y122_AQ),
.I3(CLBLM_L_X10Y121_SLICE_X13Y121_B5Q),
.I4(CLBLM_R_X5Y126_SLICE_X7Y126_CO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y122_SLICE_X5Y122_AO5),
.O6(CLBLL_L_X4Y122_SLICE_X5Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y123_SLICE_X4Y123_AO6),
.Q(CLBLL_L_X4Y123_SLICE_X4Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y123_SLICE_X4Y123_BO6),
.Q(CLBLL_L_X4Y123_SLICE_X4Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_DLUT (
.I0(CLBLL_L_X4Y122_SLICE_X4Y122_CO5),
.I1(CLBLL_L_X4Y123_SLICE_X4Y123_AQ),
.I2(CLBLL_L_X4Y123_SLICE_X5Y123_AQ),
.I3(CLBLL_L_X4Y122_SLICE_X5Y122_BQ),
.I4(CLBLL_L_X4Y123_SLICE_X4Y123_BQ),
.I5(CLBLL_L_X4Y124_SLICE_X4Y124_AQ),
.O5(CLBLL_L_X4Y123_SLICE_X4Y123_DO5),
.O6(CLBLL_L_X4Y123_SLICE_X4Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_CLUT (
.I0(CLBLM_R_X5Y123_SLICE_X6Y123_AQ),
.I1(CLBLL_L_X4Y122_SLICE_X4Y122_A5Q),
.I2(CLBLL_L_X4Y123_SLICE_X4Y123_BQ),
.I3(CLBLL_L_X4Y122_SLICE_X5Y122_BQ),
.I4(CLBLL_L_X4Y123_SLICE_X5Y123_AQ),
.I5(CLBLL_L_X4Y124_SLICE_X4Y124_AQ),
.O5(CLBLL_L_X4Y123_SLICE_X4Y123_CO5),
.O6(CLBLL_L_X4Y123_SLICE_X4Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8bbb8888b8888888)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_BLUT (
.I0(CLBLM_R_X5Y124_SLICE_X7Y124_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y122_SLICE_X4Y122_CO5),
.I3(CLBLL_L_X4Y124_SLICE_X4Y124_AQ),
.I4(CLBLM_R_X5Y124_SLICE_X6Y124_DO5),
.I5(CLBLL_L_X4Y123_SLICE_X4Y123_BQ),
.O5(CLBLL_L_X4Y123_SLICE_X4Y123_BO5),
.O6(CLBLL_L_X4Y123_SLICE_X4Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf03cc00fc30cc00)
  ) CLBLL_L_X4Y123_SLICE_X4Y123_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y123_SLICE_X4Y123_AQ),
.I3(CLBLM_R_X7Y129_SLICE_X8Y129_CQ),
.I4(CLBLM_R_X5Y124_SLICE_X6Y124_DO5),
.I5(CLBLL_L_X4Y123_SLICE_X4Y123_CO6),
.O5(CLBLL_L_X4Y123_SLICE_X4Y123_AO5),
.O6(CLBLL_L_X4Y123_SLICE_X4Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y123_SLICE_X5Y123_BO5),
.Q(CLBLL_L_X4Y123_SLICE_X5Y123_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y123_SLICE_X5Y123_AO6),
.Q(CLBLL_L_X4Y123_SLICE_X5Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y123_SLICE_X5Y123_BO6),
.Q(CLBLL_L_X4Y123_SLICE_X5Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f5f3fff1f5f3fff)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_DLUT (
.I0(CLBLL_L_X4Y123_SLICE_X4Y123_AQ),
.I1(CLBLL_L_X4Y122_SLICE_X5Y122_BQ),
.I2(CLBLL_L_X4Y124_SLICE_X4Y124_CQ),
.I3(CLBLL_L_X4Y123_SLICE_X5Y123_AQ),
.I4(CLBLL_L_X4Y124_SLICE_X4Y124_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y123_SLICE_X5Y123_DO5),
.O6(CLBLL_L_X4Y123_SLICE_X5Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff153f80008000)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_CLUT (
.I0(CLBLM_R_X5Y123_SLICE_X6Y123_AQ),
.I1(CLBLL_L_X4Y124_SLICE_X4Y124_AQ),
.I2(CLBLL_L_X4Y123_SLICE_X4Y123_BQ),
.I3(CLBLL_L_X4Y122_SLICE_X4Y122_A5Q),
.I4(CLBLL_L_X4Y123_SLICE_X5Y123_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y123_SLICE_X5Y123_CO5),
.O6(CLBLL_L_X4Y123_SLICE_X5Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1a0b1a0fafa5050)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLL_L_X4Y122_SLICE_X5Y122_BQ),
.I3(CLBLM_R_X5Y125_SLICE_X6Y125_BQ),
.I4(CLBLL_L_X4Y125_SLICE_X5Y125_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y123_SLICE_X5Y123_BO5),
.O6(CLBLL_L_X4Y123_SLICE_X5Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0affa0000a00a0)
  ) CLBLL_L_X4Y123_SLICE_X5Y123_ALUT (
.I0(CLBLM_R_X5Y124_SLICE_X6Y124_DO5),
.I1(1'b1),
.I2(CLBLL_L_X4Y123_SLICE_X5Y123_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y123_SLICE_X5Y123_CO5),
.I5(CLBLL_L_X4Y124_SLICE_X5Y124_CQ),
.O5(CLBLL_L_X4Y123_SLICE_X5Y123_AO5),
.O6(CLBLL_L_X4Y123_SLICE_X5Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X9Y124_BO6),
.Q(CLBLL_L_X4Y124_SLICE_X4Y124_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y124_SLICE_X4Y124_AO6),
.Q(CLBLL_L_X4Y124_SLICE_X4Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y124_SLICE_X4Y124_BO6),
.Q(CLBLL_L_X4Y124_SLICE_X4Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y124_SLICE_X4Y124_CO6),
.Q(CLBLL_L_X4Y124_SLICE_X4Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y124_SLICE_X4Y124_DO6),
.Q(CLBLL_L_X4Y124_SLICE_X4Y124_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa30003000)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_DLUT (
.I0(CLBLM_R_X3Y131_SLICE_X2Y131_AQ),
.I1(CLBLM_R_X5Y124_SLICE_X7Y124_CQ),
.I2(CLBLL_L_X4Y124_SLICE_X4Y124_DQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y124_SLICE_X4Y124_DO5),
.O6(CLBLL_L_X4Y124_SLICE_X4Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f06600cc00)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_CLUT (
.I0(CLBLL_L_X4Y124_SLICE_X4Y124_BQ),
.I1(CLBLL_L_X4Y124_SLICE_X4Y124_CQ),
.I2(CLBLM_R_X3Y123_SLICE_X3Y123_AQ),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_DO5),
.I4(CLBLL_L_X4Y123_SLICE_X4Y123_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y124_SLICE_X4Y124_CO5),
.O6(CLBLL_L_X4Y124_SLICE_X4Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hddcceecc11002200)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_BLUT (
.I0(CLBLL_L_X4Y123_SLICE_X4Y123_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_DO5),
.I4(CLBLL_L_X4Y124_SLICE_X4Y124_BQ),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_CQ),
.O5(CLBLL_L_X4Y124_SLICE_X4Y124_BO5),
.O6(CLBLL_L_X4Y124_SLICE_X4Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff780078ff000000)
  ) CLBLL_L_X4Y124_SLICE_X4Y124_ALUT (
.I0(CLBLM_R_X5Y123_SLICE_X6Y123_AQ),
.I1(CLBLL_L_X4Y122_SLICE_X4Y122_A5Q),
.I2(CLBLL_L_X4Y124_SLICE_X4Y124_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_DO5),
.O5(CLBLL_L_X4Y124_SLICE_X4Y124_AO5),
.O6(CLBLL_L_X4Y124_SLICE_X4Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y124_SLICE_X5Y124_AO6),
.Q(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y124_SLICE_X5Y124_BO6),
.Q(CLBLL_L_X4Y124_SLICE_X5Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y124_SLICE_X5Y124_CO6),
.Q(CLBLL_L_X4Y124_SLICE_X5Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y124_SLICE_X5Y124_DO6),
.Q(CLBLL_L_X4Y124_SLICE_X5Y124_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00e4e4e4e4)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_DLUT (
.I0(CLBLL_L_X2Y119_SLICE_X1Y119_BO6),
.I1(CLBLL_L_X4Y123_SLICE_X5Y123_B5Q),
.I2(CLBLL_L_X4Y124_SLICE_X5Y124_DQ),
.I3(CLBLL_L_X4Y122_SLICE_X5Y122_DQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y124_SLICE_X5Y124_DO5),
.O6(CLBLL_L_X4Y124_SLICE_X5Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe54fe54ae04ae04)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y124_SLICE_X5Y124_CQ),
.I2(CLBLM_R_X5Y126_SLICE_X7Y126_CO5),
.I3(CLBLM_R_X3Y124_SLICE_X3Y124_BQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_A5Q),
.O5(CLBLL_L_X4Y124_SLICE_X5Y124_CO5),
.O6(CLBLL_L_X4Y124_SLICE_X5Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaf0aaccaacc)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_BLUT (
.I0(CLBLL_L_X4Y122_SLICE_X4Y122_DQ),
.I1(CLBLL_L_X4Y124_SLICE_X5Y124_BQ),
.I2(CLBLM_R_X7Y125_SLICE_X8Y125_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X10Y129_SLICE_X13Y129_DO6),
.O5(CLBLL_L_X4Y124_SLICE_X5Y124_BO5),
.O6(CLBLL_L_X4Y124_SLICE_X5Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbea5140ffaa5500)
  ) CLBLL_L_X4Y124_SLICE_X5Y124_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.I2(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.I3(CLBLL_L_X4Y120_SLICE_X5Y120_BQ),
.I4(CLBLL_L_X4Y123_SLICE_X4Y123_AQ),
.I5(CLBLL_L_X4Y125_SLICE_X4Y125_BQ),
.O5(CLBLL_L_X4Y124_SLICE_X5Y124_AO5),
.O6(CLBLL_L_X4Y124_SLICE_X5Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y125_SLICE_X4Y125_CO5),
.Q(CLBLL_L_X4Y125_SLICE_X4Y125_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y125_SLICE_X4Y125_AO6),
.Q(CLBLL_L_X4Y125_SLICE_X4Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y125_SLICE_X4Y125_BO6),
.Q(CLBLL_L_X4Y125_SLICE_X4Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y125_SLICE_X4Y125_CO6),
.Q(CLBLL_L_X4Y125_SLICE_X4Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7350ffff73507350)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_DLUT (
.I0(CLBLL_L_X4Y126_SLICE_X4Y126_CO5),
.I1(CLBLL_L_X2Y129_SLICE_X0Y129_AO6),
.I2(CLBLM_L_X10Y121_SLICE_X12Y121_C5Q),
.I3(CLBLL_L_X4Y121_SLICE_X4Y121_AQ),
.I4(CLBLL_L_X4Y126_SLICE_X4Y126_BO6),
.I5(CLBLM_R_X3Y125_SLICE_X3Y125_AQ),
.O5(CLBLL_L_X4Y125_SLICE_X4Y125_DO5),
.O6(CLBLL_L_X4Y125_SLICE_X4Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccf0aaf0aa)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_CLUT (
.I0(CLBLM_R_X3Y130_SLICE_X3Y130_BO6),
.I1(CLBLL_L_X2Y127_SLICE_X0Y127_CO6),
.I2(CLBLM_R_X3Y123_SLICE_X3Y123_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y125_SLICE_X4Y125_CO5),
.O6(CLBLL_L_X4Y125_SLICE_X4Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff030003ff030003)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.I2(CLBLM_R_X3Y124_SLICE_X3Y124_C5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y125_SLICE_X4Y125_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y125_SLICE_X4Y125_BO5),
.O6(CLBLL_L_X4Y125_SLICE_X4Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0cfc0c0cfc0)
  ) CLBLL_L_X4Y125_SLICE_X4Y125_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y122_SLICE_X3Y122_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y121_SLICE_X10Y121_AO5),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X8Y124_SLICE_X11Y124_BQ),
.O5(CLBLL_L_X4Y125_SLICE_X4Y125_AO5),
.O6(CLBLL_L_X4Y125_SLICE_X4Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y125_SLICE_X5Y125_AO6),
.Q(CLBLL_L_X4Y125_SLICE_X5Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y125_SLICE_X5Y125_BO6),
.Q(CLBLL_L_X4Y125_SLICE_X5Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h73507350ffff7350)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_DLUT (
.I0(CLBLL_L_X4Y126_SLICE_X4Y126_CO5),
.I1(CLBLL_L_X2Y129_SLICE_X0Y129_AO6),
.I2(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.I3(CLBLM_R_X5Y122_SLICE_X6Y122_AQ),
.I4(CLBLM_R_X7Y125_SLICE_X9Y125_DQ),
.I5(CLBLL_L_X4Y126_SLICE_X4Y126_BO6),
.O5(CLBLL_L_X4Y125_SLICE_X5Y125_DO5),
.O6(CLBLL_L_X4Y125_SLICE_X5Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f00afaacfccefee)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_CLUT (
.I0(CLBLM_R_X5Y125_SLICE_X7Y125_AQ),
.I1(CLBLL_L_X4Y124_SLICE_X5Y124_BQ),
.I2(CLBLL_L_X2Y129_SLICE_X0Y129_AO6),
.I3(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.I4(CLBLM_R_X3Y130_SLICE_X3Y130_AO6),
.I5(CLBLL_L_X4Y126_SLICE_X4Y126_BO6),
.O5(CLBLL_L_X4Y125_SLICE_X5Y125_CO5),
.O6(CLBLL_L_X4Y125_SLICE_X5Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aafff0f088cc)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_BLUT (
.I0(CLBLM_R_X11Y120_SLICE_X14Y120_DO6),
.I1(CLBLL_L_X4Y125_SLICE_X5Y125_BQ),
.I2(CLBLL_L_X4Y124_SLICE_X5Y124_BQ),
.I3(CLBLM_R_X7Y123_SLICE_X9Y123_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y123_SLICE_X7Y123_BQ),
.O5(CLBLL_L_X4Y125_SLICE_X5Y125_BO5),
.O6(CLBLL_L_X4Y125_SLICE_X5Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33cc00fd31ec20)
  ) CLBLL_L_X4Y125_SLICE_X5Y125_ALUT (
.I0(CLBLM_R_X7Y123_SLICE_X9Y123_A5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y125_SLICE_X5Y125_AQ),
.I3(CLBLM_R_X5Y128_SLICE_X6Y128_A5Q),
.I4(CLBLL_L_X4Y120_SLICE_X5Y120_AQ),
.I5(CLBLM_R_X11Y120_SLICE_X14Y120_DO6),
.O5(CLBLL_L_X4Y125_SLICE_X5Y125_AO5),
.O6(CLBLL_L_X4Y125_SLICE_X5Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y126_SLICE_X4Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y126_SLICE_X4Y126_AO6),
.Q(CLBLL_L_X4Y126_SLICE_X4Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLL_L_X4Y126_SLICE_X4Y126_DLUT (
.I0(CLBLL_L_X2Y129_SLICE_X1Y129_CO6),
.I1(CLBLL_L_X2Y126_SLICE_X0Y126_BO6),
.I2(CLBLL_L_X4Y129_SLICE_X5Y129_DO6),
.I3(CLBLL_L_X4Y126_SLICE_X5Y126_DO6),
.I4(CLBLM_R_X3Y128_SLICE_X2Y128_DO6),
.I5(CLBLL_L_X4Y125_SLICE_X5Y125_DO6),
.O5(CLBLL_L_X4Y126_SLICE_X4Y126_DO5),
.O6(CLBLL_L_X4Y126_SLICE_X4Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefffefffeffffff)
  ) CLBLL_L_X4Y126_SLICE_X4Y126_CLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y126_SLICE_X4Y126_CO5),
.O6(CLBLL_L_X4Y126_SLICE_X4Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffdffffffeff)
  ) CLBLL_L_X4Y126_SLICE_X4Y126_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y126_SLICE_X4Y126_BO5),
.O6(CLBLL_L_X4Y126_SLICE_X4Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf088f000f000f000)
  ) CLBLL_L_X4Y126_SLICE_X4Y126_ALUT (
.I0(CLBLM_R_X5Y128_SLICE_X6Y128_DQ),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_A5Q),
.I2(CLBLM_R_X7Y122_SLICE_X9Y122_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y129_SLICE_X5Y129_AQ),
.I5(CLBLL_L_X4Y119_SLICE_X4Y119_DQ),
.O5(CLBLL_L_X4Y126_SLICE_X4Y126_AO5),
.O6(CLBLL_L_X4Y126_SLICE_X4Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f000f0aafaaafa)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_DLUT (
.I0(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y128_SLICE_X10Y128_CQ),
.I3(CLBLL_L_X4Y126_SLICE_X4Y126_BO5),
.I4(1'b1),
.I5(CLBLM_R_X3Y130_SLICE_X3Y130_AO6),
.O5(CLBLL_L_X4Y126_SLICE_X5Y126_DO5),
.O6(CLBLL_L_X4Y126_SLICE_X5Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000fa0accccfece)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_CLUT (
.I0(CLBLM_R_X5Y128_SLICE_X6Y128_AQ),
.I1(CLBLM_R_X5Y120_SLICE_X7Y120_BQ),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_B5Q),
.I4(CLBLL_L_X4Y126_SLICE_X4Y126_CO6),
.I5(CLBLM_R_X3Y130_SLICE_X3Y130_AO6),
.O5(CLBLL_L_X4Y126_SLICE_X5Y126_CO5),
.O6(CLBLL_L_X4Y126_SLICE_X5Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h73735050ff73ff50)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_BLUT (
.I0(CLBLL_L_X2Y129_SLICE_X0Y129_AO6),
.I1(CLBLL_L_X4Y126_SLICE_X4Y126_BO6),
.I2(CLBLL_L_X4Y124_SLICE_X5Y124_AQ),
.I3(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.I4(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.I5(CLBLL_L_X4Y126_SLICE_X4Y126_BO5),
.O5(CLBLL_L_X4Y126_SLICE_X5Y126_BO5),
.O6(CLBLL_L_X4Y126_SLICE_X5Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7755735033007350)
  ) CLBLL_L_X4Y126_SLICE_X5Y126_ALUT (
.I0(CLBLL_L_X4Y126_SLICE_X4Y126_CO6),
.I1(CLBLM_R_X3Y130_SLICE_X3Y130_AO6),
.I2(CLBLM_L_X10Y125_SLICE_X13Y125_AQ),
.I3(CLBLL_L_X4Y121_SLICE_X5Y121_BQ),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_L_X8Y126_SLICE_X11Y126_AQ),
.O5(CLBLL_L_X4Y126_SLICE_X5Y126_AO5),
.O6(CLBLL_L_X4Y126_SLICE_X5Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h020f020f02020202)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_DLUT (
.I0(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.I1(CLBLL_L_X2Y130_SLICE_X0Y130_BO6),
.I2(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.I3(CLBLL_L_X2Y130_SLICE_X0Y130_AO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.O5(CLBLL_L_X4Y127_SLICE_X4Y127_DO5),
.O6(CLBLL_L_X4Y127_SLICE_X4Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000a000a333b000a)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_CLUT (
.I0(CLBLM_R_X3Y122_SLICE_X2Y122_DQ),
.I1(CLBLL_L_X2Y130_SLICE_X0Y130_BO6),
.I2(CLBLL_L_X2Y130_SLICE_X0Y130_CO5),
.I3(CLBLL_L_X2Y128_SLICE_X1Y128_AO6),
.I4(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.I5(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.O5(CLBLL_L_X4Y127_SLICE_X4Y127_CO5),
.O6(CLBLL_L_X4Y127_SLICE_X4Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffbaba30ba)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_BLUT (
.I0(CLBLM_R_X7Y126_SLICE_X9Y126_C5Q),
.I1(CLBLL_L_X2Y126_SLICE_X0Y126_AO6),
.I2(CLBLM_R_X5Y126_SLICE_X7Y126_BQ),
.I3(RIOB33_X105Y137_IOB_X1Y137_I),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(CLBLM_R_X3Y127_SLICE_X3Y127_DO6),
.O5(CLBLL_L_X4Y127_SLICE_X4Y127_BO5),
.O6(CLBLL_L_X4Y127_SLICE_X4Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00550c5d00000c0c)
  ) CLBLL_L_X4Y127_SLICE_X4Y127_ALUT (
.I0(CLBLL_L_X2Y128_SLICE_X1Y128_AO5),
.I1(CLBLM_R_X3Y121_SLICE_X2Y121_AQ),
.I2(CLBLL_L_X2Y130_SLICE_X0Y130_CO5),
.I3(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.I4(CLBLL_L_X2Y130_SLICE_X0Y130_AO6),
.I5(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.O5(CLBLL_L_X4Y127_SLICE_X4Y127_AO5),
.O6(CLBLL_L_X4Y127_SLICE_X4Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000022ff2222)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_DLUT (
.I0(CLBLL_L_X4Y122_SLICE_X5Y122_AQ),
.I1(CLBLL_L_X2Y128_SLICE_X1Y128_AO6),
.I2(1'b1),
.I3(CLBLL_L_X2Y130_SLICE_X0Y130_BO6),
.I4(CLBLM_R_X5Y125_SLICE_X7Y125_BQ),
.I5(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.O5(CLBLL_L_X4Y127_SLICE_X5Y127_DO5),
.O6(CLBLL_L_X4Y127_SLICE_X5Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1111000051515050)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_CLUT (
.I0(CLBLL_L_X2Y130_SLICE_X0Y130_CO5),
.I1(CLBLL_L_X2Y130_SLICE_X0Y130_AO6),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(1'b1),
.I4(CLBLM_R_X3Y121_SLICE_X2Y121_C5Q),
.I5(CLBLL_L_X2Y130_SLICE_X0Y130_BO6),
.O5(CLBLL_L_X4Y127_SLICE_X5Y127_CO5),
.O6(CLBLL_L_X4Y127_SLICE_X5Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0303000003000300)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.I2(CLBLL_L_X2Y130_SLICE_X1Y130_AO6),
.I3(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I4(CLBLL_L_X4Y124_SLICE_X5Y124_CQ),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLL_L_X4Y127_SLICE_X5Y127_BO5),
.O6(CLBLL_L_X4Y127_SLICE_X5Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffafffffffe)
  ) CLBLL_L_X4Y127_SLICE_X5Y127_ALUT (
.I0(CLBLM_R_X5Y127_SLICE_X7Y127_DO6),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_CQ),
.I2(CLBLL_L_X4Y127_SLICE_X4Y127_CO6),
.I3(CLBLL_L_X4Y127_SLICE_X5Y127_BO6),
.I4(CLBLL_L_X4Y127_SLICE_X5Y127_CO6),
.I5(CLBLL_L_X2Y128_SLICE_X0Y128_AO5),
.O5(CLBLL_L_X4Y127_SLICE_X5Y127_AO5),
.O6(CLBLL_L_X4Y127_SLICE_X5Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55005500f5f0f5f0)
  ) CLBLL_L_X4Y128_SLICE_X4Y128_DLUT (
.I0(CLBLL_L_X4Y126_SLICE_X4Y126_CO5),
.I1(1'b1),
.I2(CLBLL_L_X4Y119_SLICE_X5Y119_CQ),
.I3(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y130_SLICE_X3Y130_AO6),
.O5(CLBLL_L_X4Y128_SLICE_X4Y128_DO5),
.O6(CLBLL_L_X4Y128_SLICE_X4Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1033101010331010)
  ) CLBLL_L_X4Y128_SLICE_X4Y128_CLUT (
.I0(CLBLL_L_X2Y128_SLICE_X1Y128_AO6),
.I1(CLBLL_L_X2Y130_SLICE_X0Y130_CO5),
.I2(CLBLM_R_X7Y123_SLICE_X9Y123_BQ),
.I3(CLBLL_L_X2Y130_SLICE_X0Y130_BO6),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y128_SLICE_X4Y128_CO5),
.O6(CLBLL_L_X4Y128_SLICE_X4Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffefffefe)
  ) CLBLL_L_X4Y128_SLICE_X4Y128_BLUT (
.I0(CLBLM_R_X5Y128_SLICE_X7Y128_CO6),
.I1(CLBLL_L_X4Y128_SLICE_X5Y128_DO6),
.I2(CLBLL_L_X4Y127_SLICE_X4Y127_AO6),
.I3(CLBLM_R_X3Y130_SLICE_X2Y130_BO6),
.I4(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.I5(CLBLL_L_X4Y128_SLICE_X4Y128_CO6),
.O5(CLBLL_L_X4Y128_SLICE_X4Y128_BO5),
.O6(CLBLL_L_X4Y128_SLICE_X4Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLL_L_X4Y128_SLICE_X4Y128_ALUT (
.I0(CLBLL_L_X4Y128_SLICE_X4Y128_DO6),
.I1(CLBLL_L_X4Y126_SLICE_X5Y126_BO6),
.I2(CLBLL_L_X2Y129_SLICE_X1Y129_CO6),
.I3(CLBLL_L_X4Y128_SLICE_X4Y128_BO6),
.I4(CLBLL_L_X4Y127_SLICE_X4Y127_BO6),
.I5(CLBLM_R_X3Y128_SLICE_X3Y128_DO6),
.O5(CLBLL_L_X4Y128_SLICE_X4Y128_AO5),
.O6(CLBLL_L_X4Y128_SLICE_X4Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000100000)
  ) CLBLL_L_X4Y128_SLICE_X5Y128_DLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_L_X10Y129_SLICE_X13Y129_AQ),
.I5(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.O5(CLBLL_L_X4Y128_SLICE_X5Y128_DO5),
.O6(CLBLL_L_X4Y128_SLICE_X5Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffba)
  ) CLBLL_L_X4Y128_SLICE_X5Y128_CLUT (
.I0(CLBLL_L_X4Y128_SLICE_X5Y128_AO6),
.I1(CLBLL_L_X2Y128_SLICE_X0Y128_AO5),
.I2(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I3(CLBLM_R_X5Y127_SLICE_X6Y127_DO6),
.I4(CLBLM_R_X3Y128_SLICE_X3Y128_AO6),
.I5(CLBLL_L_X4Y128_SLICE_X5Y128_BO6),
.O5(CLBLL_L_X4Y128_SLICE_X5Y128_CO5),
.O6(CLBLL_L_X4Y128_SLICE_X5Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f0022222f22)
  ) CLBLL_L_X4Y128_SLICE_X5Y128_BLUT (
.I0(CLBLM_R_X5Y123_SLICE_X7Y123_AQ),
.I1(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.I2(CLBLL_L_X2Y128_SLICE_X1Y128_AO6),
.I3(CLBLL_L_X4Y125_SLICE_X5Y125_AQ),
.I4(CLBLL_L_X2Y130_SLICE_X0Y130_CO5),
.I5(CLBLL_L_X2Y128_SLICE_X1Y128_AO5),
.O5(CLBLL_L_X4Y128_SLICE_X5Y128_BO5),
.O6(CLBLL_L_X4Y128_SLICE_X5Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000222200f022f2)
  ) CLBLL_L_X4Y128_SLICE_X5Y128_ALUT (
.I0(CLBLM_R_X7Y126_SLICE_X8Y126_CQ),
.I1(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(CLBLL_L_X2Y130_SLICE_X0Y130_CO5),
.I4(CLBLL_L_X2Y130_SLICE_X0Y130_AO6),
.I5(CLBLL_L_X2Y130_SLICE_X0Y130_BO6),
.O5(CLBLL_L_X4Y128_SLICE_X5Y128_AO5),
.O6(CLBLL_L_X4Y128_SLICE_X5Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y129_SLICE_X4Y129_AO6),
.Q(CLBLL_L_X4Y129_SLICE_X4Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fff0fcfcfffc)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_DLUT (
.I0(1'b1),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(CLBLL_L_X4Y127_SLICE_X4Y127_DO6),
.I3(CLBLL_L_X4Y120_SLICE_X5Y120_CQ),
.I4(CLBLL_L_X4Y129_SLICE_X4Y129_BO5),
.I5(CLBLM_R_X3Y129_SLICE_X3Y129_AO6),
.O5(CLBLL_L_X4Y129_SLICE_X4Y129_DO5),
.O6(CLBLL_L_X4Y129_SLICE_X4Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0003000100020000)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_CLUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(CLBLL_L_X4Y130_SLICE_X4Y130_AO5),
.I2(RIOB33_X105Y135_IOB_X1Y135_I),
.I3(CLBLL_L_X2Y130_SLICE_X0Y130_BO6),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(CLBLL_L_X4Y122_SLICE_X4Y122_AQ),
.O5(CLBLL_L_X4Y129_SLICE_X4Y129_CO5),
.O6(CLBLL_L_X4Y129_SLICE_X4Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffffffbffff)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_BLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLL_L_X2Y130_SLICE_X0Y130_CO5),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y129_SLICE_X4Y129_BO5),
.O6(CLBLL_L_X4Y129_SLICE_X4Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000fffc00fc)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y125_SLICE_X6Y125_A5Q),
.I2(CLBLL_L_X4Y129_SLICE_X4Y129_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y125_SLICE_X4Y125_AQ),
.I5(CLBLL_L_X2Y119_SLICE_X1Y119_BO6),
.O5(CLBLL_L_X4Y129_SLICE_X4Y129_AO5),
.O6(CLBLL_L_X4Y129_SLICE_X4Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y129_SLICE_X5Y129_AO6),
.Q(CLBLL_L_X4Y129_SLICE_X5Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffdc)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_DLUT (
.I0(CLBLL_L_X4Y129_SLICE_X4Y129_BO6),
.I1(CLBLL_L_X4Y129_SLICE_X4Y129_CO6),
.I2(CLBLM_R_X7Y125_SLICE_X8Y125_DQ),
.I3(CLBLL_L_X4Y129_SLICE_X5Y129_CO6),
.I4(CLBLM_R_X5Y128_SLICE_X7Y128_DO6),
.I5(CLBLL_L_X4Y129_SLICE_X5Y129_BO6),
.O5(CLBLL_L_X4Y129_SLICE_X5Y129_DO5),
.O6(CLBLL_L_X4Y129_SLICE_X5Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0537050500330000)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_CLUT (
.I0(CLBLL_L_X2Y130_SLICE_X0Y130_AO6),
.I1(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.I2(CLBLL_L_X2Y130_SLICE_X0Y130_CO5),
.I3(CLBLL_L_X2Y128_SLICE_X1Y128_AO5),
.I4(CLBLM_R_X7Y128_SLICE_X8Y128_DQ),
.I5(CLBLM_R_X3Y121_SLICE_X2Y121_BQ),
.O5(CLBLL_L_X4Y129_SLICE_X5Y129_CO5),
.O6(CLBLL_L_X4Y129_SLICE_X5Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010000000000)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(CLBLM_L_X10Y125_SLICE_X13Y125_BQ),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(RIOB33_X105Y133_IOB_X1Y133_I),
.O5(CLBLL_L_X4Y129_SLICE_X5Y129_BO5),
.O6(CLBLL_L_X4Y129_SLICE_X5Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00fcf0cc00fcf0)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y129_SLICE_X8Y129_A5Q),
.I2(CLBLL_L_X4Y129_SLICE_X5Y129_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X2Y120_SLICE_X1Y120_BO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y129_SLICE_X5Y129_AO5),
.O6(CLBLL_L_X4Y129_SLICE_X5Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8c8c8c8c8c8cff8c)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_DLUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(CLBLL_L_X4Y125_SLICE_X4Y125_C5Q),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(CLBLM_R_X5Y129_SLICE_X6Y129_CQ),
.I4(CLBLL_L_X2Y130_SLICE_X0Y130_AO6),
.I5(CLBLL_L_X2Y130_SLICE_X0Y130_CO6),
.O5(CLBLL_L_X4Y130_SLICE_X4Y130_DO5),
.O6(CLBLL_L_X4Y130_SLICE_X4Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffdc)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_CLUT (
.I0(CLBLM_R_X3Y130_SLICE_X3Y130_AO6),
.I1(CLBLL_L_X4Y130_SLICE_X5Y130_AO6),
.I2(CLBLM_R_X3Y123_SLICE_X2Y123_AQ),
.I3(CLBLL_L_X4Y131_SLICE_X4Y131_AO6),
.I4(CLBLL_L_X4Y127_SLICE_X4Y127_DO6),
.I5(CLBLL_L_X4Y130_SLICE_X4Y130_BO6),
.O5(CLBLL_L_X4Y130_SLICE_X4Y130_CO5),
.O6(CLBLL_L_X4Y130_SLICE_X4Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0545ffff0044)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_BLUT (
.I0(CLBLL_L_X2Y130_SLICE_X0Y130_CO6),
.I1(LIOB33_X0Y67_IOB_X0Y68_I),
.I2(CLBLL_L_X2Y130_SLICE_X0Y130_AO6),
.I3(CLBLL_L_X2Y130_SLICE_X0Y130_BO6),
.I4(CLBLL_L_X4Y130_SLICE_X4Y130_AO6),
.I5(CLBLM_R_X5Y129_SLICE_X6Y129_CQ),
.O5(CLBLL_L_X4Y130_SLICE_X4Y130_BO5),
.O6(CLBLL_L_X4Y130_SLICE_X4Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc4444ffffff55)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_ALUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(CLBLL_L_X4Y125_SLICE_X4Y125_C5Q),
.I2(1'b1),
.I3(RIOB33_X105Y129_IOB_X1Y130_I),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y130_SLICE_X4Y130_AO5),
.O6(CLBLL_L_X4Y130_SLICE_X4Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y130_SLICE_X5Y130_DO5),
.O6(CLBLL_L_X4Y130_SLICE_X5Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y130_SLICE_X5Y130_CO5),
.O6(CLBLL_L_X4Y130_SLICE_X5Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y130_SLICE_X5Y130_BO5),
.O6(CLBLL_L_X4Y130_SLICE_X5Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h003f000f00330000)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y130_SLICE_X0Y130_BO6),
.I2(CLBLL_L_X2Y130_SLICE_X0Y130_AO6),
.I3(CLBLL_L_X2Y130_SLICE_X0Y130_CO5),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(CLBLL_L_X4Y120_SLICE_X5Y120_CQ),
.O5(CLBLL_L_X4Y130_SLICE_X5Y130_AO5),
.O6(CLBLL_L_X4Y130_SLICE_X5Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X4Y131_DO5),
.O6(CLBLL_L_X4Y131_SLICE_X4Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X4Y131_CO5),
.O6(CLBLL_L_X4Y131_SLICE_X4Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffefeffffffff)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_BLUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(RIOB33_X105Y135_IOB_X1Y136_I),
.I2(RIOB33_X105Y129_IOB_X1Y130_I),
.I3(1'b1),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(RIOB33_X105Y137_IOB_X1Y137_I),
.O5(CLBLL_L_X4Y131_SLICE_X4Y131_BO5),
.O6(CLBLL_L_X4Y131_SLICE_X4Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000800000000)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(CLBLM_R_X7Y129_SLICE_X8Y129_DQ),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLL_L_X4Y131_SLICE_X4Y131_AO5),
.O6(CLBLL_L_X4Y131_SLICE_X4Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X5Y131_DO5),
.O6(CLBLL_L_X4Y131_SLICE_X5Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X5Y131_CO5),
.O6(CLBLL_L_X4Y131_SLICE_X5Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X5Y131_BO5),
.O6(CLBLL_L_X4Y131_SLICE_X5Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X5Y131_AO5),
.O6(CLBLL_L_X4Y131_SLICE_X5Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y124_SLICE_X54Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y124_SLICE_X54Y124_DO5),
.O6(CLBLL_L_X36Y124_SLICE_X54Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y124_SLICE_X54Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y124_SLICE_X54Y124_CO5),
.O6(CLBLL_L_X36Y124_SLICE_X54Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y124_SLICE_X54Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y124_SLICE_X54Y124_BO5),
.O6(CLBLL_L_X36Y124_SLICE_X54Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0030003000300030)
  ) CLBLL_L_X36Y124_SLICE_X54Y124_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y123_SLICE_X6Y123_BQ),
.I2(RIOB33_X105Y119_IOB_X1Y119_I),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y124_SLICE_X54Y124_AO5),
.O6(CLBLL_L_X36Y124_SLICE_X54Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y124_SLICE_X55Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y124_SLICE_X55Y124_DO5),
.O6(CLBLL_L_X36Y124_SLICE_X55Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y124_SLICE_X55Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y124_SLICE_X55Y124_CO5),
.O6(CLBLL_L_X36Y124_SLICE_X55Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y124_SLICE_X55Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y124_SLICE_X55Y124_BO5),
.O6(CLBLL_L_X36Y124_SLICE_X55Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y124_SLICE_X55Y124_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y124_SLICE_X55Y124_AO5),
.O6(CLBLL_L_X36Y124_SLICE_X55Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_DO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_CO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_BO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y123_IOB_X1Y124_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_AO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_DO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_CO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_BO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_AO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y116_SLICE_X10Y116_BO6),
.Q(CLBLM_L_X8Y116_SLICE_X10Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5c5c55555c5c5c5c)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_DLUT (
.I0(CLBLL_L_X4Y120_SLICE_X4Y120_C5Q),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_BO6),
.I2(CLBLM_R_X3Y124_SLICE_X3Y124_DO6),
.I3(1'b1),
.I4(CLBLM_R_X7Y118_SLICE_X9Y118_BO5),
.I5(CLBLM_R_X5Y118_SLICE_X7Y118_BO5),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_DO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3335ccc5333accca)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_CLUT (
.I0(CLBLM_L_X8Y116_SLICE_X10Y116_AO6),
.I1(CLBLM_L_X8Y123_SLICE_X10Y123_CQ),
.I2(CLBLM_R_X3Y124_SLICE_X3Y124_DO6),
.I3(CLBLM_R_X3Y126_SLICE_X2Y126_BO6),
.I4(CLBLM_R_X7Y124_SLICE_X8Y124_B5Q),
.I5(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_CO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaf0aac0aac0)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_BLUT (
.I0(CLBLM_R_X3Y123_SLICE_X2Y123_DQ),
.I1(CLBLM_L_X8Y116_SLICE_X10Y116_BQ),
.I2(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X5Y116_SLICE_X7Y116_BQ),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_BO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0004fffbfbfbfbfb)
  ) CLBLM_L_X8Y116_SLICE_X10Y116_ALUT (
.I0(CLBLL_L_X4Y117_SLICE_X5Y117_BQ),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_CQ),
.I2(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I3(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_DQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y116_SLICE_X10Y116_AO5),
.O6(CLBLM_L_X8Y116_SLICE_X10Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_DO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555f7045555f704)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_CLUT (
.I0(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.I1(CLBLM_R_X5Y118_SLICE_X7Y118_BO5),
.I2(CLBLM_R_X7Y118_SLICE_X9Y118_BO5),
.I3(CLBLM_R_X7Y115_SLICE_X9Y115_AO6),
.I4(CLBLM_R_X3Y124_SLICE_X3Y124_DO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_CO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0bff00f400f40bff)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_BLUT (
.I0(CLBLM_R_X7Y118_SLICE_X9Y118_BO5),
.I1(CLBLM_R_X5Y118_SLICE_X7Y118_BO5),
.I2(CLBLM_R_X3Y124_SLICE_X3Y124_DO6),
.I3(CLBLM_R_X7Y118_SLICE_X8Y118_C5Q),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_CQ),
.I5(CLBLM_L_X8Y118_SLICE_X11Y118_CO6),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_BO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X8Y116_SLICE_X11Y116_ALUT (
.I0(CLBLM_L_X8Y117_SLICE_X11Y117_BO6),
.I1(CLBLM_R_X7Y116_SLICE_X9Y116_CO6),
.I2(CLBLM_L_X8Y116_SLICE_X10Y116_CO6),
.I3(CLBLM_L_X8Y116_SLICE_X11Y116_BO6),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_DO6),
.I5(CLBLM_L_X8Y116_SLICE_X11Y116_CO6),
.O5(CLBLM_L_X8Y116_SLICE_X11Y116_AO5),
.O6(CLBLM_L_X8Y116_SLICE_X11Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y117_SLICE_X10Y117_AO6),
.Q(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y117_SLICE_X10Y117_BO6),
.Q(CLBLM_L_X8Y117_SLICE_X10Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000cccc00ff40bf)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_DLUT (
.I0(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I1(CLBLL_L_X4Y117_SLICE_X5Y117_BQ),
.I2(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I3(CLBLM_L_X10Y119_SLICE_X12Y119_DQ),
.I4(CLBLM_R_X5Y116_SLICE_X7Y116_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y117_SLICE_X10Y117_DO5),
.O6(CLBLM_L_X8Y117_SLICE_X10Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd555ffff8000ffff)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_CLUT (
.I0(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I1(CLBLL_L_X4Y117_SLICE_X5Y117_BQ),
.I2(CLBLM_R_X5Y116_SLICE_X7Y116_CQ),
.I3(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I4(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y117_SLICE_X10Y117_CO5),
.O6(CLBLM_L_X8Y117_SLICE_X10Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffe0ffe000e000e0)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_BLUT (
.I0(CLBLM_R_X7Y118_SLICE_X8Y118_DQ),
.I1(CLBLM_L_X8Y117_SLICE_X10Y117_BQ),
.I2(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y117_SLICE_X5Y117_AQ),
.O5(CLBLM_L_X8Y117_SLICE_X10Y117_BO5),
.O6(CLBLM_L_X8Y117_SLICE_X10Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffeccdc33320010)
  ) CLBLM_L_X8Y117_SLICE_X10Y117_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I4(CLBLM_R_X5Y117_SLICE_X6Y117_BQ),
.I5(CLBLM_L_X8Y116_SLICE_X10Y116_BQ),
.O5(CLBLM_L_X8Y117_SLICE_X10Y117_AO5),
.O6(CLBLM_L_X8Y117_SLICE_X10Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777bbbbddddeeee)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_DLUT (
.I0(CLBLL_L_X4Y120_SLICE_X4Y120_C5Q),
.I1(CLBLM_R_X7Y118_SLICE_X9Y118_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X8Y116_SLICE_X10Y116_BQ),
.I5(CLBLM_L_X10Y124_SLICE_X13Y124_D5Q),
.O5(CLBLM_L_X8Y117_SLICE_X11Y117_DO5),
.O6(CLBLM_L_X8Y117_SLICE_X11Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff7bdeffff7bde)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_CLUT (
.I0(CLBLM_L_X8Y118_SLICE_X11Y118_AQ),
.I1(CLBLM_L_X8Y119_SLICE_X11Y119_CQ),
.I2(CLBLM_R_X7Y118_SLICE_X8Y118_C5Q),
.I3(CLBLM_L_X8Y123_SLICE_X10Y123_CQ),
.I4(CLBLM_L_X8Y117_SLICE_X11Y117_DO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y117_SLICE_X11Y117_CO5),
.O6(CLBLM_L_X8Y117_SLICE_X11Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff01bb10ff04ee4)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_BLUT (
.I0(CLBLM_R_X3Y124_SLICE_X3Y124_DO6),
.I1(CLBLM_L_X8Y117_SLICE_X10Y117_DO5),
.I2(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.I3(CLBLM_L_X10Y124_SLICE_X13Y124_D5Q),
.I4(CLBLM_R_X3Y126_SLICE_X2Y126_BO6),
.I5(CLBLM_L_X8Y117_SLICE_X11Y117_AO5),
.O5(CLBLM_L_X8Y117_SLICE_X11Y117_BO5),
.O6(CLBLM_L_X8Y117_SLICE_X11Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff3f300ff20df)
  ) CLBLM_L_X8Y117_SLICE_X11Y117_ALUT (
.I0(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I1(CLBLL_L_X4Y117_SLICE_X5Y117_BQ),
.I2(CLBLM_R_X5Y116_SLICE_X7Y116_CQ),
.I3(CLBLM_L_X8Y117_SLICE_X10Y117_BQ),
.I4(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y117_SLICE_X11Y117_AO5),
.O6(CLBLM_L_X8Y117_SLICE_X11Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y118_SLICE_X10Y118_AO6),
.Q(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y118_SLICE_X10Y118_BO6),
.Q(CLBLM_L_X8Y118_SLICE_X10Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y118_SLICE_X10Y118_CO6),
.Q(CLBLM_L_X8Y118_SLICE_X10Y118_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333111133333131)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_DLUT (
.I0(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.I1(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(1'b1),
.I4(CLBLM_R_X3Y123_SLICE_X2Y123_DQ),
.I5(CLBLM_R_X3Y126_SLICE_X3Y126_AO6),
.O5(CLBLM_L_X8Y118_SLICE_X10Y118_DO5),
.O6(CLBLM_L_X8Y118_SLICE_X10Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaacc00cccc)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_CLUT (
.I0(CLBLM_L_X8Y118_SLICE_X10Y118_BQ),
.I1(CLBLM_L_X8Y118_SLICE_X10Y118_CQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y118_SLICE_X10Y118_CO5),
.O6(CLBLM_L_X8Y118_SLICE_X10Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ccacccac)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_BLUT (
.I0(CLBLM_R_X7Y118_SLICE_X9Y118_CO6),
.I1(CLBLM_L_X8Y118_SLICE_X10Y118_BQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I4(CLBLM_L_X8Y118_SLICE_X11Y118_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y118_SLICE_X10Y118_BO5),
.O6(CLBLM_L_X8Y118_SLICE_X10Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc05cc0000ff00f0)
  ) CLBLM_L_X8Y118_SLICE_X10Y118_ALUT (
.I0(CLBLM_L_X8Y118_SLICE_X10Y118_DO6),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_AQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y118_SLICE_X10Y118_AO5),
.O6(CLBLM_L_X8Y118_SLICE_X10Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y118_SLICE_X11Y118_AO6),
.Q(CLBLM_L_X8Y118_SLICE_X11Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y118_SLICE_X11Y118_BO6),
.Q(CLBLM_L_X8Y118_SLICE_X11Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_DLUT (
.I0(CLBLM_R_X7Y118_SLICE_X9Y118_AQ),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_BQ),
.I2(CLBLM_R_X7Y118_SLICE_X8Y118_AQ),
.I3(CLBLM_L_X8Y119_SLICE_X11Y119_CQ),
.I4(CLBLM_L_X8Y118_SLICE_X11Y118_AQ),
.I5(CLBLM_L_X8Y116_SLICE_X10Y116_BQ),
.O5(CLBLM_L_X8Y118_SLICE_X11Y118_DO5),
.O6(CLBLM_L_X8Y118_SLICE_X11Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00008800f0f0f0d2)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_CLUT (
.I0(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I1(CLBLL_L_X4Y117_SLICE_X5Y117_BQ),
.I2(CLBLM_L_X10Y119_SLICE_X13Y119_DO6),
.I3(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I4(CLBLM_R_X5Y116_SLICE_X7Y116_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y118_SLICE_X11Y118_CO5),
.O6(CLBLM_L_X8Y118_SLICE_X11Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0ffc000f000c0)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y118_SLICE_X11Y118_BQ),
.I2(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y118_SLICE_X7Y118_AQ),
.I5(CLBLM_L_X8Y119_SLICE_X11Y119_CQ),
.O5(CLBLM_L_X8Y118_SLICE_X11Y118_BO5),
.O6(CLBLM_L_X8Y118_SLICE_X11Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcff0000fc0000)
  ) CLBLM_L_X8Y118_SLICE_X11Y118_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y118_SLICE_X9Y118_AQ),
.I2(CLBLM_L_X8Y118_SLICE_X11Y118_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I5(CLBLM_R_X11Y120_SLICE_X14Y120_AQ),
.O5(CLBLM_L_X8Y118_SLICE_X11Y118_AO5),
.O6(CLBLM_L_X8Y118_SLICE_X11Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y119_SLICE_X10Y119_AO6),
.Q(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y119_SLICE_X10Y119_BO6),
.Q(CLBLM_L_X8Y119_SLICE_X10Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_DLUT (
.I0(CLBLM_R_X5Y116_SLICE_X6Y116_AQ),
.I1(CLBLM_L_X10Y119_SLICE_X12Y119_CQ),
.I2(CLBLM_R_X7Y119_SLICE_X8Y119_CQ),
.I3(CLBLM_L_X10Y119_SLICE_X12Y119_DQ),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_DQ),
.I5(CLBLM_L_X8Y119_SLICE_X11Y119_BQ),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_DO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000556600000f0f)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_CLUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_DQ),
.I1(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I2(CLBLM_L_X8Y123_SLICE_X10Y123_CQ),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_AO5),
.I4(CLBLM_L_X8Y125_SLICE_X10Y125_DQ),
.I5(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_CO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf088f088f088f088)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y119_SLICE_X10Y119_BQ),
.I2(CLBLM_R_X3Y120_SLICE_X2Y120_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_BO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf555cccca000)
  ) CLBLM_L_X8Y119_SLICE_X10Y119_ALUT (
.I0(CLBLM_L_X8Y123_SLICE_X10Y123_DO6),
.I1(CLBLM_R_X5Y117_SLICE_X6Y117_CQ),
.I2(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y120_SLICE_X12Y120_CQ),
.O5(CLBLM_L_X8Y119_SLICE_X10Y119_AO5),
.O6(CLBLM_L_X8Y119_SLICE_X10Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y119_SLICE_X11Y119_AO6),
.Q(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y119_SLICE_X11Y119_BO6),
.Q(CLBLM_L_X8Y119_SLICE_X11Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y119_SLICE_X11Y119_CO6),
.Q(CLBLM_L_X8Y119_SLICE_X11Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000003a30000f353)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_DLUT (
.I0(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I1(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.I2(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I3(CLBLM_L_X8Y116_SLICE_X10Y116_AO5),
.I4(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.I5(CLBLM_L_X8Y117_SLICE_X10Y117_BQ),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_DO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0eef0eef000f000)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_CLUT (
.I0(CLBLM_L_X8Y118_SLICE_X11Y118_AQ),
.I1(CLBLM_L_X8Y119_SLICE_X11Y119_CQ),
.I2(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_CO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500eeaa4400)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y119_SLICE_X11Y119_BQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I4(CLBLL_L_X4Y122_SLICE_X4Y122_A5Q),
.I5(CLBLM_L_X10Y119_SLICE_X13Y119_DO6),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_BO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc55550505)
  ) CLBLM_L_X8Y119_SLICE_X11Y119_ALUT (
.I0(CLBLM_L_X8Y119_SLICE_X11Y119_DO6),
.I1(CLBLM_R_X11Y120_SLICE_X14Y120_BQ),
.I2(RIOB33_X105Y141_IOB_X1Y142_I),
.I3(1'b1),
.I4(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y119_SLICE_X11Y119_AO5),
.O6(CLBLM_L_X8Y119_SLICE_X11Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X10Y120_AO6),
.Q(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y120_SLICE_X10Y120_BO6),
.Q(CLBLM_L_X8Y120_SLICE_X10Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5ff55ff5affaaffa)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_DLUT (
.I0(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y120_SLICE_X8Y120_CQ),
.I3(CLBLM_L_X12Y121_SLICE_X16Y121_AQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y120_SLICE_X12Y120_CQ),
.O5(CLBLM_L_X8Y120_SLICE_X10Y120_DO5),
.O6(CLBLM_L_X8Y120_SLICE_X10Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996666999966)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_CLUT (
.I0(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I1(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y119_SLICE_X7Y119_BQ),
.I4(CLBLM_R_X7Y120_SLICE_X8Y120_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y120_SLICE_X10Y120_CO5),
.O6(CLBLM_L_X8Y120_SLICE_X10Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ccaacc00ccaa)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_BLUT (
.I0(CLBLM_L_X10Y122_SLICE_X13Y122_CQ),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_CQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y120_SLICE_X10Y120_BO5),
.O6(CLBLM_L_X8Y120_SLICE_X10Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffe3332ccdc0010)
  ) CLBLM_L_X8Y120_SLICE_X10Y120_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I4(CLBLM_L_X8Y126_SLICE_X11Y126_CQ),
.I5(CLBLM_R_X5Y119_SLICE_X7Y119_CQ),
.O5(CLBLM_L_X8Y120_SLICE_X10Y120_AO5),
.O6(CLBLM_L_X8Y120_SLICE_X10Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h77bb77bbddeeddee)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_DLUT (
.I0(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.I1(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y123_SLICE_X13Y123_AQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y122_SLICE_X15Y122_AQ),
.O5(CLBLM_L_X8Y120_SLICE_X11Y120_DO5),
.O6(CLBLM_L_X8Y120_SLICE_X11Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h66ffff6666ffff66)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_CLUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I1(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.I4(CLBLM_L_X10Y124_SLICE_X13Y124_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y120_SLICE_X11Y120_CO5),
.O6(CLBLM_L_X8Y120_SLICE_X11Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5aa5a5a5a55a5a)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_BLUT (
.I0(CLBLM_L_X8Y117_SLICE_X10Y117_AQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y123_SLICE_X13Y123_AQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y118_SLICE_X8Y118_BQ),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.O5(CLBLM_L_X8Y120_SLICE_X11Y120_BO5),
.O6(CLBLM_L_X8Y120_SLICE_X11Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffbbeebbee)
  ) CLBLM_L_X8Y120_SLICE_X11Y120_ALUT (
.I0(CLBLM_L_X8Y120_SLICE_X11Y120_DO6),
.I1(CLBLM_R_X7Y118_SLICE_X8Y118_BQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y121_SLICE_X12Y121_BQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y120_SLICE_X11Y120_CO6),
.O5(CLBLM_L_X8Y120_SLICE_X11Y120_AO5),
.O6(CLBLM_L_X8Y120_SLICE_X11Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X10Y121_BO6),
.Q(CLBLM_L_X8Y121_SLICE_X10Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X10Y121_CO6),
.Q(CLBLM_L_X8Y121_SLICE_X10Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aa00fc00fc00)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_DLUT (
.I0(CLBLM_R_X3Y122_SLICE_X2Y122_A5Q),
.I1(CLBLM_L_X8Y121_SLICE_X10Y121_CQ),
.I2(CLBLL_L_X4Y122_SLICE_X5Y122_DQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X10Y122_SLICE_X13Y122_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y121_SLICE_X10Y121_DO5),
.O6(CLBLM_L_X8Y121_SLICE_X10Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heafac0f0faeaf0c0)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y121_SLICE_X10Y121_CQ),
.I2(CLBLM_L_X8Y118_SLICE_X10Y118_AO5),
.I3(CLBLM_L_X8Y124_SLICE_X10Y124_CO6),
.I4(CLBLM_R_X7Y119_SLICE_X9Y119_AQ),
.I5(CLBLM_R_X7Y119_SLICE_X9Y119_CO6),
.O5(CLBLM_L_X8Y121_SLICE_X10Y121_CO5),
.O6(CLBLM_L_X8Y121_SLICE_X10Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff001111ff002222)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_BLUT (
.I0(CLBLM_L_X8Y121_SLICE_X10Y121_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(CLBLM_L_X8Y126_SLICE_X11Y126_B5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y119_SLICE_X4Y119_CQ),
.O5(CLBLM_L_X8Y121_SLICE_X10Y121_BO5),
.O6(CLBLM_L_X8Y121_SLICE_X10Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0cc88cc88cc88)
  ) CLBLM_L_X8Y121_SLICE_X10Y121_ALUT (
.I0(CLBLM_R_X11Y122_SLICE_X14Y122_DQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.I3(CLBLM_L_X10Y126_SLICE_X12Y126_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y121_SLICE_X10Y121_AO5),
.O6(CLBLM_L_X8Y121_SLICE_X10Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X11Y121_AO6),
.Q(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X11Y121_BO6),
.Q(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X11Y121_CO6),
.Q(CLBLM_L_X8Y121_SLICE_X11Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heaeafbea11111111)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_DLUT (
.I0(CLBLM_R_X3Y123_SLICE_X2Y123_DQ),
.I1(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.I2(CLBLM_L_X8Y121_SLICE_X10Y121_DO6),
.I3(CLBLL_L_X4Y128_SLICE_X4Y128_AO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y121_SLICE_X11Y121_DO5),
.O6(CLBLM_L_X8Y121_SLICE_X11Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff888800008888)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y121_SLICE_X11Y121_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y120_SLICE_X8Y120_AQ),
.O5(CLBLM_L_X8Y121_SLICE_X11Y121_CO5),
.O6(CLBLM_L_X8Y121_SLICE_X11Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccf044f044)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.I2(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.O5(CLBLM_L_X8Y121_SLICE_X11Y121_BO5),
.O6(CLBLM_L_X8Y121_SLICE_X11Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccca0ffa000)
  ) CLBLM_L_X8Y121_SLICE_X11Y121_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y120_SLICE_X7Y120_BQ),
.I2(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.I3(CLBLM_L_X8Y123_SLICE_X10Y123_DO6),
.I4(CLBLM_R_X11Y122_SLICE_X15Y122_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y121_SLICE_X11Y121_AO5),
.O6(CLBLM_L_X8Y121_SLICE_X11Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X10Y122_AO5),
.Q(CLBLM_L_X8Y122_SLICE_X10Y122_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X10Y122_AO6),
.Q(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X13Y122_BO6),
.Q(CLBLM_L_X8Y122_SLICE_X10Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffcfffc)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y122_SLICE_X13Y122_CQ),
.I2(CLBLM_L_X8Y122_SLICE_X10Y122_A5Q),
.I3(CLBLM_R_X5Y123_SLICE_X6Y123_CQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y122_SLICE_X12Y122_BQ),
.O5(CLBLM_L_X8Y122_SLICE_X10Y122_DO5),
.O6(CLBLM_L_X8Y122_SLICE_X10Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffafffa)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_CLUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_BQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y121_SLICE_X9Y121_B5Q),
.I3(CLBLM_L_X10Y122_SLICE_X13Y122_DQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y124_SLICE_X10Y124_BQ),
.O5(CLBLM_L_X8Y122_SLICE_X10Y122_CO5),
.O6(CLBLM_L_X8Y122_SLICE_X10Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_BLUT (
.I0(CLBLM_L_X8Y122_SLICE_X11Y122_CO6),
.I1(CLBLM_L_X10Y126_SLICE_X12Y126_CQ),
.I2(CLBLM_R_X5Y124_SLICE_X7Y124_C5Q),
.I3(CLBLL_L_X4Y122_SLICE_X4Y122_DQ),
.I4(CLBLM_L_X8Y122_SLICE_X11Y122_AQ),
.I5(CLBLM_L_X8Y122_SLICE_X10Y122_CO6),
.O5(CLBLM_L_X8Y122_SLICE_X10Y122_BO5),
.O6(CLBLM_L_X8Y122_SLICE_X10Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00f00c5c5c0c0)
  ) CLBLM_L_X8Y122_SLICE_X10Y122_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y122_SLICE_X7Y122_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(CLBLM_L_X8Y120_SLICE_X10Y120_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y122_SLICE_X10Y122_AO5),
.O6(CLBLM_L_X8Y122_SLICE_X10Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X11Y122_AO5),
.Q(CLBLM_L_X8Y122_SLICE_X11Y122_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y122_SLICE_X11Y122_AO6),
.Q(CLBLM_L_X8Y122_SLICE_X11Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffefefefe)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_DLUT (
.I0(CLBLM_L_X10Y122_SLICE_X13Y122_C5Q),
.I1(CLBLM_L_X10Y119_SLICE_X12Y119_BQ),
.I2(CLBLM_L_X10Y126_SLICE_X13Y126_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y125_SLICE_X6Y125_BQ),
.O5(CLBLM_L_X8Y122_SLICE_X11Y122_DO5),
.O6(CLBLM_L_X8Y122_SLICE_X11Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_CLUT (
.I0(CLBLM_L_X8Y123_SLICE_X11Y123_BQ),
.I1(CLBLM_L_X10Y122_SLICE_X12Y122_DO6),
.I2(CLBLM_L_X8Y122_SLICE_X10Y122_DO6),
.I3(CLBLM_L_X10Y121_SLICE_X12Y121_DQ),
.I4(CLBLM_L_X8Y122_SLICE_X11Y122_DO6),
.I5(CLBLL_L_X4Y123_SLICE_X5Y123_BQ),
.O5(CLBLM_L_X8Y122_SLICE_X11Y122_CO5),
.O6(CLBLM_L_X8Y122_SLICE_X11Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa8faf00000000)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_BLUT (
.I0(CLBLM_L_X8Y123_SLICE_X11Y123_DO5),
.I1(CLBLL_L_X4Y128_SLICE_X4Y128_AO6),
.I2(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X3Y123_SLICE_X2Y123_DQ),
.I5(CLBLM_L_X8Y118_SLICE_X10Y118_AO5),
.O5(CLBLM_L_X8Y122_SLICE_X11Y122_BO5),
.O6(CLBLM_L_X8Y122_SLICE_X11Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0cc00ff00aaaa)
  ) CLBLM_L_X8Y122_SLICE_X11Y122_ALUT (
.I0(CLBLM_R_X5Y128_SLICE_X7Y128_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y118_SLICE_X8Y118_AQ),
.I3(CLBLM_L_X10Y122_SLICE_X13Y122_C5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y122_SLICE_X11Y122_AO5),
.O6(CLBLM_L_X8Y122_SLICE_X11Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X10Y123_CO5),
.Q(CLBLM_L_X8Y123_SLICE_X10Y123_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X10Y123_AO6),
.Q(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X10Y123_BO6),
.Q(CLBLM_L_X8Y123_SLICE_X10Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X10Y123_CO6),
.Q(CLBLM_L_X8Y123_SLICE_X10Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0004000400040004)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_DLUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.I1(CLBLL_L_X2Y121_SLICE_X0Y121_AQ),
.I2(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y123_SLICE_X10Y123_DO5),
.O6(CLBLM_L_X8Y123_SLICE_X10Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaff00ccccf0f0)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_CLUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.I1(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(CLBLM_L_X8Y122_SLICE_X10Y122_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y123_SLICE_X10Y123_CO5),
.O6(CLBLM_L_X8Y123_SLICE_X10Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0afaca0a0)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_BLUT (
.I0(CLBLM_R_X11Y124_SLICE_X14Y124_CQ),
.I1(CLBLM_L_X8Y123_SLICE_X10Y123_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y122_SLICE_X9Y122_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.O5(CLBLM_L_X8Y123_SLICE_X10Y123_BO5),
.O6(CLBLM_L_X8Y123_SLICE_X10Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffcfc0cac0)
  ) CLBLM_L_X8Y123_SLICE_X10Y123_ALUT (
.I0(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I1(CLBLL_L_X4Y123_SLICE_X5Y123_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X7Y120_SLICE_X9Y120_BO6),
.O5(CLBLM_L_X8Y123_SLICE_X10Y123_AO5),
.O6(CLBLM_L_X8Y123_SLICE_X10Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X11Y123_CO5),
.Q(CLBLM_L_X8Y123_SLICE_X11Y123_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X11Y123_AO6),
.Q(CLBLM_L_X8Y123_SLICE_X11Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X11Y123_BO6),
.Q(CLBLM_L_X8Y123_SLICE_X11Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y123_SLICE_X11Y123_CO6),
.Q(CLBLM_L_X8Y123_SLICE_X11Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f000acacacac)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_DLUT (
.I0(CLBLM_L_X10Y126_SLICE_X12Y126_CQ),
.I1(CLBLM_L_X10Y123_SLICE_X12Y123_BQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.I4(CLBLM_L_X8Y124_SLICE_X10Y124_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y123_SLICE_X11Y123_DO5),
.O6(CLBLM_L_X8Y123_SLICE_X11Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0f000fa0a)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_CLUT (
.I0(CLBLM_L_X8Y123_SLICE_X11Y123_C5Q),
.I1(CLBLM_L_X8Y123_SLICE_X10Y123_C5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y127_SLICE_X12Y127_DQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y123_SLICE_X11Y123_CO5),
.O6(CLBLM_L_X8Y123_SLICE_X11Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aaaacccc)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_BLUT (
.I0(CLBLM_L_X8Y123_SLICE_X11Y123_CQ),
.I1(CLBLM_L_X10Y126_SLICE_X12Y126_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y123_SLICE_X11Y123_BO5),
.O6(CLBLM_L_X8Y123_SLICE_X11Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f5f5f000050500)
  ) CLBLM_L_X8Y123_SLICE_X11Y123_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y123_SLICE_X11Y123_DO5),
.I4(CLBLM_R_X3Y120_SLICE_X2Y120_CQ),
.I5(CLBLM_L_X10Y124_SLICE_X13Y124_C5Q),
.O5(CLBLM_L_X8Y123_SLICE_X11Y123_AO5),
.O6(CLBLM_L_X8Y123_SLICE_X11Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X10Y124_BO5),
.Q(CLBLM_L_X8Y124_SLICE_X10Y124_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X10Y124_AO6),
.Q(CLBLM_L_X8Y124_SLICE_X10Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X10Y124_BO6),
.Q(CLBLM_L_X8Y124_SLICE_X10Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb8bbbbb88b88888)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_DLUT (
.I0(CLBLM_L_X8Y124_SLICE_X10Y124_BQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.I3(CLBLL_L_X4Y124_SLICE_X4Y124_DQ),
.I4(CLBLM_L_X10Y124_SLICE_X12Y124_DO6),
.I5(CLBLM_R_X7Y124_SLICE_X9Y124_AQ),
.O5(CLBLM_L_X8Y124_SLICE_X10Y124_DO5),
.O6(CLBLM_L_X8Y124_SLICE_X10Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6966a5aa6999a555)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_CLUT (
.I0(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.I1(CLBLM_R_X7Y124_SLICE_X8Y124_CO6),
.I2(CLBLM_R_X11Y125_SLICE_X14Y125_CQ),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_CQ),
.I4(CLBLM_L_X10Y124_SLICE_X12Y124_DO6),
.I5(CLBLM_R_X7Y124_SLICE_X9Y124_CO6),
.O5(CLBLM_L_X8Y124_SLICE_X10Y124_CO5),
.O6(CLBLM_L_X8Y124_SLICE_X10Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0cfc0c0fafa0a0a)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_BLUT (
.I0(CLBLM_L_X8Y126_SLICE_X11Y126_B5Q),
.I1(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y122_SLICE_X13Y122_DQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y124_SLICE_X10Y124_BO5),
.O6(CLBLM_L_X8Y124_SLICE_X10Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00a0000000a0)
  ) CLBLM_L_X8Y124_SLICE_X10Y124_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(CLBLM_L_X8Y124_SLICE_X10Y124_AQ),
.I3(CLBLM_R_X5Y124_SLICE_X7Y124_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y124_SLICE_X9Y124_AQ),
.O5(CLBLM_L_X8Y124_SLICE_X10Y124_AO5),
.O6(CLBLM_L_X8Y124_SLICE_X10Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X11Y124_AO6),
.Q(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X11Y124_BO6),
.Q(CLBLM_L_X8Y124_SLICE_X11Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff08f000ff08f000)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X3Y128_SLICE_X2Y128_AO6),
.I2(CLBLM_R_X3Y123_SLICE_X2Y123_DQ),
.I3(CLBLM_L_X8Y121_SLICE_X10Y121_DO5),
.I4(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y124_SLICE_X11Y124_DO5),
.O6(CLBLM_L_X8Y124_SLICE_X11Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfa00fa00fa00)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_CLUT (
.I0(CLBLM_L_X8Y123_SLICE_X10Y123_AQ),
.I1(CLBLM_L_X10Y124_SLICE_X13Y124_BQ),
.I2(CLBLM_R_X5Y124_SLICE_X6Y124_CQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y124_SLICE_X11Y124_CO5),
.O6(CLBLM_L_X8Y124_SLICE_X11Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf101f404f101f404)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y123_SLICE_X11Y123_BQ),
.I4(CLBLM_L_X8Y124_SLICE_X11Y124_CO5),
.I5(1'b1),
.O5(CLBLM_L_X8Y124_SLICE_X11Y124_BO5),
.O6(CLBLM_L_X8Y124_SLICE_X11Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00a0cccc00a0)
  ) CLBLM_L_X8Y124_SLICE_X11Y124_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y126_SLICE_X11Y126_BQ),
.I2(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.I3(CLBLM_R_X5Y124_SLICE_X7Y124_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y124_SLICE_X11Y124_AO5),
.O6(CLBLM_L_X8Y124_SLICE_X11Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X10Y125_AO6),
.Q(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X10Y125_CO6),
.Q(CLBLM_L_X8Y125_SLICE_X10Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X10Y125_DO6),
.Q(CLBLM_L_X8Y125_SLICE_X10Y125_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff00f3f3)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_DLUT (
.I0(1'b1),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_DQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y119_SLICE_X10Y119_CO6),
.O5(CLBLM_L_X8Y125_SLICE_X10Y125_DO5),
.O6(CLBLM_L_X8Y125_SLICE_X10Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc05055050)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.I2(CLBLM_L_X10Y125_SLICE_X12Y125_CQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y125_SLICE_X10Y125_BO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y125_SLICE_X10Y125_CO5),
.O6(CLBLM_L_X8Y125_SLICE_X10Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcf80c08cc88cc88)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_BLUT (
.I0(CLBLM_L_X10Y125_SLICE_X12Y125_DQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y122_SLICE_X10Y122_A5Q),
.I4(CLBLM_R_X7Y118_SLICE_X8Y118_DQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y125_SLICE_X10Y125_BO5),
.O6(CLBLM_L_X8Y125_SLICE_X10Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55aa00fe54ba10)
  ) CLBLM_L_X8Y125_SLICE_X10Y125_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I2(CLBLM_L_X8Y125_SLICE_X10Y125_AQ),
.I3(CLBLM_R_X11Y126_SLICE_X15Y126_CQ),
.I4(CLBLM_R_X7Y122_SLICE_X9Y122_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X8Y125_SLICE_X10Y125_AO5),
.O6(CLBLM_L_X8Y125_SLICE_X10Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X11Y125_AO6),
.Q(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X11Y125_BO6),
.Q(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X11Y125_CO6),
.Q(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcfcfcfcdcfcdc)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X3Y123_SLICE_X2Y123_DQ),
.I2(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.I3(CLBLM_R_X3Y128_SLICE_X2Y128_AO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y125_SLICE_X6Y125_CO6),
.O5(CLBLM_L_X8Y125_SLICE_X11Y125_DO5),
.O6(CLBLM_L_X8Y125_SLICE_X11Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafacacafa0aca0)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_CLUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_CQ),
.I1(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y124_SLICE_X11Y124_DO6),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.O5(CLBLM_L_X8Y125_SLICE_X11Y125_CO5),
.O6(CLBLM_L_X8Y125_SLICE_X11Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeee00000eee0)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_BLUT (
.I0(CLBLM_R_X7Y124_SLICE_X8Y124_DO6),
.I1(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.I2(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y127_SLICE_X11Y127_CQ),
.O5(CLBLM_L_X8Y125_SLICE_X11Y125_BO5),
.O6(CLBLM_L_X8Y125_SLICE_X11Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd11dd11dc10dc10)
  ) CLBLM_L_X8Y125_SLICE_X11Y125_ALUT (
.I0(CLBLM_L_X10Y129_SLICE_X13Y129_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.I3(CLBLM_L_X10Y119_SLICE_X12Y119_BQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y126_SLICE_X9Y126_DQ),
.O5(CLBLM_L_X8Y125_SLICE_X11Y125_AO5),
.O6(CLBLM_L_X8Y125_SLICE_X11Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X5Y118_SLICE_X7Y118_AQ),
.Q(CLBLM_L_X8Y126_SLICE_X10Y126_AQ),
.R(CLBLM_L_X8Y131_SLICE_X11Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffefffeff)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_DLUT (
.I0(CLBLM_L_X10Y125_SLICE_X13Y125_AQ),
.I1(CLBLM_L_X8Y127_SLICE_X10Y127_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_DQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y127_SLICE_X12Y127_CQ),
.O5(CLBLM_L_X8Y126_SLICE_X10Y126_DO5),
.O6(CLBLM_L_X8Y126_SLICE_X10Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000800000008000)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_CLUT (
.I0(CLBLM_R_X7Y125_SLICE_X8Y125_CQ),
.I1(CLBLM_L_X8Y127_SLICE_X10Y127_CQ),
.I2(CLBLM_L_X8Y127_SLICE_X11Y127_DQ),
.I3(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.I4(CLBLM_L_X8Y126_SLICE_X10Y126_DO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y126_SLICE_X10Y126_CO5),
.O6(CLBLM_L_X8Y126_SLICE_X10Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffefe)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_BLUT (
.I0(CLBLM_R_X7Y119_SLICE_X9Y119_AQ),
.I1(CLBLM_L_X8Y124_SLICE_X11Y124_BQ),
.I2(CLBLL_L_X4Y125_SLICE_X4Y125_AQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y126_SLICE_X10Y126_AO6),
.I5(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.O5(CLBLM_L_X8Y126_SLICE_X10Y126_BO5),
.O6(CLBLM_L_X8Y126_SLICE_X10Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffeff55005500)
  ) CLBLM_L_X8Y126_SLICE_X10Y126_ALUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_L_X10Y125_SLICE_X12Y125_CQ),
.I2(CLBLM_L_X8Y125_SLICE_X10Y125_CQ),
.I3(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.I4(CLBLM_L_X10Y124_SLICE_X13Y124_DQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y126_SLICE_X10Y126_AO5),
.O6(CLBLM_L_X8Y126_SLICE_X10Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y126_SLICE_X11Y126_BO5),
.Q(CLBLM_L_X8Y126_SLICE_X11Y126_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y126_SLICE_X11Y126_AO6),
.Q(CLBLM_L_X8Y126_SLICE_X11Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y126_SLICE_X11Y126_BO6),
.Q(CLBLM_L_X8Y126_SLICE_X11Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y126_SLICE_X11Y126_CO6),
.Q(CLBLM_L_X8Y126_SLICE_X11Y126_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y126_SLICE_X11Y126_DO6),
.Q(CLBLM_L_X8Y126_SLICE_X11Y126_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa33aa30aa00aa00)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_DLUT (
.I0(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X8Y126_SLICE_X11Y126_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y125_SLICE_X11Y125_DO6),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.O5(CLBLM_L_X8Y126_SLICE_X11Y126_DO5),
.O6(CLBLM_L_X8Y126_SLICE_X11Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f0f3f003000300)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y127_SLICE_X15Y127_BO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y126_SLICE_X11Y126_BQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y124_SLICE_X11Y124_BQ),
.O5(CLBLM_L_X8Y126_SLICE_X11Y126_CO5),
.O6(CLBLM_L_X8Y126_SLICE_X11Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf2f20202ff0ff000)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_BLUT (
.I0(CLBLM_L_X10Y127_SLICE_X13Y127_DQ),
.I1(CLBLM_R_X11Y127_SLICE_X15Y127_BO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y124_SLICE_X10Y124_BQ),
.I4(CLBLM_R_X5Y126_SLICE_X7Y126_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y126_SLICE_X11Y126_BO5),
.O6(CLBLM_L_X8Y126_SLICE_X11Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f2f22222)
  ) CLBLM_L_X8Y126_SLICE_X11Y126_ALUT (
.I0(CLBLM_L_X8Y126_SLICE_X10Y126_CO6),
.I1(CLBLM_L_X8Y126_SLICE_X10Y126_BO6),
.I2(CLBLM_L_X8Y126_SLICE_X11Y126_AQ),
.I3(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y126_SLICE_X11Y126_AO5),
.O6(CLBLM_L_X8Y126_SLICE_X11Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X10Y127_AO6),
.Q(CLBLM_L_X8Y127_SLICE_X10Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X10Y127_BO6),
.Q(CLBLM_L_X8Y127_SLICE_X10Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X10Y127_CO6),
.Q(CLBLM_L_X8Y127_SLICE_X10Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0ff0f0f0f0)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X4Y125_SLICE_X4Y125_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.O5(CLBLM_L_X8Y127_SLICE_X10Y127_DO5),
.O6(CLBLM_L_X8Y127_SLICE_X10Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00000f000f00)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X8Y127_SLICE_X10Y127_BQ),
.I4(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y127_SLICE_X10Y127_CO5),
.O6(CLBLM_L_X8Y127_SLICE_X10Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0300c03c)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_BLUT (
.I0(CLBLM_R_X5Y128_SLICE_X7Y128_AQ),
.I1(CLBLM_L_X8Y127_SLICE_X10Y127_BQ),
.I2(CLBLM_L_X10Y127_SLICE_X12Y127_CQ),
.I3(CLBLM_L_X8Y127_SLICE_X10Y127_DO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y127_SLICE_X10Y127_BO5),
.O6(CLBLM_L_X8Y127_SLICE_X10Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5500ccccf5a0)
  ) CLBLM_L_X8Y127_SLICE_X10Y127_ALUT (
.I0(CLBLM_R_X5Y130_SLICE_X7Y130_DO6),
.I1(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.I2(CLBLM_L_X8Y127_SLICE_X10Y127_AQ),
.I3(CLBLM_R_X7Y127_SLICE_X9Y127_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y130_SLICE_X8Y130_CO6),
.O5(CLBLM_L_X8Y127_SLICE_X10Y127_AO5),
.O6(CLBLM_L_X8Y127_SLICE_X10Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X11Y127_AO6),
.Q(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X11Y127_BO6),
.Q(CLBLM_L_X8Y127_SLICE_X11Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X11Y127_CO6),
.Q(CLBLM_L_X8Y127_SLICE_X11Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y127_SLICE_X11Y127_DO6),
.Q(CLBLM_L_X8Y127_SLICE_X11Y127_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0000c3c3)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_DLUT (
.I0(CLBLM_R_X7Y127_SLICE_X9Y127_CQ),
.I1(CLBLM_R_X7Y119_SLICE_X9Y119_AQ),
.I2(CLBLM_L_X10Y124_SLICE_X12Y124_BO5),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y127_SLICE_X11Y127_DO5),
.O6(CLBLM_L_X8Y127_SLICE_X11Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff000c0c0c0c)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y124_SLICE_X6Y124_A5Q),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X8Y127_SLICE_X11Y127_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y127_SLICE_X11Y127_CO5),
.O6(CLBLM_L_X8Y127_SLICE_X11Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf505f000fd0df808)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_BLUT (
.I0(CLBLM_R_X5Y130_SLICE_X7Y130_DO6),
.I1(CLBLM_L_X8Y127_SLICE_X11Y127_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y118_SLICE_X11Y118_BQ),
.I4(CLBLM_L_X8Y128_SLICE_X11Y128_AQ),
.I5(CLBLM_R_X7Y130_SLICE_X8Y130_CO6),
.O5(CLBLM_L_X8Y127_SLICE_X11Y127_BO5),
.O6(CLBLM_L_X8Y127_SLICE_X11Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00ccaaaaf0cc)
  ) CLBLM_L_X8Y127_SLICE_X11Y127_ALUT (
.I0(CLBLM_R_X7Y123_SLICE_X9Y123_CQ),
.I1(CLBLM_L_X8Y127_SLICE_X11Y127_BQ),
.I2(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I3(CLBLM_R_X5Y130_SLICE_X7Y130_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y130_SLICE_X8Y130_CO6),
.O5(CLBLM_L_X8Y127_SLICE_X11Y127_AO5),
.O6(CLBLM_L_X8Y127_SLICE_X11Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X10Y128_AO6),
.Q(CLBLM_L_X8Y128_SLICE_X10Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X10Y128_BO6),
.Q(CLBLM_L_X8Y128_SLICE_X10Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X10Y128_CO6),
.Q(CLBLM_L_X8Y128_SLICE_X10Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00ff00ff0a5f00f)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_DLUT (
.I0(CLBLM_L_X8Y127_SLICE_X11Y127_BQ),
.I1(1'b1),
.I2(CLBLM_L_X8Y128_SLICE_X10Y128_BQ),
.I3(CLBLM_R_X7Y131_SLICE_X9Y131_CO6),
.I4(CLBLM_L_X8Y129_SLICE_X10Y129_DO6),
.I5(CLBLM_R_X7Y128_SLICE_X9Y128_DO6),
.O5(CLBLM_L_X8Y128_SLICE_X10Y128_DO5),
.O6(CLBLM_L_X8Y128_SLICE_X10Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000d0c0d0c0)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_CLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_L_X8Y128_SLICE_X10Y128_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.I4(CLBLM_R_X5Y120_SLICE_X7Y120_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y128_SLICE_X10Y128_CO5),
.O6(CLBLM_L_X8Y128_SLICE_X10Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4044f0ff4044f0ff)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_BLUT (
.I0(CLBLM_L_X8Y128_SLICE_X10Y128_DO6),
.I1(CLBLM_R_X7Y131_SLICE_X9Y131_BO6),
.I2(CLBLL_L_X4Y120_SLICE_X5Y120_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y131_SLICE_X8Y131_CO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y128_SLICE_X10Y128_BO5),
.O6(CLBLM_L_X8Y128_SLICE_X10Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4500cfcf4500cfcf)
  ) CLBLM_L_X8Y128_SLICE_X10Y128_ALUT (
.I0(CLBLM_L_X8Y129_SLICE_X10Y129_CO6),
.I1(CLBLL_L_X2Y121_SLICE_X0Y121_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y131_SLICE_X9Y131_BO6),
.I4(CLBLM_R_X7Y131_SLICE_X8Y131_CO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y128_SLICE_X10Y128_AO5),
.O6(CLBLM_L_X8Y128_SLICE_X10Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X11Y128_AO6),
.Q(CLBLM_L_X8Y128_SLICE_X11Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X11Y128_BO6),
.Q(CLBLM_L_X8Y128_SLICE_X11Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X11Y128_CO6),
.Q(CLBLM_L_X8Y128_SLICE_X11Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y128_SLICE_X11Y128_DO6),
.Q(CLBLM_L_X8Y128_SLICE_X11Y128_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0cfc0cfc0c0c0c0)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y127_SLICE_X11Y127_DQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y127_SLICE_X11Y127_CQ),
.O5(CLBLM_L_X8Y128_SLICE_X11Y128_DO5),
.O6(CLBLM_L_X8Y128_SLICE_X11Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7700550077775555)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_CLUT (
.I0(CLBLM_R_X7Y131_SLICE_X8Y131_CO6),
.I1(CLBLM_L_X8Y129_SLICE_X11Y129_CO6),
.I2(1'b1),
.I3(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.I4(CLBLM_R_X7Y131_SLICE_X9Y131_BO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y128_SLICE_X11Y128_CO5),
.O6(CLBLM_L_X8Y128_SLICE_X11Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0f5a0e4e4f5a0)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y128_SLICE_X11Y128_BQ),
.I2(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I3(CLBLM_R_X7Y128_SLICE_X9Y128_AQ),
.I4(CLBLM_R_X5Y130_SLICE_X7Y130_DO6),
.I5(CLBLM_R_X7Y130_SLICE_X8Y130_CO6),
.O5(CLBLM_L_X8Y128_SLICE_X11Y128_BO5),
.O6(CLBLM_L_X8Y128_SLICE_X11Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff3bff08003b0008)
  ) CLBLM_L_X8Y128_SLICE_X11Y128_ALUT (
.I0(CLBLM_L_X8Y128_SLICE_X11Y128_AQ),
.I1(CLBLM_R_X5Y130_SLICE_X7Y130_DO6),
.I2(CLBLM_R_X7Y130_SLICE_X8Y130_CO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.I5(CLBLM_R_X5Y128_SLICE_X6Y128_DQ),
.O5(CLBLM_L_X8Y128_SLICE_X11Y128_AO5),
.O6(CLBLM_L_X8Y128_SLICE_X11Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X5Y124_SLICE_X6Y124_A5Q),
.Q(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.R(CLBLM_L_X8Y131_SLICE_X11Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h222a000000004440)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_DLUT (
.I0(CLBLM_L_X8Y129_SLICE_X11Y129_AQ),
.I1(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.I2(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.I3(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I4(CLBLM_L_X8Y128_SLICE_X10Y128_AQ),
.I5(CLBLM_R_X7Y129_SLICE_X9Y129_AQ),
.O5(CLBLM_L_X8Y129_SLICE_X10Y129_DO5),
.O6(CLBLM_L_X8Y129_SLICE_X10Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff2000dfff0200fd)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_CLUT (
.I0(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.I1(CLBLM_R_X7Y128_SLICE_X9Y128_DO6),
.I2(CLBLM_R_X7Y130_SLICE_X9Y130_CO6),
.I3(CLBLM_R_X7Y131_SLICE_X9Y131_CO6),
.I4(CLBLM_L_X8Y128_SLICE_X10Y128_AQ),
.I5(CLBLM_L_X8Y129_SLICE_X11Y129_AQ),
.O5(CLBLM_L_X8Y129_SLICE_X10Y129_CO5),
.O6(CLBLM_L_X8Y129_SLICE_X10Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4555555555555455)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_BLUT (
.I0(CLBLM_R_X7Y131_SLICE_X9Y131_CO6),
.I1(CLBLM_R_X7Y128_SLICE_X9Y128_DO6),
.I2(CLBLM_L_X8Y128_SLICE_X10Y128_AQ),
.I3(CLBLM_L_X8Y128_SLICE_X11Y128_AQ),
.I4(CLBLM_L_X8Y129_SLICE_X11Y129_AQ),
.I5(CLBLM_R_X7Y130_SLICE_X9Y130_CO6),
.O5(CLBLM_L_X8Y129_SLICE_X10Y129_BO5),
.O6(CLBLM_L_X8Y129_SLICE_X10Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000001)
  ) CLBLM_L_X8Y129_SLICE_X10Y129_ALUT (
.I0(CLBLM_R_X7Y130_SLICE_X9Y130_CO6),
.I1(CLBLM_L_X8Y128_SLICE_X10Y128_BQ),
.I2(CLBLM_L_X8Y128_SLICE_X10Y128_AQ),
.I3(CLBLM_R_X7Y129_SLICE_X9Y129_AQ),
.I4(CLBLM_L_X8Y129_SLICE_X11Y129_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X10Y129_AO5),
.O6(CLBLM_L_X8Y129_SLICE_X10Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y129_SLICE_X11Y129_BO5),
.Q(CLBLM_L_X8Y129_SLICE_X11Y129_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y129_SLICE_X11Y129_AO6),
.Q(CLBLM_L_X8Y129_SLICE_X11Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y129_SLICE_X11Y129_BO6),
.Q(CLBLM_L_X8Y129_SLICE_X11Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc66cc66cc33cc33)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_DLUT (
.I0(CLBLM_R_X7Y128_SLICE_X9Y128_DO6),
.I1(CLBLM_L_X8Y129_SLICE_X11Y129_AQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y131_SLICE_X9Y131_CO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.O5(CLBLM_L_X8Y129_SLICE_X11Y129_DO5),
.O6(CLBLM_L_X8Y129_SLICE_X11Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa55a55595)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_CLUT (
.I0(CLBLM_L_X8Y128_SLICE_X11Y128_CQ),
.I1(CLBLM_L_X8Y129_SLICE_X10Y129_AO5),
.I2(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I3(CLBLM_R_X7Y128_SLICE_X9Y128_DO6),
.I4(CLBLM_L_X8Y129_SLICE_X10Y129_AO6),
.I5(CLBLM_R_X7Y131_SLICE_X9Y131_CO6),
.O5(CLBLM_L_X8Y129_SLICE_X11Y129_CO5),
.O6(CLBLM_L_X8Y129_SLICE_X11Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa0ffa0ffffc0c0)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_BLUT (
.I0(CLBLM_R_X7Y127_SLICE_X9Y127_AQ),
.I1(CLBLM_R_X5Y129_SLICE_X6Y129_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y128_SLICE_X13Y128_DO6),
.I4(CLBLM_R_X5Y129_SLICE_X7Y129_BO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y129_SLICE_X11Y129_BO5),
.O6(CLBLM_L_X8Y129_SLICE_X11Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5500ffff05000f0f)
  ) CLBLM_L_X8Y129_SLICE_X11Y129_ALUT (
.I0(CLBLM_L_X8Y129_SLICE_X11Y129_DO6),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y131_SLICE_X9Y131_BO6),
.I4(CLBLM_R_X7Y131_SLICE_X8Y131_CO6),
.I5(CLBLM_R_X7Y123_SLICE_X9Y123_BQ),
.O5(CLBLM_L_X8Y129_SLICE_X11Y129_AO5),
.O6(CLBLM_L_X8Y129_SLICE_X11Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X10Y130_AO6),
.Q(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X10Y130_BO6),
.Q(CLBLM_L_X8Y130_SLICE_X10Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X10Y130_CO6),
.Q(CLBLM_L_X8Y130_SLICE_X10Y130_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cd00ef00ff00ff)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_DLUT (
.I0(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I1(CLBLM_R_X7Y128_SLICE_X9Y128_DO6),
.I2(CLBLM_L_X8Y131_SLICE_X10Y131_BO5),
.I3(CLBLM_R_X7Y131_SLICE_X9Y131_CO6),
.I4(CLBLM_L_X8Y131_SLICE_X10Y131_AO5),
.I5(CLBLM_R_X7Y127_SLICE_X9Y127_CQ),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_DO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd0d770755055505)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_CLUT (
.I0(CLBLM_R_X7Y131_SLICE_X8Y131_CO6),
.I1(CLBLM_L_X8Y130_SLICE_X10Y130_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y125_SLICE_X12Y125_DQ),
.I4(CLBLM_L_X8Y130_SLICE_X10Y130_DO6),
.I5(CLBLM_R_X7Y131_SLICE_X9Y131_BO6),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_CO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff0fcc0cff0f)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y131_SLICE_X9Y131_BO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y124_SLICE_X13Y124_A5Q),
.I4(CLBLM_R_X7Y131_SLICE_X8Y131_CO6),
.I5(CLBLM_L_X8Y131_SLICE_X10Y131_CO6),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_BO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaf0aafcaafc)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_ALUT (
.I0(CLBLM_L_X8Y130_SLICE_X10Y130_CQ),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_AO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000c000c555d000c)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_DLUT (
.I0(CLBLM_L_X8Y130_SLICE_X11Y130_AO6),
.I1(CLBLM_R_X7Y129_SLICE_X8Y129_CQ),
.I2(CLBLM_L_X8Y130_SLICE_X11Y130_CO6),
.I3(CLBLM_L_X8Y130_SLICE_X11Y130_AO5),
.I4(CLBLM_R_X7Y125_SLICE_X8Y125_AQ),
.I5(CLBLM_L_X8Y130_SLICE_X11Y130_BO6),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_DO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffd)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_CLUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(RIOB33_X105Y129_IOB_X1Y130_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y135_IOB_X1Y135_I),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_CO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffff7f)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y135_IOB_X1Y136_I),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(RIOB33_X105Y129_IOB_X1Y130_I),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(RIOB33_X105Y135_IOB_X1Y135_I),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_BO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fffffffff0fff)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_AO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.Q(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.R(CLBLM_L_X8Y131_SLICE_X11Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0d05050508000000)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_DLUT (
.I0(CLBLM_L_X8Y130_SLICE_X10Y130_BQ),
.I1(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I2(CLBLM_R_X7Y128_SLICE_X9Y128_DO6),
.I3(CLBLM_L_X8Y131_SLICE_X10Y131_AO5),
.I4(CLBLM_L_X8Y130_SLICE_X10Y130_CQ),
.I5(CLBLM_L_X8Y131_SLICE_X10Y131_BO6),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_DO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0e000000f1ff)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_CLUT (
.I0(CLBLM_L_X8Y131_SLICE_X10Y131_AO6),
.I1(CLBLM_L_X8Y131_SLICE_X10Y131_BO6),
.I2(CLBLM_R_X7Y128_SLICE_X9Y128_DO6),
.I3(CLBLM_L_X8Y127_SLICE_X10Y127_AQ),
.I4(CLBLM_R_X7Y131_SLICE_X9Y131_CO6),
.I5(CLBLM_L_X8Y130_SLICE_X10Y130_BQ),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_CO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010011001100)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_BLUT (
.I0(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I1(CLBLM_L_X8Y128_SLICE_X11Y128_CQ),
.I2(CLBLM_L_X8Y130_SLICE_X10Y130_CQ),
.I3(CLBLM_L_X8Y129_SLICE_X10Y129_AO5),
.I4(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_BO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000088008800)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_ALUT (
.I0(CLBLM_L_X8Y129_SLICE_X10Y129_AO6),
.I1(CLBLM_L_X8Y128_SLICE_X11Y128_CQ),
.I2(CLBLM_L_X8Y130_SLICE_X10Y130_CQ),
.I3(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I4(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_AO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X11Y131_AO6),
.Q(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5511551155115511)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(1'b1),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_DO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00005400abff)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_CLUT (
.I0(CLBLM_R_X7Y128_SLICE_X9Y128_DO6),
.I1(CLBLM_L_X8Y131_SLICE_X10Y131_AO5),
.I2(CLBLM_L_X8Y131_SLICE_X10Y131_BO5),
.I3(CLBLM_L_X8Y128_SLICE_X11Y128_BQ),
.I4(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I5(CLBLM_R_X7Y131_SLICE_X9Y131_CO6),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_CO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff004f00ff007f)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_BLUT (
.I0(CLBLM_L_X8Y129_SLICE_X10Y129_AO6),
.I1(CLBLM_L_X8Y128_SLICE_X11Y128_CQ),
.I2(CLBLM_R_X7Y128_SLICE_X9Y128_AQ),
.I3(CLBLM_R_X7Y131_SLICE_X9Y131_CO6),
.I4(CLBLM_R_X7Y128_SLICE_X9Y128_DO6),
.I5(CLBLM_L_X8Y129_SLICE_X10Y129_AO5),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_BO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33033303bb0bbb0b)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_ALUT (
.I0(CLBLM_R_X7Y131_SLICE_X9Y131_BO6),
.I1(CLBLM_R_X7Y131_SLICE_X8Y131_CO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y130_SLICE_X14Y130_AQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y131_SLICE_X11Y131_CO6),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_AO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y117_SLICE_X12Y117_AO6),
.Q(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y117_SLICE_X12Y117_DO5),
.O6(CLBLM_L_X10Y117_SLICE_X12Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y117_SLICE_X12Y117_CO5),
.O6(CLBLM_L_X10Y117_SLICE_X12Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y117_SLICE_X12Y117_BO5),
.O6(CLBLM_L_X10Y117_SLICE_X12Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cca0cc00cc0a)
  ) CLBLM_L_X10Y117_SLICE_X12Y117_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X12Y126_SLICE_X16Y126_BQ),
.I2(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y126_SLICE_X9Y126_BQ),
.I5(CLBLM_L_X8Y117_SLICE_X10Y117_CO6),
.O5(CLBLM_L_X10Y117_SLICE_X12Y117_AO5),
.O6(CLBLM_L_X10Y117_SLICE_X12Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y117_SLICE_X13Y117_DO5),
.O6(CLBLM_L_X10Y117_SLICE_X13Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y117_SLICE_X13Y117_CO5),
.O6(CLBLM_L_X10Y117_SLICE_X13Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y117_SLICE_X13Y117_BO5),
.O6(CLBLM_L_X10Y117_SLICE_X13Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y117_SLICE_X13Y117_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y117_SLICE_X13Y117_AO5),
.O6(CLBLM_L_X10Y117_SLICE_X13Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y118_SLICE_X12Y118_AO6),
.Q(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_DO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055ffff0055ffff)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_CLUT (
.I0(CLBLM_L_X8Y118_SLICE_X11Y118_CO5),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X10Y121_SLICE_X12Y121_CQ),
.I4(CLBLM_R_X3Y125_SLICE_X2Y125_BO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_CO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f0f5f0f5f0fff0)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_BLUT (
.I0(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I1(1'b1),
.I2(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.I3(CLBLM_R_X7Y118_SLICE_X9Y118_BO6),
.I4(CLBLM_L_X8Y118_SLICE_X11Y118_CO5),
.I5(CLBLM_L_X10Y121_SLICE_X12Y121_CQ),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_BO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf888f888f888f8f8)
  ) CLBLM_L_X10Y118_SLICE_X12Y118_ALUT (
.I0(CLBLM_L_X10Y128_SLICE_X12Y128_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y131_SLICE_X11Y131_DO6),
.I3(CLBLM_L_X10Y118_SLICE_X12Y118_BO6),
.I4(CLBLM_L_X8Y116_SLICE_X11Y116_AO6),
.I5(CLBLM_R_X7Y118_SLICE_X9Y118_BO6),
.O5(CLBLM_L_X10Y118_SLICE_X12Y118_AO5),
.O6(CLBLM_L_X10Y118_SLICE_X12Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y118_SLICE_X13Y118_AO6),
.Q(CLBLM_L_X10Y118_SLICE_X13Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_DO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_CO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0101010d0d0d0d01)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_BLUT (
.I0(CLBLM_L_X10Y120_SLICE_X13Y120_A5Q),
.I1(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I2(CLBLM_L_X10Y118_SLICE_X13Y118_AQ),
.I3(CLBLM_L_X8Y117_SLICE_X11Y117_AO6),
.I4(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I5(CLBLM_R_X5Y119_SLICE_X6Y119_CQ),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_BO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88dd88dd888888dd)
  ) CLBLM_L_X10Y118_SLICE_X13Y118_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y118_SLICE_X13Y118_BO6),
.I4(RIOB33_X105Y141_IOB_X1Y142_I),
.I5(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.O5(CLBLM_L_X10Y118_SLICE_X13Y118_AO5),
.O6(CLBLM_L_X10Y118_SLICE_X13Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y119_SLICE_X12Y119_AO6),
.Q(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y119_SLICE_X12Y119_BO6),
.Q(CLBLM_L_X10Y119_SLICE_X12Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y119_SLICE_X12Y119_CO6),
.Q(CLBLM_L_X10Y119_SLICE_X12Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y119_SLICE_X12Y119_DO6),
.Q(CLBLM_L_X10Y119_SLICE_X12Y119_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefe5454aaaa0000)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y119_SLICE_X12Y119_CQ),
.I2(CLBLM_L_X10Y119_SLICE_X12Y119_DQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y127_SLICE_X10Y127_CQ),
.I5(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_DO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5e4e4a0a0a0a0)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y119_SLICE_X12Y119_CQ),
.I2(CLBLM_R_X11Y122_SLICE_X14Y122_DQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y119_SLICE_X6Y119_CQ),
.I5(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_CO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd1d1c0c0d1d1c0c0)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y118_SLICE_X3Y118_BQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y122_SLICE_X12Y122_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_BO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeaafbaafc00f300)
  ) CLBLM_L_X10Y119_SLICE_X12Y119_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y118_SLICE_X12Y118_CO6),
.I2(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.I3(CLBLM_L_X8Y131_SLICE_X11Y131_DO6),
.I4(CLBLM_L_X8Y116_SLICE_X11Y116_AO6),
.I5(CLBLM_L_X10Y121_SLICE_X12Y121_CQ),
.O5(CLBLM_L_X10Y119_SLICE_X12Y119_AO5),
.O6(CLBLM_L_X10Y119_SLICE_X12Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y119_SLICE_X13Y119_AO6),
.Q(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y119_SLICE_X13Y119_BO6),
.Q(CLBLM_L_X10Y119_SLICE_X13Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333cfcfcccc)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y120_SLICE_X13Y120_CQ),
.I2(CLBLM_L_X10Y120_SLICE_X13Y120_DO6),
.I3(1'b1),
.I4(CLBLM_L_X8Y119_SLICE_X10Y119_DO6),
.I5(CLBLM_L_X10Y121_SLICE_X13Y121_AQ),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_DO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h005000af00330033)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_CLUT (
.I0(CLBLM_L_X8Y117_SLICE_X11Y117_AO6),
.I1(CLBLM_L_X10Y124_SLICE_X13Y124_D5Q),
.I2(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I3(CLBLM_L_X10Y123_SLICE_X13Y123_BQ),
.I4(CLBLM_L_X10Y119_SLICE_X12Y119_DQ),
.I5(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_CO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00f0f0cc00)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y119_SLICE_X13Y119_BQ),
.I2(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.I3(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y117_SLICE_X10Y117_BQ),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_BO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaccaac0aac0)
  ) CLBLM_L_X10Y119_SLICE_X13Y119_ALUT (
.I0(CLBLM_L_X10Y120_SLICE_X13Y120_BQ),
.I1(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I2(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y119_SLICE_X11Y119_CQ),
.O5(CLBLM_L_X10Y119_SLICE_X13Y119_AO5),
.O6(CLBLM_L_X10Y119_SLICE_X13Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X12Y120_AO6),
.Q(CLBLM_L_X10Y120_SLICE_X12Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X12Y120_BO6),
.Q(CLBLM_L_X10Y120_SLICE_X12Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X12Y120_CO6),
.Q(CLBLM_L_X10Y120_SLICE_X12Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2211112211222211)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_DLUT (
.I0(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_AQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y120_SLICE_X10Y120_CO6),
.I4(CLBLM_R_X11Y123_SLICE_X14Y123_AQ),
.I5(CLBLM_L_X8Y120_SLICE_X11Y120_BO6),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_DO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff8f8000008f80)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_CQ),
.I2(CLBLM_L_X8Y123_SLICE_X10Y123_DO6),
.I3(CLBLM_L_X10Y121_SLICE_X12Y121_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y128_SLICE_X10Y128_BQ),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_CO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcff0cfff8ff08)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X10Y120_SLICE_X12Y120_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y120_SLICE_X9Y120_AO6),
.I4(CLBLM_L_X10Y119_SLICE_X13Y119_BQ),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_BO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff500f5ffc400c4)
  ) CLBLM_L_X10Y120_SLICE_X12Y120_ALUT (
.I0(CLBLM_L_X10Y120_SLICE_X12Y120_DO6),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X7Y118_SLICE_X9Y118_BO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.O5(CLBLM_L_X10Y120_SLICE_X12Y120_AO5),
.O6(CLBLM_L_X10Y120_SLICE_X12Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X13Y120_AO5),
.Q(CLBLM_L_X10Y120_SLICE_X13Y120_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X13Y120_AO6),
.Q(CLBLM_L_X10Y120_SLICE_X13Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X13Y120_BO6),
.Q(CLBLM_L_X10Y120_SLICE_X13Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y120_SLICE_X13Y120_CO6),
.Q(CLBLM_L_X10Y120_SLICE_X13Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffeffff)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_DLUT (
.I0(CLBLM_L_X10Y122_SLICE_X13Y122_AQ),
.I1(CLBLM_R_X5Y119_SLICE_X6Y119_CQ),
.I2(CLBLM_R_X7Y118_SLICE_X8Y118_DQ),
.I3(CLBLM_L_X8Y117_SLICE_X10Y117_BQ),
.I4(CLBLM_L_X10Y120_SLICE_X13Y120_BO5),
.I5(CLBLM_L_X10Y124_SLICE_X13Y124_AQ),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_DO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ff00cc00)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y121_SLICE_X13Y121_AQ),
.I2(CLBLM_R_X7Y125_SLICE_X9Y125_B5Q),
.I3(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I4(CLBLM_L_X10Y120_SLICE_X13Y120_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_CO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafc0003030303)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_BLUT (
.I0(CLBLM_L_X10Y121_SLICE_X12Y121_BQ),
.I1(CLBLM_L_X10Y120_SLICE_X13Y120_BQ),
.I2(CLBLM_L_X10Y119_SLICE_X13Y119_BQ),
.I3(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_BO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0ff00aaaa)
  ) CLBLM_L_X10Y120_SLICE_X13Y120_ALUT (
.I0(CLBLM_R_X7Y125_SLICE_X9Y125_B5Q),
.I1(CLBLM_L_X10Y121_SLICE_X13Y121_AQ),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y120_SLICE_X13Y120_AO5),
.O6(CLBLM_L_X10Y120_SLICE_X13Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y121_SLICE_X12Y121_CO5),
.Q(CLBLM_L_X10Y121_SLICE_X12Y121_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y121_SLICE_X12Y121_AO6),
.Q(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y121_SLICE_X12Y121_BO6),
.Q(CLBLM_L_X10Y121_SLICE_X12Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y121_SLICE_X12Y121_CO6),
.Q(CLBLM_L_X10Y121_SLICE_X12Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y121_SLICE_X12Y121_DO6),
.Q(CLBLM_L_X10Y121_SLICE_X12Y121_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0afa0afa0)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_DLUT (
.I0(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y123_SLICE_X5Y123_BQ),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y121_SLICE_X12Y121_DO5),
.O6(CLBLM_L_X10Y121_SLICE_X12Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3c0f3c0bbbb8888)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_CLUT (
.I0(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I3(CLBLM_L_X10Y126_SLICE_X12Y126_A5Q),
.I4(CLBLM_R_X11Y127_SLICE_X14Y127_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y121_SLICE_X12Y121_CO5),
.O6(CLBLM_L_X10Y121_SLICE_X12Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaacfc0aaaa0f00)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_BLUT (
.I0(CLBLL_L_X4Y121_SLICE_X4Y121_DQ),
.I1(CLBLM_L_X10Y121_SLICE_X12Y121_BQ),
.I2(CLBLM_L_X8Y123_SLICE_X10Y123_DO6),
.I3(CLBLM_R_X11Y121_SLICE_X14Y121_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y121_SLICE_X12Y121_BO5),
.O6(CLBLM_L_X10Y121_SLICE_X12Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfafaccccfa00)
  ) CLBLM_L_X10Y121_SLICE_X12Y121_ALUT (
.I0(CLBLM_L_X8Y121_SLICE_X11Y121_DO6),
.I1(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.I2(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.O5(CLBLM_L_X10Y121_SLICE_X12Y121_AO5),
.O6(CLBLM_L_X10Y121_SLICE_X12Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y121_SLICE_X13Y121_BO5),
.Q(CLBLM_L_X10Y121_SLICE_X13Y121_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y121_SLICE_X13Y121_AO6),
.Q(CLBLM_L_X10Y121_SLICE_X13Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y121_SLICE_X13Y121_BO6),
.Q(CLBLM_L_X10Y121_SLICE_X13Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y121_SLICE_X13Y121_CO6),
.Q(CLBLM_L_X10Y121_SLICE_X13Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdffddffdeffeeffe)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_DLUT (
.I0(CLBLM_R_X11Y123_SLICE_X14Y123_AQ),
.I1(CLBLM_L_X8Y120_SLICE_X10Y120_DO6),
.I2(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.I3(CLBLM_R_X11Y122_SLICE_X15Y122_BQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y121_SLICE_X14Y121_CQ),
.O5(CLBLM_L_X10Y121_SLICE_X13Y121_DO5),
.O6(CLBLM_L_X10Y121_SLICE_X13Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fcfcff00a8a8)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_CLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X10Y121_SLICE_X13Y121_CQ),
.I2(CLBLM_R_X5Y120_SLICE_X7Y120_DO6),
.I3(CLBLL_L_X4Y119_SLICE_X4Y119_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.O5(CLBLM_L_X10Y121_SLICE_X13Y121_CO5),
.O6(CLBLM_L_X10Y121_SLICE_X13Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa00aaf0ccf0cc)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(CLBLM_L_X8Y122_SLICE_X11Y122_A5Q),
.I2(CLBLM_R_X7Y117_SLICE_X8Y117_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y123_SLICE_X14Y123_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y121_SLICE_X13Y121_BO5),
.O6(CLBLM_L_X10Y121_SLICE_X13Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haafcaafcaa00aa00)
  ) CLBLM_L_X10Y121_SLICE_X13Y121_ALUT (
.I0(CLBLM_L_X8Y125_SLICE_X10Y125_CQ),
.I1(CLBLM_L_X10Y124_SLICE_X13Y124_AQ),
.I2(CLBLM_L_X10Y121_SLICE_X13Y121_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X3Y125_SLICE_X2Y125_BO6),
.O5(CLBLM_L_X10Y121_SLICE_X13Y121_AO5),
.O6(CLBLM_L_X10Y121_SLICE_X13Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X12Y122_AO6),
.Q(CLBLM_L_X10Y122_SLICE_X12Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X12Y122_BO6),
.Q(CLBLM_L_X10Y122_SLICE_X12Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffefefefe)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_DLUT (
.I0(CLBLL_L_X4Y122_SLICE_X5Y122_DQ),
.I1(CLBLM_L_X10Y123_SLICE_X12Y123_CQ),
.I2(CLBLM_R_X11Y123_SLICE_X14Y123_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_CQ),
.O5(CLBLM_L_X10Y122_SLICE_X12Y122_DO5),
.O6(CLBLM_L_X10Y122_SLICE_X12Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00f0ff0f03c3c)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y122_SLICE_X12Y122_AQ),
.I2(CLBLM_L_X10Y122_SLICE_X12Y122_BQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y126_SLICE_X13Y126_DQ),
.I5(CLBLM_L_X8Y122_SLICE_X10Y122_BO6),
.O5(CLBLM_L_X10Y122_SLICE_X12Y122_CO5),
.O6(CLBLM_L_X10Y122_SLICE_X12Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf303f303f000f000)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y124_SLICE_X13Y124_D5Q),
.I4(1'b1),
.I5(CLBLM_L_X10Y123_SLICE_X12Y123_CQ),
.O5(CLBLM_L_X10Y122_SLICE_X12Y122_BO5),
.O6(CLBLM_L_X10Y122_SLICE_X12Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc005acccc05a0)
  ) CLBLM_L_X10Y122_SLICE_X12Y122_ALUT (
.I0(CLBLM_L_X10Y123_SLICE_X12Y123_CQ),
.I1(CLBLM_L_X8Y123_SLICE_X11Y123_C5Q),
.I2(CLBLM_L_X10Y122_SLICE_X12Y122_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y122_SLICE_X12Y122_CO6),
.O5(CLBLM_L_X10Y122_SLICE_X12Y122_AO5),
.O6(CLBLM_L_X10Y122_SLICE_X12Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X13Y122_CO5),
.Q(CLBLM_L_X10Y122_SLICE_X13Y122_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X13Y122_AO6),
.Q(CLBLM_L_X10Y122_SLICE_X13Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X13Y122_CO6),
.Q(CLBLM_L_X10Y122_SLICE_X13Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y122_SLICE_X13Y122_DO6),
.Q(CLBLM_L_X10Y122_SLICE_X13Y122_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00ff55aa00)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_B5Q),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y122_SLICE_X13Y122_DO5),
.O6(CLBLM_L_X10Y122_SLICE_X13Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf505f000f4f40404)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLL_L_X4Y122_SLICE_X4Y122_DQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y123_SLICE_X13Y123_BQ),
.I4(CLBLM_L_X10Y122_SLICE_X12Y122_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y122_SLICE_X13Y122_CO5),
.O6(CLBLM_L_X10Y122_SLICE_X13Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcac0c0ffaa0000)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_BLUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_B5Q),
.I1(CLBLM_L_X10Y119_SLICE_X12Y119_DQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y121_SLICE_X13Y121_CQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y122_SLICE_X13Y122_BO5),
.O6(CLBLM_L_X10Y122_SLICE_X13Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaccc0aaaaccc0)
  ) CLBLM_L_X10Y122_SLICE_X13Y122_ALUT (
.I0(CLBLM_L_X10Y128_SLICE_X12Y128_CQ),
.I1(CLBLM_R_X3Y125_SLICE_X2Y125_BO6),
.I2(CLBLM_L_X10Y122_SLICE_X13Y122_AQ),
.I3(CLBLM_L_X10Y120_SLICE_X13Y120_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y122_SLICE_X13Y122_AO5),
.O6(CLBLM_L_X10Y122_SLICE_X13Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X12Y123_AO6),
.Q(CLBLM_L_X10Y123_SLICE_X12Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X12Y123_BO6),
.Q(CLBLM_L_X10Y123_SLICE_X12Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X12Y123_CO6),
.Q(CLBLM_L_X10Y123_SLICE_X12Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcf80c08cc88cc88)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_DLUT (
.I0(CLBLM_L_X10Y121_SLICE_X12Y121_AQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y122_SLICE_X13Y122_CQ),
.I4(CLBLM_R_X3Y125_SLICE_X2Y125_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_DO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacacaca0a0a0a0)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_CLUT (
.I0(CLBLM_R_X7Y119_SLICE_X9Y119_BQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y119_SLICE_X12Y119_BQ),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_CO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff4fe000f040e)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_BLUT (
.I0(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I1(CLBLM_L_X10Y123_SLICE_X12Y123_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y123_SLICE_X9Y123_DO6),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X10Y123_SLICE_X13Y123_CQ),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_BO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccaaccf0ccf0)
  ) CLBLM_L_X10Y123_SLICE_X12Y123_ALUT (
.I0(CLBLM_L_X8Y127_SLICE_X10Y127_CQ),
.I1(CLBLM_R_X11Y121_SLICE_X14Y121_CQ),
.I2(CLBLM_L_X10Y123_SLICE_X12Y123_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X10Y129_SLICE_X13Y129_DO6),
.O5(CLBLM_L_X10Y123_SLICE_X12Y123_AO5),
.O6(CLBLM_L_X10Y123_SLICE_X12Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X13Y123_AO6),
.Q(CLBLM_L_X10Y123_SLICE_X13Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X13Y123_BO6),
.Q(CLBLM_L_X10Y123_SLICE_X13Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X13Y123_CO6),
.Q(CLBLM_L_X10Y123_SLICE_X13Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00cc00fa00fa)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_DLUT (
.I0(CLBLM_L_X8Y118_SLICE_X10Y118_AQ),
.I1(CLBLM_L_X10Y123_SLICE_X13Y123_CQ),
.I2(CLBLL_L_X4Y121_SLICE_X5Y121_CQ),
.I3(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.I4(CLBLL_L_X4Y117_SLICE_X4Y117_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_DO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffc8ff00ffc8)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_CLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X10Y123_SLICE_X13Y123_CQ),
.I2(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I3(CLBLM_R_X7Y121_SLICE_X9Y121_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y126_SLICE_X14Y126_BQ),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_CO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000ccccf5f5)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_BLUT (
.I0(RIOB33_X105Y141_IOB_X1Y142_I),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y119_SLICE_X13Y119_CO6),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_BO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33fe32cc00dc10)
  ) CLBLM_L_X10Y123_SLICE_X13Y123_ALUT (
.I0(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y123_SLICE_X13Y123_AQ),
.I3(CLBLM_L_X10Y121_SLICE_X13Y121_CQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X10Y126_SLICE_X13Y126_CQ),
.O5(CLBLM_L_X10Y123_SLICE_X13Y123_AO5),
.O6(CLBLM_L_X10Y123_SLICE_X13Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X10Y121_SLICE_X13Y121_BQ),
.Q(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.R(CLBLM_L_X8Y131_SLICE_X11Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000aaaaaaaa)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_DLUT (
.I0(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y124_SLICE_X10Y124_AQ),
.O5(CLBLM_L_X10Y124_SLICE_X12Y124_DO5),
.O6(CLBLM_L_X10Y124_SLICE_X12Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf000002222)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_CLUT (
.I0(CLBLM_L_X8Y126_SLICE_X11Y126_CQ),
.I1(CLBLM_L_X10Y125_SLICE_X12Y125_BQ),
.I2(CLBLM_L_X10Y124_SLICE_X13Y124_B5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y124_SLICE_X13Y124_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y124_SLICE_X12Y124_CO5),
.O6(CLBLM_L_X10Y124_SLICE_X12Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00c8c837373737)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_BLUT (
.I0(CLBLM_R_X11Y124_SLICE_X14Y124_CQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLL_L_X4Y123_SLICE_X5Y123_BQ),
.I3(CLBLM_R_X11Y122_SLICE_X15Y122_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y124_SLICE_X12Y124_BO5),
.O6(CLBLM_L_X10Y124_SLICE_X12Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00bebe0c0c0c0c)
  ) CLBLM_L_X10Y124_SLICE_X12Y124_ALUT (
.I0(CLBLM_L_X10Y128_SLICE_X13Y128_CO6),
.I1(CLBLM_L_X8Y126_SLICE_X11Y126_CQ),
.I2(CLBLM_L_X10Y124_SLICE_X13Y124_C5Q),
.I3(CLBLM_L_X8Y121_SLICE_X11Y121_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y124_SLICE_X12Y124_AO5),
.O6(CLBLM_L_X10Y124_SLICE_X12Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y123_SLICE_X12Y123_DO6),
.Q(CLBLM_L_X10Y124_SLICE_X13Y124_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X12Y124_BO6),
.Q(CLBLM_L_X10Y124_SLICE_X13Y124_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X12Y124_AO6),
.Q(CLBLM_L_X10Y124_SLICE_X13Y124_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X12Y124_CO6),
.Q(CLBLM_L_X10Y124_SLICE_X13Y124_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X13Y124_AO6),
.Q(CLBLM_L_X10Y124_SLICE_X13Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X13Y124_BO6),
.Q(CLBLM_L_X10Y124_SLICE_X13Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X13Y124_CO6),
.Q(CLBLM_L_X10Y124_SLICE_X13Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y124_SLICE_X13Y124_DO6),
.Q(CLBLM_L_X10Y124_SLICE_X13Y124_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000030c030c)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y125_SLICE_X10Y125_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y122_SLICE_X13Y122_BO5),
.I4(CLBLM_L_X10Y124_SLICE_X13Y124_B5Q),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y124_SLICE_X13Y124_DO5),
.O6(CLBLM_L_X10Y124_SLICE_X13Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa003000cc)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_CLUT (
.I0(CLBLM_R_X11Y119_SLICE_X14Y119_BQ),
.I1(CLBLM_L_X10Y124_SLICE_X13Y124_CQ),
.I2(CLBLM_L_X10Y125_SLICE_X13Y125_CQ),
.I3(CLBLM_L_X10Y128_SLICE_X13Y128_CO6),
.I4(CLBLM_L_X10Y124_SLICE_X12Y124_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y124_SLICE_X13Y124_CO5),
.O6(CLBLM_L_X10Y124_SLICE_X13Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacafa0a0a0afa0)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_BLUT (
.I0(CLBLM_R_X7Y129_SLICE_X9Y129_AQ),
.I1(CLBLM_L_X10Y124_SLICE_X13Y124_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.I4(CLBLM_L_X8Y123_SLICE_X10Y123_DO6),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y124_SLICE_X13Y124_BO5),
.O6(CLBLM_L_X10Y124_SLICE_X13Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaac0aaccaac0)
  ) CLBLM_L_X10Y124_SLICE_X13Y124_ALUT (
.I0(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I1(CLBLM_R_X3Y125_SLICE_X2Y125_BO6),
.I2(CLBLM_L_X10Y124_SLICE_X13Y124_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y122_SLICE_X13Y122_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y124_SLICE_X13Y124_AO5),
.O6(CLBLM_L_X10Y124_SLICE_X13Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y125_SLICE_X12Y125_AO6),
.Q(CLBLM_L_X10Y125_SLICE_X12Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y125_SLICE_X12Y125_BO6),
.Q(CLBLM_L_X10Y125_SLICE_X12Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y125_SLICE_X12Y125_CO6),
.Q(CLBLM_L_X10Y125_SLICE_X12Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y125_SLICE_X12Y125_DO6),
.Q(CLBLM_L_X10Y125_SLICE_X12Y125_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55fa50ee44ea40)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X10Y125_SLICE_X12Y125_DQ),
.I3(CLBLM_L_X10Y124_SLICE_X13Y124_AQ),
.I4(CLBLM_L_X8Y125_SLICE_X11Y125_DO6),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.O5(CLBLM_L_X10Y125_SLICE_X12Y125_DO5),
.O6(CLBLM_L_X10Y125_SLICE_X12Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc05500550)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X11Y129_SLICE_X14Y129_BQ),
.I2(CLBLM_L_X8Y127_SLICE_X10Y127_CQ),
.I3(CLBLM_L_X10Y123_SLICE_X12Y123_DO5),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y125_SLICE_X12Y125_CO5),
.O6(CLBLM_L_X10Y125_SLICE_X12Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff1400000014)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_BLUT (
.I0(CLBLM_L_X10Y128_SLICE_X13Y128_CO6),
.I1(CLBLM_L_X10Y125_SLICE_X12Y125_BQ),
.I2(CLBLM_L_X10Y124_SLICE_X12Y124_AO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y125_SLICE_X13Y125_DO5),
.I5(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.O5(CLBLM_L_X10Y125_SLICE_X12Y125_BO5),
.O6(CLBLM_L_X10Y125_SLICE_X12Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff003232ff000000)
  ) CLBLM_L_X10Y125_SLICE_X12Y125_ALUT (
.I0(CLBLM_L_X8Y121_SLICE_X11Y121_DO6),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X10Y125_SLICE_X12Y125_AQ),
.I3(CLBLM_R_X7Y125_SLICE_X9Y125_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.O5(CLBLM_L_X10Y125_SLICE_X12Y125_AO5),
.O6(CLBLM_L_X10Y125_SLICE_X12Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y125_SLICE_X13Y125_AO6),
.Q(CLBLM_L_X10Y125_SLICE_X13Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y125_SLICE_X13Y125_BO6),
.Q(CLBLM_L_X10Y125_SLICE_X13Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y125_SLICE_X13Y125_CO6),
.Q(CLBLM_L_X10Y125_SLICE_X13Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000a00000002)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_DLUT (
.I0(CLBLM_L_X8Y126_SLICE_X11Y126_CQ),
.I1(CLBLM_L_X10Y125_SLICE_X13Y125_CQ),
.I2(CLBLM_L_X10Y125_SLICE_X12Y125_BQ),
.I3(CLBLM_L_X10Y124_SLICE_X13Y124_CQ),
.I4(CLBLM_L_X10Y124_SLICE_X13Y124_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y125_SLICE_X13Y125_DO5),
.O6(CLBLM_L_X10Y125_SLICE_X13Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfb51fe54fb51fe54)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y125_SLICE_X13Y125_CQ),
.I2(CLBLM_L_X10Y128_SLICE_X13Y128_CO6),
.I3(CLBLL_L_X4Y120_SLICE_X4Y120_DQ),
.I4(CLBLM_L_X10Y125_SLICE_X13Y125_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y125_SLICE_X13Y125_CO5),
.O6(CLBLM_L_X10Y125_SLICE_X13Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f05555f0f04444)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_BLUT (
.I0(CLBLM_L_X10Y129_SLICE_X13Y129_DO6),
.I1(CLBLM_L_X10Y125_SLICE_X13Y125_BQ),
.I2(CLBLM_L_X10Y125_SLICE_X13Y125_CQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y125_SLICE_X10Y125_CQ),
.O5(CLBLM_L_X10Y125_SLICE_X13Y125_BO5),
.O6(CLBLM_L_X10Y125_SLICE_X13Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50aa00fe54aa00)
  ) CLBLM_L_X10Y125_SLICE_X13Y125_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.I2(CLBLM_L_X10Y125_SLICE_X13Y125_AQ),
.I3(CLBLM_L_X8Y117_SLICE_X10Y117_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_L_X10Y125_SLICE_X13Y125_AO5),
.O6(CLBLM_L_X10Y125_SLICE_X13Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y126_SLICE_X12Y126_BO6),
.Q(CLBLM_L_X10Y126_SLICE_X12Y126_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y126_SLICE_X12Y126_AO6),
.Q(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y126_SLICE_X12Y126_CO6),
.Q(CLBLM_L_X10Y126_SLICE_X12Y126_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00fc00fc00ff00aa)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_DLUT (
.I0(CLBLM_L_X10Y125_SLICE_X12Y125_AQ),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_AQ),
.I2(CLBLM_L_X8Y126_SLICE_X11Y126_DQ),
.I3(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.I4(CLBLM_L_X10Y120_SLICE_X12Y120_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y126_SLICE_X12Y126_DO5),
.O6(CLBLM_L_X10Y126_SLICE_X12Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f08888f0f08888)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X11Y123_SLICE_X14Y123_DQ),
.I2(CLBLM_L_X8Y126_SLICE_X11Y126_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y126_SLICE_X12Y126_CO5),
.O6(CLBLM_L_X10Y126_SLICE_X12Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbb88888fff00000)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_BLUT (
.I0(CLBLM_L_X10Y126_SLICE_X13Y126_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y125_SLICE_X11Y125_CQ),
.I3(CLBLL_L_X4Y122_SLICE_X5Y122_DQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y126_SLICE_X12Y126_BO5),
.O6(CLBLM_L_X10Y126_SLICE_X12Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff220022ffe200e2)
  ) CLBLM_L_X10Y126_SLICE_X12Y126_ALUT (
.I0(CLBLM_L_X10Y128_SLICE_X12Y128_CQ),
.I1(CLBLM_R_X11Y126_SLICE_X15Y126_DO5),
.I2(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y125_SLICE_X12Y125_AQ),
.I5(CLBLM_L_X10Y128_SLICE_X13Y128_CO6),
.O5(CLBLM_L_X10Y126_SLICE_X12Y126_AO5),
.O6(CLBLM_L_X10Y126_SLICE_X12Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y126_SLICE_X13Y126_AO6),
.Q(CLBLM_L_X10Y126_SLICE_X13Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y126_SLICE_X13Y126_BO6),
.Q(CLBLM_L_X10Y126_SLICE_X13Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y126_SLICE_X13Y126_CO6),
.Q(CLBLM_L_X10Y126_SLICE_X13Y126_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y126_SLICE_X13Y126_DO6),
.Q(CLBLM_L_X10Y126_SLICE_X13Y126_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f055550000)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(CLBLM_L_X12Y127_SLICE_X16Y127_AQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y122_SLICE_X5Y122_DQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y126_SLICE_X13Y126_DO5),
.O6(CLBLM_L_X10Y126_SLICE_X13Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fe000ef0f00000)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_CLUT (
.I0(CLBLM_L_X10Y123_SLICE_X13Y123_BQ),
.I1(CLBLM_L_X10Y126_SLICE_X13Y126_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X10Y126_SLICE_X13Y126_AQ),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.O5(CLBLM_L_X10Y126_SLICE_X13Y126_CO5),
.O6(CLBLM_L_X10Y126_SLICE_X13Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf044f0fff044f000)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_BLUT (
.I0(CLBLM_L_X10Y128_SLICE_X13Y128_CO6),
.I1(CLBLM_L_X10Y126_SLICE_X13Y126_BQ),
.I2(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y126_SLICE_X15Y126_DO5),
.I5(CLBLM_R_X11Y126_SLICE_X14Y126_DQ),
.O5(CLBLM_L_X10Y126_SLICE_X13Y126_BO5),
.O6(CLBLM_L_X10Y126_SLICE_X13Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88bb8888b8bbb888)
  ) CLBLM_L_X10Y126_SLICE_X13Y126_ALUT (
.I0(CLBLM_R_X3Y119_SLICE_X2Y119_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y126_SLICE_X13Y126_AQ),
.I3(CLBLM_R_X11Y126_SLICE_X15Y126_DO5),
.I4(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.I5(CLBLM_L_X10Y128_SLICE_X13Y128_CO6),
.O5(CLBLM_L_X10Y126_SLICE_X13Y126_AO5),
.O6(CLBLM_L_X10Y126_SLICE_X13Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X12Y127_AO6),
.Q(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X12Y127_BO6),
.Q(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X12Y127_CO6),
.Q(CLBLM_L_X10Y127_SLICE_X12Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X12Y127_DO6),
.Q(CLBLM_L_X10Y127_SLICE_X12Y127_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcacfcfcfcfcfcf)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_DLUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(CLBLM_L_X10Y126_SLICE_X12Y126_A5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y129_SLICE_X12Y129_CO6),
.I4(RIOB33_X105Y135_IOB_X1Y135_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_L_X10Y127_SLICE_X12Y127_DO5),
.O6(CLBLM_L_X10Y127_SLICE_X12Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0d1d1c0c0d1d1c0)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.I3(CLBLM_L_X10Y126_SLICE_X12Y126_BO5),
.I4(CLBLL_L_X4Y125_SLICE_X4Y125_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y127_SLICE_X12Y127_CO5),
.O6(CLBLM_L_X10Y127_SLICE_X12Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5e4e4f5f5e4e4)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y126_SLICE_X11Y126_CQ),
.I2(CLBLM_R_X3Y121_SLICE_X2Y121_CQ),
.I3(1'b1),
.I4(CLBLM_R_X11Y127_SLICE_X15Y127_BO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y127_SLICE_X12Y127_BO5),
.O6(CLBLM_L_X10Y127_SLICE_X12Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55fe54aa00ba10)
  ) CLBLM_L_X10Y127_SLICE_X12Y127_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X10Y127_SLICE_X12Y127_AQ),
.I3(CLBLM_L_X10Y127_SLICE_X13Y127_BQ),
.I4(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I5(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.O5(CLBLM_L_X10Y127_SLICE_X12Y127_AO5),
.O6(CLBLM_L_X10Y127_SLICE_X12Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X13Y127_AO6),
.Q(CLBLM_L_X10Y127_SLICE_X13Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X13Y127_BO6),
.Q(CLBLM_L_X10Y127_SLICE_X13Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X13Y127_CO6),
.Q(CLBLM_L_X10Y127_SLICE_X13Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y127_SLICE_X13Y127_DO6),
.Q(CLBLM_L_X10Y127_SLICE_X13Y127_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0055550000)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_DLUT (
.I0(CLBLM_R_X11Y127_SLICE_X15Y127_BO6),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X4Y125_SLICE_X4Y125_CQ),
.I4(CLBLM_L_X10Y127_SLICE_X13Y127_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y127_SLICE_X13Y127_DO5),
.O6(CLBLM_L_X10Y127_SLICE_X13Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aafeff000000)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_CLUT (
.I0(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.I1(CLBLM_R_X11Y128_SLICE_X15Y128_AQ),
.I2(CLBLM_L_X10Y128_SLICE_X12Y128_AQ),
.I3(CLBLM_R_X11Y126_SLICE_X15Y126_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y127_SLICE_X12Y127_BQ),
.O5(CLBLM_L_X10Y127_SLICE_X13Y127_CO5),
.O6(CLBLM_L_X10Y127_SLICE_X13Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00fa50ee44fa50)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y127_SLICE_X13Y127_BQ),
.I2(CLBLM_R_X11Y126_SLICE_X15Y126_CQ),
.I3(CLBLM_L_X8Y128_SLICE_X11Y128_AQ),
.I4(CLBLM_R_X11Y126_SLICE_X15Y126_DO5),
.I5(CLBLM_L_X10Y128_SLICE_X13Y128_CO6),
.O5(CLBLM_L_X10Y127_SLICE_X13Y127_BO5),
.O6(CLBLM_L_X10Y127_SLICE_X13Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaffaaffaa3f)
  ) CLBLM_L_X10Y127_SLICE_X13Y127_ALUT (
.I0(CLBLM_L_X10Y127_SLICE_X13Y127_CQ),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y135_IOB_X1Y135_I),
.I5(CLBLM_L_X10Y129_SLICE_X12Y129_CO6),
.O5(CLBLM_L_X10Y127_SLICE_X13Y127_AO5),
.O6(CLBLM_L_X10Y127_SLICE_X13Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y128_SLICE_X12Y128_AO6),
.Q(CLBLM_L_X10Y128_SLICE_X12Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y128_SLICE_X12Y128_BO6),
.Q(CLBLM_L_X10Y128_SLICE_X12Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y128_SLICE_X12Y128_CO6),
.Q(CLBLM_L_X10Y128_SLICE_X12Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y128_SLICE_X12Y128_DO6),
.Q(CLBLM_L_X10Y128_SLICE_X12Y128_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff44ff4500440045)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_DLUT (
.I0(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.I1(CLBLM_R_X11Y126_SLICE_X15Y126_BQ),
.I2(CLBLM_L_X10Y128_SLICE_X12Y128_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y128_SLICE_X15Y128_AQ),
.I5(CLBLM_L_X8Y129_SLICE_X11Y129_BQ),
.O5(CLBLM_L_X10Y128_SLICE_X12Y128_DO5),
.O6(CLBLM_L_X10Y128_SLICE_X12Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haafaeefa00504450)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y128_SLICE_X12Y128_CQ),
.I2(CLBLM_L_X10Y126_SLICE_X13Y126_BQ),
.I3(CLBLM_R_X11Y126_SLICE_X15Y126_DO5),
.I4(CLBLM_L_X10Y128_SLICE_X13Y128_CO6),
.I5(CLBLM_R_X7Y126_SLICE_X8Y126_CQ),
.O5(CLBLM_L_X10Y128_SLICE_X12Y128_CO5),
.O6(CLBLM_L_X10Y128_SLICE_X12Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaaf0f0ffee)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_BLUT (
.I0(CLBLM_L_X10Y128_SLICE_X13Y128_CO6),
.I1(CLBLM_L_X10Y128_SLICE_X12Y128_BQ),
.I2(CLBLM_L_X8Y128_SLICE_X10Y128_CQ),
.I3(CLBLM_L_X10Y127_SLICE_X13Y127_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y126_SLICE_X15Y126_DO5),
.O5(CLBLM_L_X10Y128_SLICE_X12Y128_BO5),
.O6(CLBLM_L_X10Y128_SLICE_X12Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddcc1100dcdc1010)
  ) CLBLM_L_X10Y128_SLICE_X12Y128_ALUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y128_SLICE_X12Y128_AQ),
.I3(CLBLM_R_X11Y128_SLICE_X15Y128_AQ),
.I4(CLBLM_R_X5Y127_SLICE_X7Y127_B5Q),
.I5(CLBLM_R_X11Y127_SLICE_X15Y127_CO5),
.O5(CLBLM_L_X10Y128_SLICE_X12Y128_AO5),
.O6(CLBLM_L_X10Y128_SLICE_X12Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y128_SLICE_X13Y128_AO6),
.Q(CLBLM_L_X10Y128_SLICE_X13Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y128_SLICE_X13Y128_BO6),
.Q(CLBLM_L_X10Y128_SLICE_X13Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033000300320032)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_DLUT (
.I0(CLBLM_L_X10Y128_SLICE_X13Y128_CO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y127_SLICE_X13Y127_BQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X11Y126_SLICE_X15Y126_DO5),
.I5(CLBLM_L_X8Y129_SLICE_X11Y129_BQ),
.O5(CLBLM_L_X10Y128_SLICE_X13Y128_DO5),
.O6(CLBLM_L_X10Y128_SLICE_X13Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000500000400)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_CLUT (
.I0(CLBLM_R_X11Y128_SLICE_X15Y128_AQ),
.I1(CLBLM_L_X10Y125_SLICE_X13Y125_DO5),
.I2(CLBLM_L_X10Y128_SLICE_X12Y128_AQ),
.I3(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.I4(CLBLM_R_X11Y126_SLICE_X15Y126_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y128_SLICE_X13Y128_CO5),
.O6(CLBLM_L_X10Y128_SLICE_X13Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff005050ff00d8d8)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_BLUT (
.I0(CLBLM_R_X11Y126_SLICE_X15Y126_DO5),
.I1(CLBLM_L_X10Y128_SLICE_X13Y128_BQ),
.I2(CLBLM_L_X10Y126_SLICE_X13Y126_AQ),
.I3(CLBLM_R_X7Y125_SLICE_X8Y125_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y128_SLICE_X13Y128_CO6),
.O5(CLBLM_L_X10Y128_SLICE_X13Y128_BO5),
.O6(CLBLM_L_X10Y128_SLICE_X13Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0afa0a0a0afa0)
  ) CLBLM_L_X10Y128_SLICE_X13Y128_ALUT (
.I0(CLBLM_L_X8Y128_SLICE_X11Y128_DQ),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y128_SLICE_X14Y128_BO6),
.I4(CLBLM_R_X11Y127_SLICE_X15Y127_BO5),
.I5(1'b1),
.O5(CLBLM_L_X10Y128_SLICE_X13Y128_AO5),
.O6(CLBLM_L_X10Y128_SLICE_X13Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y124_SLICE_X11Y124_CO6),
.Q(CLBLM_L_X10Y129_SLICE_X12Y129_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y129_SLICE_X12Y129_AO6),
.Q(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y129_SLICE_X12Y129_BO6),
.Q(CLBLM_L_X10Y129_SLICE_X12Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y129_SLICE_X12Y129_DO5),
.O6(CLBLM_L_X10Y129_SLICE_X12Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_CLUT (
.I0(RIOB33_X105Y129_IOB_X1Y130_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y127_IOB_X1Y128_I),
.I5(RIOB33_X105Y133_IOB_X1Y134_I),
.O5(CLBLM_L_X10Y129_SLICE_X12Y129_CO5),
.O6(CLBLM_L_X10Y129_SLICE_X12Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffd0f0f0f0d)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_BLUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(CLBLM_L_X10Y129_SLICE_X12Y129_CO6),
.I5(CLBLM_L_X10Y129_SLICE_X12Y129_A5Q),
.O5(CLBLM_L_X10Y129_SLICE_X12Y129_BO5),
.O6(CLBLM_L_X10Y129_SLICE_X12Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888d8d88dd8)
  ) CLBLM_L_X10Y129_SLICE_X12Y129_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y129_SLICE_X12Y129_BQ),
.I2(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.I3(CLBLM_R_X11Y127_SLICE_X15Y127_CO5),
.I4(CLBLM_L_X10Y129_SLICE_X13Y129_BO6),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_L_X10Y129_SLICE_X12Y129_AO5),
.O6(CLBLM_L_X10Y129_SLICE_X12Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y129_SLICE_X13Y129_AO6),
.Q(CLBLM_L_X10Y129_SLICE_X13Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0202ffff0202ffff)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_DLUT (
.I0(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X10Y125_SLICE_X13Y125_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y129_SLICE_X13Y129_DO5),
.O6(CLBLM_L_X10Y129_SLICE_X13Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000fffffffdffff)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_CLUT (
.I0(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.I1(CLBLM_R_X11Y126_SLICE_X15Y126_BQ),
.I2(CLBLM_L_X10Y128_SLICE_X12Y128_AQ),
.I3(CLBLM_R_X11Y128_SLICE_X15Y128_AQ),
.I4(CLBLM_L_X10Y125_SLICE_X13Y125_DO5),
.I5(CLBLM_L_X8Y129_SLICE_X11Y129_BQ),
.O5(CLBLM_L_X10Y129_SLICE_X13Y129_CO5),
.O6(CLBLM_L_X10Y129_SLICE_X13Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf453333ccccc0c0)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_BLUT (
.I0(CLBLM_R_X11Y126_SLICE_X15Y126_BQ),
.I1(CLBLM_L_X10Y128_SLICE_X12Y128_AQ),
.I2(CLBLM_R_X11Y128_SLICE_X15Y128_AQ),
.I3(CLBLM_L_X8Y129_SLICE_X11Y129_BQ),
.I4(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y129_SLICE_X13Y129_BO5),
.O6(CLBLM_L_X10Y129_SLICE_X13Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff555000005550)
  ) CLBLM_L_X10Y129_SLICE_X13Y129_ALUT (
.I0(CLBLM_L_X10Y129_SLICE_X13Y129_DO6),
.I1(1'b1),
.I2(CLBLM_L_X10Y129_SLICE_X13Y129_AQ),
.I3(CLBLM_L_X10Y124_SLICE_X13Y124_DQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y121_SLICE_X14Y121_BQ),
.O5(CLBLM_L_X10Y129_SLICE_X13Y129_AO5),
.O6(CLBLM_L_X10Y129_SLICE_X13Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X11Y128_SLICE_X15Y128_AQ),
.Q(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.R(CLBLM_L_X8Y131_SLICE_X11Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_DO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_CO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_BO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_AO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_DO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_CO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_BO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_AO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y136_SLICE_X12Y136_BO5),
.Q(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y136_SLICE_X12Y136_AO6),
.Q(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y135_SLICE_X12Y135_DO5),
.O6(CLBLM_L_X10Y135_SLICE_X12Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y135_SLICE_X12Y135_CO5),
.O6(CLBLM_L_X10Y135_SLICE_X12Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y135_SLICE_X12Y135_BO5),
.O6(CLBLM_L_X10Y135_SLICE_X12Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y135_SLICE_X12Y135_AO5),
.O6(CLBLM_L_X10Y135_SLICE_X12Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y135_SLICE_X13Y135_DO5),
.O6(CLBLM_L_X10Y135_SLICE_X13Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y135_SLICE_X13Y135_CO5),
.O6(CLBLM_L_X10Y135_SLICE_X13Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y135_SLICE_X13Y135_BO5),
.O6(CLBLM_L_X10Y135_SLICE_X13Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y135_SLICE_X13Y135_AO5),
.O6(CLBLM_L_X10Y135_SLICE_X13Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y136_SLICE_X12Y136_DO5),
.O6(CLBLM_L_X10Y136_SLICE_X12Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y136_SLICE_X12Y136_CO5),
.O6(CLBLM_L_X10Y136_SLICE_X12Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ff55ff00cccc)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_BLUT (
.I0(RIOB33_X105Y143_IOB_X1Y143_I),
.I1(CLBLM_L_X10Y129_SLICE_X12Y129_A5Q),
.I2(1'b1),
.I3(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y136_SLICE_X12Y136_BO5),
.O6(CLBLM_L_X10Y136_SLICE_X12Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0acc0accccffff)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_ALUT (
.I0(CLBLM_R_X7Y126_SLICE_X9Y126_DQ),
.I1(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y136_SLICE_X12Y136_AO5),
.O6(CLBLM_L_X10Y136_SLICE_X12Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y136_SLICE_X13Y136_DO5),
.O6(CLBLM_L_X10Y136_SLICE_X13Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y136_SLICE_X13Y136_CO5),
.O6(CLBLM_L_X10Y136_SLICE_X13Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y136_SLICE_X13Y136_BO5),
.O6(CLBLM_L_X10Y136_SLICE_X13Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y136_SLICE_X13Y136_AO5),
.O6(CLBLM_L_X10Y136_SLICE_X13Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y121_SLICE_X16Y121_AO6),
.Q(CLBLM_L_X12Y121_SLICE_X16Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y121_SLICE_X16Y121_BO6),
.Q(CLBLM_L_X12Y121_SLICE_X16Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y121_SLICE_X16Y121_DO5),
.O6(CLBLM_L_X12Y121_SLICE_X16Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y121_SLICE_X16Y121_CO5),
.O6(CLBLM_L_X12Y121_SLICE_X16Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hef45ef45ee44ee44)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y121_SLICE_X16Y121_BQ),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.I3(CLBLM_L_X10Y120_SLICE_X13Y120_A5Q),
.I4(1'b1),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_L_X12Y121_SLICE_X16Y121_BO5),
.O6(CLBLM_L_X12Y121_SLICE_X16Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d888dd888888dd)
  ) CLBLM_L_X12Y121_SLICE_X16Y121_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y121_SLICE_X16Y121_BQ),
.I2(CLBLM_L_X12Y121_SLICE_X16Y121_AQ),
.I3(CLBLM_R_X11Y121_SLICE_X15Y121_CO6),
.I4(CLBLM_L_X8Y123_SLICE_X10Y123_DO6),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X12Y121_SLICE_X16Y121_AO5),
.O6(CLBLM_L_X12Y121_SLICE_X16Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y121_SLICE_X17Y121_DO5),
.O6(CLBLM_L_X12Y121_SLICE_X17Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y121_SLICE_X17Y121_CO5),
.O6(CLBLM_L_X12Y121_SLICE_X17Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y121_SLICE_X17Y121_BO5),
.O6(CLBLM_L_X12Y121_SLICE_X17Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y121_SLICE_X17Y121_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y121_SLICE_X17Y121_AO5),
.O6(CLBLM_L_X12Y121_SLICE_X17Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y126_SLICE_X16Y126_AO6),
.Q(CLBLM_L_X12Y126_SLICE_X16Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y126_SLICE_X16Y126_BO6),
.Q(CLBLM_L_X12Y126_SLICE_X16Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y126_SLICE_X16Y126_DO5),
.O6(CLBLM_L_X12Y126_SLICE_X16Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y126_SLICE_X16Y126_CO5),
.O6(CLBLM_L_X12Y126_SLICE_X16Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0cfcfcac5)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_BLUT (
.I0(CLBLM_L_X12Y126_SLICE_X16Y126_BQ),
.I1(CLBLM_R_X7Y127_SLICE_X8Y127_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y127_SLICE_X16Y127_BO6),
.I4(CLBLM_R_X11Y130_SLICE_X14Y130_BO5),
.I5(CLBLM_R_X11Y127_SLICE_X15Y127_BO5),
.O5(CLBLM_L_X12Y126_SLICE_X16Y126_BO5),
.O6(CLBLM_L_X12Y126_SLICE_X16Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8bbb8b8b8bbb8b8)
  ) CLBLM_L_X12Y126_SLICE_X16Y126_ALUT (
.I0(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y126_SLICE_X16Y126_AQ),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.I4(RIOB33_X105Y141_IOB_X1Y142_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y126_SLICE_X16Y126_AO5),
.O6(CLBLM_L_X12Y126_SLICE_X16Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y126_SLICE_X17Y126_DO5),
.O6(CLBLM_L_X12Y126_SLICE_X17Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y126_SLICE_X17Y126_CO5),
.O6(CLBLM_L_X12Y126_SLICE_X17Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y126_SLICE_X17Y126_BO5),
.O6(CLBLM_L_X12Y126_SLICE_X17Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y126_SLICE_X17Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y126_SLICE_X17Y126_AO5),
.O6(CLBLM_L_X12Y126_SLICE_X17Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y127_SLICE_X16Y127_AO6),
.Q(CLBLM_L_X12Y127_SLICE_X16Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff6633ffff6666)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_DLUT (
.I0(CLBLM_L_X10Y129_SLICE_X13Y129_CO6),
.I1(CLBLM_L_X12Y127_SLICE_X16Y127_AQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y128_SLICE_X14Y128_AO5),
.I4(CLBLM_R_X11Y130_SLICE_X14Y130_BO5),
.I5(CLBLM_L_X10Y128_SLICE_X12Y128_BQ),
.O5(CLBLM_L_X12Y127_SLICE_X16Y127_DO5),
.O6(CLBLM_L_X12Y127_SLICE_X16Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000010000)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_CLUT (
.I0(CLBLM_L_X12Y126_SLICE_X16Y126_BQ),
.I1(CLBLM_R_X11Y126_SLICE_X15Y126_AQ),
.I2(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.I3(CLBLM_R_X11Y126_SLICE_X14Y126_CQ),
.I4(CLBLM_R_X11Y128_SLICE_X15Y128_DO6),
.I5(CLBLM_L_X10Y128_SLICE_X13Y128_AQ),
.O5(CLBLM_L_X12Y127_SLICE_X16Y127_CO5),
.O6(CLBLM_L_X12Y127_SLICE_X16Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000bbbf0000ffbf)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_BLUT (
.I0(CLBLM_R_X11Y128_SLICE_X14Y128_AO5),
.I1(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.I2(CLBLM_R_X11Y128_SLICE_X15Y128_DO6),
.I3(CLBLM_L_X10Y128_SLICE_X13Y128_AQ),
.I4(CLBLM_L_X10Y129_SLICE_X13Y129_CO6),
.I5(CLBLM_R_X11Y128_SLICE_X14Y128_DO6),
.O5(CLBLM_L_X12Y127_SLICE_X16Y127_BO5),
.O6(CLBLM_L_X12Y127_SLICE_X16Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0cacacaca)
  ) CLBLM_L_X12Y127_SLICE_X16Y127_ALUT (
.I0(CLBLM_L_X12Y127_SLICE_X16Y127_DO6),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X11Y127_SLICE_X15Y127_BO5),
.O5(CLBLM_L_X12Y127_SLICE_X16Y127_AO5),
.O6(CLBLM_L_X12Y127_SLICE_X16Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000022)
  ) CLBLM_L_X12Y127_SLICE_X17Y127_DLUT (
.I0(CLBLM_R_X11Y128_SLICE_X15Y128_DO6),
.I1(CLBLM_R_X11Y126_SLICE_X14Y126_CQ),
.I2(1'b1),
.I3(CLBLM_L_X12Y126_SLICE_X16Y126_BQ),
.I4(CLBLM_R_X11Y126_SLICE_X15Y126_AQ),
.I5(CLBLM_L_X10Y128_SLICE_X13Y128_AQ),
.O5(CLBLM_L_X12Y127_SLICE_X17Y127_DO5),
.O6(CLBLM_L_X12Y127_SLICE_X17Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff7fffffffffff)
  ) CLBLM_L_X12Y127_SLICE_X17Y127_CLUT (
.I0(CLBLM_L_X12Y126_SLICE_X16Y126_BQ),
.I1(CLBLM_R_X11Y126_SLICE_X14Y126_CQ),
.I2(CLBLM_R_X11Y126_SLICE_X15Y126_AQ),
.I3(CLBLM_R_X11Y128_SLICE_X14Y128_DO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y128_SLICE_X13Y128_AQ),
.O5(CLBLM_L_X12Y127_SLICE_X17Y127_CO5),
.O6(CLBLM_L_X12Y127_SLICE_X17Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X12Y127_SLICE_X17Y127_BLUT (
.I0(CLBLM_R_X11Y126_SLICE_X15Y126_AQ),
.I1(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.I2(CLBLM_L_X12Y126_SLICE_X16Y126_BQ),
.I3(CLBLM_L_X10Y128_SLICE_X13Y128_AQ),
.I4(CLBLM_R_X11Y128_SLICE_X14Y128_DO6),
.I5(CLBLM_R_X11Y126_SLICE_X14Y126_CQ),
.O5(CLBLM_L_X12Y127_SLICE_X17Y127_BO5),
.O6(CLBLM_L_X12Y127_SLICE_X17Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffdf2000ffcf30)
  ) CLBLM_L_X12Y127_SLICE_X17Y127_ALUT (
.I0(CLBLM_L_X12Y127_SLICE_X17Y127_DO6),
.I1(CLBLM_R_X11Y128_SLICE_X14Y128_AO5),
.I2(CLBLM_R_X11Y126_SLICE_X15Y126_CQ),
.I3(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.I4(CLBLM_L_X10Y129_SLICE_X13Y129_CO6),
.I5(CLBLM_L_X12Y127_SLICE_X17Y127_CO6),
.O5(CLBLM_L_X12Y127_SLICE_X17Y127_AO5),
.O6(CLBLM_L_X12Y127_SLICE_X17Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y118_SLICE_X2Y118_AO6),
.Q(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_DO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff7ffffffffffff)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_CLUT (
.I0(CLBLM_R_X3Y119_SLICE_X2Y119_AQ),
.I1(CLBLL_L_X2Y119_SLICE_X1Y119_AQ),
.I2(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I3(CLBLM_R_X7Y117_SLICE_X9Y117_DO6),
.I4(CLBLM_R_X3Y119_SLICE_X3Y119_BO5),
.I5(CLBLM_R_X3Y119_SLICE_X2Y119_BQ),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_CO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h80800000cc80cc00)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_BLUT (
.I0(CLBLL_L_X2Y119_SLICE_X1Y119_AQ),
.I1(CLBLM_R_X3Y119_SLICE_X2Y119_BQ),
.I2(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y119_SLICE_X2Y119_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_BO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccca0a000aa)
  ) CLBLM_R_X3Y118_SLICE_X2Y118_ALUT (
.I0(CLBLM_R_X3Y119_SLICE_X2Y119_CO6),
.I1(CLBLM_R_X5Y119_SLICE_X7Y119_CQ),
.I2(CLBLM_R_X3Y118_SLICE_X2Y118_AQ),
.I3(CLBLM_R_X3Y118_SLICE_X2Y118_BO6),
.I4(CLBLM_R_X3Y118_SLICE_X2Y118_CO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y118_SLICE_X2Y118_AO5),
.O6(CLBLM_R_X3Y118_SLICE_X2Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y118_SLICE_X3Y118_AO6),
.Q(CLBLM_R_X3Y118_SLICE_X3Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y118_SLICE_X3Y118_BO6),
.Q(CLBLM_R_X3Y118_SLICE_X3Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_DO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7ff77fff7ffffff)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_CLUT (
.I0(CLBLL_L_X4Y118_SLICE_X5Y118_BQ),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_BQ),
.I2(CLBLM_R_X3Y118_SLICE_X3Y118_BQ),
.I3(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I4(CLBLM_R_X3Y118_SLICE_X3Y118_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_CO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0040405050)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_BLUT (
.I0(CLBLM_L_X8Y123_SLICE_X11Y123_CQ),
.I1(CLBLM_R_X3Y118_SLICE_X3Y118_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I4(CLBLM_R_X3Y118_SLICE_X3Y118_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_BO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdc10cc00cd01cc00)
  ) CLBLM_R_X3Y118_SLICE_X3Y118_ALUT (
.I0(CLBLM_L_X8Y123_SLICE_X11Y123_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y118_SLICE_X3Y118_AQ),
.I3(CLBLL_L_X2Y125_SLICE_X1Y125_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X3Y118_SLICE_X3Y118_CO6),
.O5(CLBLM_R_X3Y118_SLICE_X3Y118_AO5),
.O6(CLBLM_R_X3Y118_SLICE_X3Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y119_SLICE_X2Y119_AO6),
.Q(CLBLM_R_X3Y119_SLICE_X2Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y119_SLICE_X2Y119_BO6),
.Q(CLBLM_R_X3Y119_SLICE_X2Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcfffcfffffffff)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y117_SLICE_X9Y117_DO6),
.I2(CLBLM_R_X3Y119_SLICE_X3Y119_BO5),
.I3(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I4(1'b1),
.I5(CLBLL_L_X2Y119_SLICE_X1Y119_AQ),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_DO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc44c400f000f0)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_CLUT (
.I0(CLBLM_L_X8Y123_SLICE_X11Y123_CQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLL_L_X2Y118_SLICE_X1Y118_B5Q),
.I3(CLBLL_L_X2Y118_SLICE_X1Y118_A5Q),
.I4(CLBLM_R_X5Y120_SLICE_X7Y120_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_CO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff009c9cff000000)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_BLUT (
.I0(CLBLM_R_X3Y119_SLICE_X2Y119_DO6),
.I1(CLBLM_R_X3Y119_SLICE_X2Y119_BQ),
.I2(CLBLM_R_X3Y119_SLICE_X2Y119_AQ),
.I3(CLBLM_L_X10Y119_SLICE_X12Y119_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X3Y119_SLICE_X2Y119_CO6),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_BO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hedfc2130cccc0000)
  ) CLBLM_R_X3Y119_SLICE_X2Y119_ALUT (
.I0(CLBLM_R_X3Y119_SLICE_X3Y119_CO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y119_SLICE_X2Y119_AQ),
.I3(CLBLL_L_X2Y119_SLICE_X1Y119_AQ),
.I4(CLBLL_L_X4Y119_SLICE_X4Y119_DQ),
.I5(CLBLM_R_X3Y119_SLICE_X2Y119_CO6),
.O5(CLBLM_R_X3Y119_SLICE_X2Y119_AO5),
.O6(CLBLM_R_X3Y119_SLICE_X2Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y119_SLICE_X3Y119_AO6),
.Q(CLBLM_R_X3Y119_SLICE_X3Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff3f5515ffff5555)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_DLUT (
.I0(CLBLL_L_X2Y127_SLICE_X0Y127_CO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X3Y123_SLICE_X3Y123_CQ),
.I3(CLBLL_L_X4Y120_SLICE_X4Y120_CQ),
.I4(CLBLM_L_X10Y120_SLICE_X12Y120_AQ),
.I5(CLBLM_R_X3Y128_SLICE_X3Y128_BO6),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_DO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdfffffffffffff)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_CLUT (
.I0(CLBLL_L_X4Y119_SLICE_X4Y119_BQ),
.I1(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I2(CLBLM_R_X3Y118_SLICE_X3Y118_AQ),
.I3(CLBLM_R_X7Y117_SLICE_X9Y117_DO6),
.I4(CLBLL_L_X4Y118_SLICE_X5Y118_BQ),
.I5(CLBLM_R_X3Y118_SLICE_X3Y118_BQ),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_CO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbf3f3f3fa0000000)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_BLUT (
.I0(CLBLM_R_X3Y118_SLICE_X3Y118_AQ),
.I1(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I2(CLBLL_L_X4Y118_SLICE_X5Y118_BQ),
.I3(CLBLM_R_X3Y118_SLICE_X3Y118_BQ),
.I4(CLBLL_L_X4Y119_SLICE_X4Y119_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_BO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00c0c0f0f0)
  ) CLBLM_R_X3Y119_SLICE_X3Y119_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I2(CLBLM_R_X3Y119_SLICE_X3Y119_AQ),
.I3(CLBLM_R_X3Y124_SLICE_X2Y124_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y119_SLICE_X3Y119_AO5),
.O6(CLBLM_R_X3Y119_SLICE_X3Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y120_SLICE_X2Y120_AO6),
.Q(CLBLM_R_X3Y120_SLICE_X2Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y120_SLICE_X2Y120_BO6),
.Q(CLBLM_R_X3Y120_SLICE_X2Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y120_SLICE_X2Y120_CO6),
.Q(CLBLM_R_X3Y120_SLICE_X2Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaff00ff00ff)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_DLUT (
.I0(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(1'b1),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_CQ),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_DO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f055f0aa)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_CLUT (
.I0(CLBLL_L_X4Y120_SLICE_X4Y120_BQ),
.I1(1'b1),
.I2(CLBLL_L_X2Y121_SLICE_X1Y121_B5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y120_SLICE_X2Y120_DO6),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_CO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000cc00cc)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y120_SLICE_X2Y120_BQ),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLL_L_X4Y120_SLICE_X4Y120_C5Q),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_BO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddc1110fffc3330)
  ) CLBLM_R_X3Y120_SLICE_X2Y120_ALUT (
.I0(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y120_SLICE_X2Y120_AQ),
.I3(CLBLM_R_X3Y121_SLICE_X3Y121_BQ),
.I4(CLBLM_R_X3Y118_SLICE_X3Y118_AQ),
.I5(CLBLL_L_X4Y125_SLICE_X4Y125_BQ),
.O5(CLBLM_R_X3Y120_SLICE_X2Y120_AO5),
.O6(CLBLM_R_X3Y120_SLICE_X2Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y120_SLICE_X3Y120_AO6),
.Q(CLBLM_R_X3Y120_SLICE_X3Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y120_SLICE_X3Y120_BO6),
.Q(CLBLM_R_X3Y120_SLICE_X3Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffa0a0a0a0a0a0)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_DLUT (
.I0(CLBLM_R_X3Y126_SLICE_X3Y126_AO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y121_SLICE_X2Y121_CQ),
.I3(1'b1),
.I4(CLBLM_R_X3Y125_SLICE_X2Y125_AQ),
.I5(CLBLM_R_X3Y130_SLICE_X3Y130_BO6),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_DO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1155b1f55555f5f5)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLL_L_X4Y125_SLICE_X4Y125_BQ),
.I2(CLBLM_R_X3Y119_SLICE_X3Y119_DO6),
.I3(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.I4(CLBLM_R_X3Y120_SLICE_X3Y120_DO6),
.I5(CLBLM_R_X3Y127_SLICE_X2Y127_DO6),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_CO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0f3c0c0c0f3c0)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y120_SLICE_X3Y120_AQ),
.I3(CLBLM_R_X5Y121_SLICE_X7Y121_AQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_BO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0074743030)
  ) CLBLM_R_X3Y120_SLICE_X3Y120_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLL_L_X4Y117_SLICE_X4Y117_AO5),
.I2(CLBLM_R_X3Y120_SLICE_X3Y120_AQ),
.I3(CLBLL_L_X4Y120_SLICE_X4Y120_BQ),
.I4(CLBLM_R_X3Y126_SLICE_X3Y126_AO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y120_SLICE_X3Y120_AO5),
.O6(CLBLM_R_X3Y120_SLICE_X3Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y121_SLICE_X2Y121_CO5),
.Q(CLBLM_R_X3Y121_SLICE_X2Y121_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y121_SLICE_X2Y121_AO6),
.Q(CLBLM_R_X3Y121_SLICE_X2Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y121_SLICE_X2Y121_BO6),
.Q(CLBLM_R_X3Y121_SLICE_X2Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y121_SLICE_X2Y121_CO6),
.Q(CLBLM_R_X3Y121_SLICE_X2Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000aa6aaaaa)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_DLUT (
.I0(CLBLM_R_X3Y121_SLICE_X2Y121_C5Q),
.I1(CLBLL_L_X2Y121_SLICE_X0Y121_BQ),
.I2(CLBLM_R_X3Y121_SLICE_X2Y121_BQ),
.I3(CLBLM_R_X11Y120_SLICE_X14Y120_DO6),
.I4(CLBLM_R_X3Y121_SLICE_X2Y121_AQ),
.I5(CLBLL_L_X2Y121_SLICE_X1Y121_CO6),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_DO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf303f303ffffa0a0)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_CLUT (
.I0(CLBLL_L_X4Y119_SLICE_X4Y119_AQ),
.I1(CLBLM_R_X11Y120_SLICE_X14Y120_DO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y120_SLICE_X12Y120_CQ),
.I4(CLBLM_R_X3Y121_SLICE_X2Y121_DO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_CO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hefcc2300dccc1000)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_BLUT (
.I0(CLBLL_L_X2Y121_SLICE_X1Y121_AO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y121_SLICE_X2Y121_AQ),
.I3(CLBLL_L_X2Y121_SLICE_X1Y121_DO6),
.I4(CLBLM_L_X10Y125_SLICE_X13Y125_BQ),
.I5(CLBLM_R_X3Y121_SLICE_X2Y121_BQ),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_BO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcca5cca5cc00cc00)
  ) CLBLM_R_X3Y121_SLICE_X2Y121_ALUT (
.I0(CLBLL_L_X2Y121_SLICE_X1Y121_AO5),
.I1(CLBLM_R_X3Y120_SLICE_X2Y120_BQ),
.I2(CLBLM_R_X3Y121_SLICE_X2Y121_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLL_L_X2Y121_SLICE_X1Y121_DO6),
.O5(CLBLM_R_X3Y121_SLICE_X2Y121_AO5),
.O6(CLBLM_R_X3Y121_SLICE_X2Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y121_SLICE_X3Y121_AO6),
.Q(CLBLM_R_X3Y121_SLICE_X3Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y121_SLICE_X3Y121_BO6),
.Q(CLBLM_R_X3Y121_SLICE_X3Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc000000cc000000)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y122_SLICE_X7Y122_AQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I4(CLBLM_R_X5Y122_SLICE_X6Y122_DO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_DO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000080008000)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_CLUT (
.I0(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I1(CLBLM_R_X5Y122_SLICE_X7Y122_AQ),
.I2(CLBLM_R_X3Y121_SLICE_X3Y121_BQ),
.I3(CLBLM_R_X5Y122_SLICE_X6Y122_DO6),
.I4(CLBLM_R_X3Y121_SLICE_X3Y121_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_CO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f000fe0e)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_BLUT (
.I0(CLBLM_R_X3Y121_SLICE_X3Y121_DO6),
.I1(CLBLM_R_X3Y121_SLICE_X3Y121_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.I4(CLBLM_R_X3Y121_SLICE_X3Y121_CO5),
.I5(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_BO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00cc55cc50)
  ) CLBLM_R_X3Y121_SLICE_X3Y121_ALUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.I1(CLBLM_R_X5Y123_SLICE_X7Y123_BQ),
.I2(CLBLM_R_X3Y121_SLICE_X3Y121_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y121_SLICE_X3Y121_CO5),
.I5(CLBLM_R_X3Y121_SLICE_X3Y121_CO6),
.O5(CLBLM_R_X3Y121_SLICE_X3Y121_AO5),
.O6(CLBLM_R_X3Y121_SLICE_X3Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y122_SLICE_X2Y122_BO6),
.Q(CLBLM_R_X3Y122_SLICE_X2Y122_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y122_SLICE_X2Y122_AO6),
.Q(CLBLM_R_X3Y122_SLICE_X2Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y122_SLICE_X2Y122_CO6),
.Q(CLBLM_R_X3Y122_SLICE_X2Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y122_SLICE_X2Y122_DO6),
.Q(CLBLM_R_X3Y122_SLICE_X2Y122_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ddd0ddd0)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_DLUT (
.I0(CLBLM_R_X7Y123_SLICE_X9Y123_A5Q),
.I1(CLBLM_R_X11Y120_SLICE_X14Y120_DO6),
.I2(CLBLM_R_X3Y122_SLICE_X2Y122_DQ),
.I3(CLBLM_R_X5Y122_SLICE_X7Y122_AQ),
.I4(CLBLM_R_X3Y121_SLICE_X3Y121_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_DO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa003c00cc)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_CLUT (
.I0(CLBLM_L_X10Y121_SLICE_X12Y121_C5Q),
.I1(CLBLM_R_X3Y122_SLICE_X2Y122_CQ),
.I2(CLBLM_R_X5Y123_SLICE_X7Y123_BQ),
.I3(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.I4(CLBLM_R_X3Y122_SLICE_X2Y122_BO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_CO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00fe3250505050)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_BLUT (
.I0(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLL_L_X2Y126_SLICE_X1Y126_AQ),
.I4(CLBLM_R_X7Y122_SLICE_X8Y122_DO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_BO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaaaaaffa0a0a0)
  ) CLBLM_R_X3Y122_SLICE_X2Y122_ALUT (
.I0(CLBLM_R_X5Y126_SLICE_X7Y126_CO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y122_SLICE_X2Y122_AQ),
.I3(CLBLL_L_X4Y122_SLICE_X5Y122_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.O5(CLBLM_R_X3Y122_SLICE_X2Y122_AO5),
.O6(CLBLM_R_X3Y122_SLICE_X2Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y122_SLICE_X3Y122_AO6),
.Q(CLBLM_R_X3Y122_SLICE_X3Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y122_SLICE_X3Y122_BO6),
.Q(CLBLM_R_X3Y122_SLICE_X3Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ffffffffffffff)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_DLUT (
.I0(CLBLM_R_X3Y121_SLICE_X3Y121_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X3Y122_SLICE_X2Y122_CQ),
.I4(CLBLM_R_X5Y123_SLICE_X7Y123_BQ),
.I5(CLBLM_R_X3Y121_SLICE_X3Y121_BQ),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_DO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f3f5ff3333ffff)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_CLUT (
.I0(CLBLM_R_X3Y121_SLICE_X3Y121_AQ),
.I1(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I2(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.I3(CLBLM_R_X3Y121_SLICE_X3Y121_BQ),
.I4(CLBLM_R_X5Y122_SLICE_X7Y122_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_CO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haafcaafcaa00aafc)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_BLUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_DQ),
.I1(CLBLM_R_X3Y122_SLICE_X3Y122_BQ),
.I2(CLBLM_R_X3Y123_SLICE_X3Y123_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y123_SLICE_X9Y123_A5Q),
.I5(CLBLM_R_X11Y120_SLICE_X14Y120_DO6),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_BO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3afa3afa3afa0a0)
  ) CLBLM_R_X3Y122_SLICE_X3Y122_ALUT (
.I0(CLBLM_R_X5Y123_SLICE_X6Y123_B5Q),
.I1(CLBLL_L_X4Y125_SLICE_X4Y125_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.I4(CLBLM_R_X3Y121_SLICE_X3Y121_AQ),
.I5(CLBLM_R_X3Y122_SLICE_X3Y122_AQ),
.O5(CLBLM_R_X3Y122_SLICE_X3Y122_AO5),
.O6(CLBLM_R_X3Y122_SLICE_X3Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y123_SLICE_X2Y123_AO6),
.Q(CLBLM_R_X3Y123_SLICE_X2Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y123_SLICE_X2Y123_BO6),
.Q(CLBLM_R_X3Y123_SLICE_X2Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y123_SLICE_X2Y123_CO6),
.Q(CLBLM_R_X3Y123_SLICE_X2Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y123_SLICE_X2Y123_DO6),
.Q(CLBLM_R_X3Y123_SLICE_X2Y123_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ccccd8d8)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_DLUT (
.I0(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I1(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.I2(CLBLM_R_X3Y123_SLICE_X2Y123_DQ),
.I3(CLBLM_R_X3Y132_SLICE_X2Y132_A5Q),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_DO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'habaeaaaa01040000)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y123_SLICE_X2Y123_CQ),
.I2(CLBLL_L_X2Y118_SLICE_X1Y118_AQ),
.I3(CLBLM_R_X3Y132_SLICE_X2Y132_A5Q),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X5Y117_SLICE_X6Y117_A5Q),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_CO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaacfcfc0c0)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_BLUT (
.I0(CLBLM_R_X3Y122_SLICE_X2Y122_DQ),
.I1(CLBLM_R_X3Y123_SLICE_X2Y123_BQ),
.I2(CLBLM_R_X5Y126_SLICE_X7Y126_CO5),
.I3(1'b1),
.I4(CLBLL_L_X4Y120_SLICE_X4Y120_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_BO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f7f78080)
  ) CLBLM_R_X3Y123_SLICE_X2Y123_ALUT (
.I0(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.I1(CLBLL_L_X4Y125_SLICE_X4Y125_BQ),
.I2(CLBLM_R_X3Y123_SLICE_X2Y123_AQ),
.I3(CLBLM_R_X3Y122_SLICE_X2Y122_AQ),
.I4(CLBLM_R_X3Y122_SLICE_X2Y122_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y123_SLICE_X2Y123_AO5),
.O6(CLBLM_R_X3Y123_SLICE_X2Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y123_SLICE_X3Y123_AO6),
.Q(CLBLM_R_X3Y123_SLICE_X3Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y123_SLICE_X3Y123_BO6),
.Q(CLBLM_R_X3Y123_SLICE_X3Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y123_SLICE_X3Y123_CO6),
.Q(CLBLM_R_X3Y123_SLICE_X3Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4040000040400000)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_DLUT (
.I0(CLBLL_L_X4Y120_SLICE_X5Y120_BQ),
.I1(CLBLM_R_X3Y123_SLICE_X3Y123_AQ),
.I2(CLBLM_R_X5Y123_SLICE_X6Y123_B5Q),
.I3(1'b1),
.I4(CLBLL_L_X4Y120_SLICE_X5Y120_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_DO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb888888888888888)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_CLUT (
.I0(CLBLM_R_X5Y124_SLICE_X7Y124_C5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y121_SLICE_X2Y121_C5Q),
.I3(CLBLL_L_X2Y121_SLICE_X0Y121_BQ),
.I4(CLBLM_R_X3Y121_SLICE_X2Y121_AQ),
.I5(CLBLM_R_X3Y121_SLICE_X2Y121_BQ),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_CO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0000002020)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_BLUT (
.I0(CLBLM_R_X3Y123_SLICE_X3Y123_DO6),
.I1(CLBLM_R_X3Y122_SLICE_X3Y122_DO6),
.I2(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.I3(CLBLM_R_X5Y126_SLICE_X7Y126_BQ),
.I4(CLBLM_R_X3Y122_SLICE_X3Y122_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_BO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcd01cd01dc10dc10)
  ) CLBLM_R_X3Y123_SLICE_X3Y123_ALUT (
.I0(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y123_SLICE_X3Y123_AQ),
.I3(CLBLM_R_X3Y125_SLICE_X3Y125_AQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y121_SLICE_X3Y121_CO6),
.O5(CLBLM_R_X3Y123_SLICE_X3Y123_AO5),
.O6(CLBLM_R_X3Y123_SLICE_X3Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y124_SLICE_X2Y124_AO5),
.Q(CLBLM_R_X3Y124_SLICE_X2Y124_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y124_SLICE_X2Y124_BO5),
.Q(CLBLM_R_X3Y124_SLICE_X2Y124_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y124_SLICE_X2Y124_AO6),
.Q(CLBLM_R_X3Y124_SLICE_X2Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y124_SLICE_X2Y124_BO6),
.Q(CLBLM_R_X3Y124_SLICE_X2Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y124_SLICE_X2Y124_CO6),
.Q(CLBLM_R_X3Y124_SLICE_X2Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y124_SLICE_X2Y124_DO6),
.Q(CLBLM_R_X3Y124_SLICE_X2Y124_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefeaaaafcfc0000)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y120_SLICE_X5Y120_A5Q),
.I2(CLBLM_R_X3Y124_SLICE_X2Y124_DQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y126_SLICE_X7Y126_CO6),
.I5(CLBLM_R_X3Y132_SLICE_X2Y132_BQ),
.O5(CLBLM_R_X3Y124_SLICE_X2Y124_DO5),
.O6(CLBLM_R_X3Y124_SLICE_X2Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0f5a0a0a0a0a0a0)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLL_L_X4Y121_SLICE_X4Y121_BQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.I5(CLBLL_L_X4Y125_SLICE_X4Y125_BQ),
.O5(CLBLM_R_X3Y124_SLICE_X2Y124_CO5),
.O6(CLBLM_R_X3Y124_SLICE_X2Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0acacacac)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_BLUT (
.I0(CLBLL_L_X2Y118_SLICE_X1Y118_AQ),
.I1(CLBLM_R_X5Y123_SLICE_X6Y123_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X3Y126_SLICE_X3Y126_AO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X2Y124_BO5),
.O6(CLBLM_R_X3Y124_SLICE_X2Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacacacfff00f00)
  ) CLBLM_R_X3Y124_SLICE_X2Y124_ALUT (
.I0(CLBLM_R_X3Y124_SLICE_X2Y124_CQ),
.I1(CLBLM_R_X3Y127_SLICE_X2Y127_DO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y128_SLICE_X3Y128_BO6),
.I4(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X2Y124_AO5),
.O6(CLBLM_R_X3Y124_SLICE_X2Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y124_SLICE_X3Y124_CO5),
.Q(CLBLM_R_X3Y124_SLICE_X3Y124_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y124_SLICE_X3Y124_AO6),
.Q(CLBLM_R_X3Y124_SLICE_X3Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y124_SLICE_X3Y124_BO6),
.Q(CLBLM_R_X3Y124_SLICE_X3Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y124_SLICE_X3Y124_CO6),
.Q(CLBLM_R_X3Y124_SLICE_X3Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffbfffb)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_DLUT (
.I0(CLBLM_R_X3Y125_SLICE_X3Y125_CO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X3Y124_SLICE_X2Y124_B5Q),
.I3(CLBLL_L_X4Y123_SLICE_X5Y123_B5Q),
.I4(1'b1),
.I5(CLBLM_R_X5Y125_SLICE_X6Y125_A5Q),
.O5(CLBLM_R_X3Y124_SLICE_X3Y124_DO5),
.O6(CLBLM_R_X3Y124_SLICE_X3Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbaba1010f5a0f5a0)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLL_L_X4Y120_SLICE_X5Y120_A5Q),
.I3(CLBLM_R_X3Y124_SLICE_X2Y124_CQ),
.I4(CLBLL_L_X4Y124_SLICE_X4Y124_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y124_SLICE_X3Y124_CO5),
.O6(CLBLM_R_X3Y124_SLICE_X3Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0eeeef0f04444)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_BLUT (
.I0(CLBLM_R_X5Y126_SLICE_X7Y126_CO5),
.I1(CLBLM_R_X3Y124_SLICE_X3Y124_BQ),
.I2(CLBLM_R_X3Y124_SLICE_X3Y124_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y121_SLICE_X4Y121_DQ),
.O5(CLBLM_R_X3Y124_SLICE_X3Y124_BO5),
.O6(CLBLM_R_X3Y124_SLICE_X3Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf0ccffcc00)
  ) CLBLM_R_X3Y124_SLICE_X3Y124_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y124_SLICE_X4Y124_AQ),
.I2(CLBLM_R_X3Y124_SLICE_X3Y124_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y124_SLICE_X11Y124_BQ),
.I5(CLBLM_L_X10Y129_SLICE_X13Y129_DO6),
.O5(CLBLM_R_X3Y124_SLICE_X3Y124_AO5),
.O6(CLBLM_R_X3Y124_SLICE_X3Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y125_SLICE_X2Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y125_SLICE_X2Y125_AO6),
.Q(CLBLM_R_X3Y125_SLICE_X2Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffaaaaaaaa)
  ) CLBLM_R_X3Y125_SLICE_X2Y125_DLUT (
.I0(CLBLM_R_X5Y123_SLICE_X7Y123_C5Q),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X3Y124_SLICE_X2Y124_B5Q),
.O5(CLBLM_R_X3Y125_SLICE_X2Y125_DO5),
.O6(CLBLM_R_X3Y125_SLICE_X2Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffef)
  ) CLBLM_R_X3Y125_SLICE_X2Y125_CLUT (
.I0(CLBLL_L_X2Y121_SLICE_X1Y121_BQ),
.I1(CLBLM_R_X5Y123_SLICE_X7Y123_C5Q),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X3Y124_SLICE_X2Y124_B5Q),
.I4(CLBLM_R_X5Y127_SLICE_X7Y127_B5Q),
.I5(CLBLM_R_X7Y126_SLICE_X9Y126_D5Q),
.O5(CLBLM_R_X3Y125_SLICE_X2Y125_CO5),
.O6(CLBLM_R_X3Y125_SLICE_X2Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000010000)
  ) CLBLM_R_X3Y125_SLICE_X2Y125_BLUT (
.I0(CLBLM_R_X3Y125_SLICE_X2Y125_DO6),
.I1(CLBLM_R_X3Y126_SLICE_X2Y126_BO6),
.I2(CLBLM_R_X5Y127_SLICE_X7Y127_B5Q),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_D5Q),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLL_L_X2Y125_SLICE_X1Y125_DO6),
.O5(CLBLM_R_X3Y125_SLICE_X2Y125_BO5),
.O6(CLBLM_R_X3Y125_SLICE_X2Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff007878ff00f0f0)
  ) CLBLM_R_X3Y125_SLICE_X2Y125_ALUT (
.I0(CLBLL_L_X2Y126_SLICE_X1Y126_AQ),
.I1(CLBLM_R_X3Y130_SLICE_X2Y130_AO5),
.I2(CLBLL_L_X2Y118_SLICE_X1Y118_AQ),
.I3(CLBLM_R_X3Y122_SLICE_X2Y122_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X2Y125_SLICE_X1Y125_AQ),
.O5(CLBLM_R_X3Y125_SLICE_X2Y125_AO5),
.O6(CLBLM_R_X3Y125_SLICE_X2Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y125_SLICE_X3Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y125_SLICE_X3Y125_AO6),
.Q(CLBLM_R_X3Y125_SLICE_X3Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y125_SLICE_X3Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y125_SLICE_X3Y125_BO6),
.Q(CLBLM_R_X3Y125_SLICE_X3Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0aff0aff0a0a0a0a)
  ) CLBLM_R_X3Y125_SLICE_X3Y125_DLUT (
.I0(CLBLM_R_X3Y124_SLICE_X3Y124_AQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y126_SLICE_X4Y126_BO6),
.I3(CLBLL_L_X2Y129_SLICE_X0Y129_AO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y120_SLICE_X2Y120_AQ),
.O5(CLBLM_R_X3Y125_SLICE_X3Y125_DO5),
.O6(CLBLM_R_X3Y125_SLICE_X3Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X3Y125_SLICE_X3Y125_CLUT (
.I0(CLBLM_R_X5Y127_SLICE_X7Y127_B5Q),
.I1(CLBLM_R_X7Y126_SLICE_X9Y126_D5Q),
.I2(CLBLM_R_X3Y126_SLICE_X2Y126_A5Q),
.I3(CLBLL_L_X2Y122_SLICE_X1Y122_A5Q),
.I4(CLBLM_R_X5Y123_SLICE_X7Y123_C5Q),
.I5(CLBLL_L_X2Y121_SLICE_X1Y121_BQ),
.O5(CLBLM_R_X3Y125_SLICE_X3Y125_CO5),
.O6(CLBLM_R_X3Y125_SLICE_X3Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000fe0efe0e)
  ) CLBLM_R_X3Y125_SLICE_X3Y125_BLUT (
.I0(CLBLM_R_X5Y122_SLICE_X6Y122_CQ),
.I1(CLBLM_R_X3Y125_SLICE_X3Y125_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X2Y125_SLICE_X1Y125_AQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y126_SLICE_X7Y126_CO6),
.O5(CLBLM_R_X3Y125_SLICE_X3Y125_BO5),
.O6(CLBLM_R_X3Y125_SLICE_X3Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffa500000fa50)
  ) CLBLM_R_X3Y125_SLICE_X3Y125_ALUT (
.I0(CLBLM_L_X10Y129_SLICE_X13Y129_DO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y125_SLICE_X3Y125_AQ),
.I3(CLBLL_L_X4Y125_SLICE_X4Y125_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X2Y121_SLICE_X0Y121_BQ),
.O5(CLBLM_R_X3Y125_SLICE_X3Y125_AO5),
.O6(CLBLM_R_X3Y125_SLICE_X3Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y126_SLICE_X2Y126_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y130_SLICE_X2Y130_AO6),
.Q(CLBLM_R_X3Y126_SLICE_X2Y126_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y126_SLICE_X2Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y126_SLICE_X2Y126_AO6),
.Q(CLBLM_R_X3Y126_SLICE_X2Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55f5ddfd00f0ccfc)
  ) CLBLM_R_X3Y126_SLICE_X2Y126_DLUT (
.I0(CLBLL_L_X2Y126_SLICE_X0Y126_AO6),
.I1(CLBLL_L_X4Y119_SLICE_X4Y119_DQ),
.I2(LIOB33_X0Y63_IOB_X0Y63_I),
.I3(CLBLL_L_X2Y130_SLICE_X1Y130_BO6),
.I4(CLBLL_L_X2Y126_SLICE_X0Y126_AO5),
.I5(CLBLL_L_X4Y124_SLICE_X5Y124_DQ),
.O5(CLBLM_R_X3Y126_SLICE_X2Y126_DO5),
.O6(CLBLM_R_X3Y126_SLICE_X2Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00aaaeae0cae)
  ) CLBLM_R_X3Y126_SLICE_X2Y126_CLUT (
.I0(CLBLM_R_X3Y124_SLICE_X2Y124_AQ),
.I1(CLBLM_R_X3Y126_SLICE_X2Y126_AQ),
.I2(CLBLL_L_X2Y130_SLICE_X0Y130_CO6),
.I3(RIOB33_X105Y137_IOB_X1Y137_I),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(CLBLL_L_X2Y128_SLICE_X1Y128_AO6),
.O5(CLBLM_R_X3Y126_SLICE_X2Y126_CO5),
.O6(CLBLM_R_X3Y126_SLICE_X2Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000002)
  ) CLBLM_R_X3Y126_SLICE_X2Y126_BLUT (
.I0(CLBLM_R_X3Y129_SLICE_X2Y129_CO6),
.I1(CLBLL_L_X4Y126_SLICE_X4Y126_DO6),
.I2(CLBLM_R_X3Y126_SLICE_X3Y126_AO6),
.I3(CLBLM_R_X3Y128_SLICE_X3Y128_BO6),
.I4(CLBLL_L_X4Y128_SLICE_X4Y128_AO6),
.I5(CLBLL_L_X2Y127_SLICE_X1Y127_CO6),
.O5(CLBLM_R_X3Y126_SLICE_X2Y126_BO5),
.O6(CLBLM_R_X3Y126_SLICE_X2Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccfc00330030)
  ) CLBLM_R_X3Y126_SLICE_X2Y126_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y126_SLICE_X2Y126_AQ),
.I3(CLBLL_L_X2Y119_SLICE_X1Y119_BO6),
.I4(CLBLM_R_X3Y126_SLICE_X2Y126_A5Q),
.I5(CLBLM_R_X3Y124_SLICE_X2Y124_A5Q),
.O5(CLBLM_R_X3Y126_SLICE_X2Y126_AO5),
.O6(CLBLM_R_X3Y126_SLICE_X2Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5d5d5d5d0c0c0c0c)
  ) CLBLM_R_X3Y126_SLICE_X3Y126_DLUT (
.I0(CLBLM_R_X3Y130_SLICE_X3Y130_AO6),
.I1(CLBLM_L_X10Y128_SLICE_X12Y128_DQ),
.I2(CLBLL_L_X4Y126_SLICE_X4Y126_BO5),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X3Y120_SLICE_X3Y120_AQ),
.O5(CLBLM_R_X3Y126_SLICE_X3Y126_DO5),
.O6(CLBLM_R_X3Y126_SLICE_X3Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff1100ffff3130)
  ) CLBLM_R_X3Y126_SLICE_X3Y126_CLUT (
.I0(CLBLL_L_X2Y130_SLICE_X0Y130_BO6),
.I1(CLBLL_L_X2Y130_SLICE_X0Y130_CO6),
.I2(CLBLM_R_X5Y126_SLICE_X6Y126_DQ),
.I3(LIOB33_X0Y65_IOB_X0Y66_I),
.I4(CLBLL_L_X2Y125_SLICE_X1Y125_CO5),
.I5(CLBLL_L_X2Y128_SLICE_X1Y128_AO6),
.O5(CLBLM_R_X3Y126_SLICE_X3Y126_CO5),
.O6(CLBLM_R_X3Y126_SLICE_X3Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffcceefcfe)
  ) CLBLM_R_X3Y126_SLICE_X3Y126_BLUT (
.I0(CLBLM_R_X7Y126_SLICE_X8Y126_AQ),
.I1(CLBLM_R_X3Y127_SLICE_X3Y127_CO6),
.I2(CLBLM_R_X3Y122_SLICE_X3Y122_AQ),
.I3(CLBLL_L_X4Y126_SLICE_X4Y126_BO6),
.I4(CLBLL_L_X2Y129_SLICE_X0Y129_AO6),
.I5(CLBLM_R_X3Y126_SLICE_X3Y126_CO6),
.O5(CLBLM_R_X3Y126_SLICE_X3Y126_BO5),
.O6(CLBLM_R_X3Y126_SLICE_X3Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X3Y126_SLICE_X3Y126_ALUT (
.I0(CLBLM_R_X3Y126_SLICE_X3Y126_DO6),
.I1(CLBLM_R_X3Y126_SLICE_X2Y126_DO6),
.I2(CLBLL_L_X2Y129_SLICE_X1Y129_CO6),
.I3(CLBLL_L_X4Y127_SLICE_X5Y127_AO6),
.I4(CLBLL_L_X4Y125_SLICE_X4Y125_DO6),
.I5(CLBLL_L_X2Y126_SLICE_X1Y126_DO6),
.O5(CLBLM_R_X3Y126_SLICE_X3Y126_AO5),
.O6(CLBLM_R_X3Y126_SLICE_X3Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffbbffbb)
  ) CLBLM_R_X3Y127_SLICE_X2Y127_DLUT (
.I0(CLBLM_R_X3Y127_SLICE_X2Y127_CO6),
.I1(CLBLL_L_X2Y129_SLICE_X1Y129_BO6),
.I2(1'b1),
.I3(CLBLL_L_X4Y125_SLICE_X5Y125_CO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y127_SLICE_X2Y127_BO6),
.O5(CLBLM_R_X3Y127_SLICE_X2Y127_DO5),
.O6(CLBLM_R_X3Y127_SLICE_X2Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffceffcece)
  ) CLBLM_R_X3Y127_SLICE_X2Y127_CLUT (
.I0(CLBLM_R_X3Y122_SLICE_X3Y122_BQ),
.I1(CLBLM_R_X3Y126_SLICE_X2Y126_CO6),
.I2(CLBLL_L_X4Y129_SLICE_X4Y129_BO6),
.I3(CLBLM_R_X3Y130_SLICE_X2Y130_BO6),
.I4(CLBLM_R_X3Y125_SLICE_X3Y125_BQ),
.I5(CLBLL_L_X2Y127_SLICE_X1Y127_DO6),
.O5(CLBLM_R_X3Y127_SLICE_X2Y127_CO5),
.O6(CLBLM_R_X3Y127_SLICE_X2Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ace0aceffff0ace)
  ) CLBLM_R_X3Y127_SLICE_X2Y127_BLUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(CLBLL_L_X4Y125_SLICE_X5Y125_BQ),
.I2(CLBLM_R_X3Y129_SLICE_X3Y129_AO6),
.I3(CLBLL_L_X4Y129_SLICE_X4Y129_BO5),
.I4(CLBLL_L_X4Y120_SLICE_X4Y120_AQ),
.I5(CLBLL_L_X2Y128_SLICE_X0Y128_AO6),
.O5(CLBLM_R_X3Y127_SLICE_X2Y127_BO5),
.O6(CLBLM_R_X3Y127_SLICE_X2Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0004000400050000)
  ) CLBLM_R_X3Y127_SLICE_X2Y127_ALUT (
.I0(CLBLL_L_X2Y130_SLICE_X0Y130_AO6),
.I1(CLBLL_L_X4Y125_SLICE_X5Y125_BQ),
.I2(CLBLL_L_X4Y130_SLICE_X4Y130_AO5),
.I3(RIOB33_X105Y135_IOB_X1Y135_I),
.I4(CLBLL_L_X4Y120_SLICE_X4Y120_AQ),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLM_R_X3Y127_SLICE_X2Y127_AO5),
.O6(CLBLM_R_X3Y127_SLICE_X2Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1111515100005050)
  ) CLBLM_R_X3Y127_SLICE_X3Y127_DLUT (
.I0(CLBLL_L_X2Y130_SLICE_X0Y130_CO6),
.I1(CLBLL_L_X2Y128_SLICE_X1Y128_AO5),
.I2(CLBLM_R_X3Y119_SLICE_X2Y119_AQ),
.I3(1'b1),
.I4(CLBLL_L_X2Y130_SLICE_X0Y130_AO6),
.I5(LIOB33_X0Y71_IOB_X0Y71_I),
.O5(CLBLM_R_X3Y127_SLICE_X3Y127_DO5),
.O6(CLBLM_R_X3Y127_SLICE_X3Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000f0222222f2)
  ) CLBLM_R_X3Y127_SLICE_X3Y127_CLUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I1(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(CLBLL_L_X2Y130_SLICE_X0Y130_BO6),
.I4(CLBLL_L_X2Y130_SLICE_X0Y130_CO5),
.I5(CLBLL_L_X2Y128_SLICE_X1Y128_AO6),
.O5(CLBLM_R_X3Y127_SLICE_X3Y127_CO5),
.O6(CLBLM_R_X3Y127_SLICE_X3Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffaaeefafe)
  ) CLBLM_R_X3Y127_SLICE_X3Y127_BLUT (
.I0(CLBLL_L_X4Y127_SLICE_X5Y127_DO6),
.I1(CLBLL_L_X4Y121_SLICE_X4Y121_BQ),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(CLBLL_L_X2Y128_SLICE_X0Y128_AO6),
.I4(CLBLM_R_X3Y129_SLICE_X3Y129_AO6),
.I5(CLBLM_R_X3Y127_SLICE_X3Y127_AO6),
.O5(CLBLM_R_X3Y127_SLICE_X3Y127_BO5),
.O6(CLBLM_R_X3Y127_SLICE_X3Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000020)
  ) CLBLM_R_X3Y127_SLICE_X3Y127_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_L_X10Y123_SLICE_X12Y123_AQ),
.I3(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X3Y127_SLICE_X3Y127_AO5),
.O6(CLBLM_R_X3Y127_SLICE_X3Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5fdf5fdf0fcf0fc)
  ) CLBLM_R_X3Y128_SLICE_X2Y128_DLUT (
.I0(CLBLL_L_X2Y128_SLICE_X0Y128_BO6),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y129_SLICE_X3Y129_DO6),
.I3(CLBLL_L_X2Y130_SLICE_X1Y130_BO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y119_SLICE_X2Y119_BQ),
.O5(CLBLM_R_X3Y128_SLICE_X2Y128_DO5),
.O6(CLBLM_R_X3Y128_SLICE_X2Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf4fff4fff4f4f4f4)
  ) CLBLM_R_X3Y128_SLICE_X2Y128_CLUT (
.I0(CLBLL_L_X2Y126_SLICE_X0Y126_AO6),
.I1(CLBLM_R_X5Y127_SLICE_X7Y127_CQ),
.I2(CLBLL_L_X2Y129_SLICE_X0Y129_DO6),
.I3(CLBLM_R_X3Y129_SLICE_X3Y129_AO5),
.I4(1'b1),
.I5(RIOB33_X105Y113_IOB_X1Y114_I),
.O5(CLBLM_R_X3Y128_SLICE_X2Y128_CO5),
.O6(CLBLM_R_X3Y128_SLICE_X2Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffeefeaafa)
  ) CLBLM_R_X3Y128_SLICE_X2Y128_BLUT (
.I0(CLBLL_L_X2Y129_SLICE_X0Y129_CO6),
.I1(CLBLL_L_X4Y124_SLICE_X4Y124_A5Q),
.I2(CLBLL_L_X4Y129_SLICE_X5Y129_AQ),
.I3(CLBLL_L_X2Y126_SLICE_X0Y126_AO5),
.I4(CLBLL_L_X2Y118_SLICE_X1Y118_CO6),
.I5(CLBLL_L_X2Y128_SLICE_X0Y128_DO6),
.O5(CLBLM_R_X3Y128_SLICE_X2Y128_BO5),
.O6(CLBLM_R_X3Y128_SLICE_X2Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X3Y128_SLICE_X2Y128_ALUT (
.I0(CLBLM_L_X8Y130_SLICE_X11Y130_DO6),
.I1(CLBLL_L_X4Y126_SLICE_X5Y126_AO6),
.I2(CLBLM_R_X3Y128_SLICE_X2Y128_BO6),
.I3(CLBLL_L_X4Y128_SLICE_X5Y128_CO6),
.I4(CLBLL_L_X2Y129_SLICE_X1Y129_CO6),
.I5(CLBLM_R_X3Y128_SLICE_X2Y128_CO6),
.O5(CLBLM_R_X3Y128_SLICE_X2Y128_AO5),
.O6(CLBLM_R_X3Y128_SLICE_X2Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff3300f3f0)
  ) CLBLM_R_X3Y128_SLICE_X3Y128_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y129_SLICE_X3Y129_AO5),
.I2(CLBLM_R_X5Y128_SLICE_X6Y128_DQ),
.I3(RIOB33_X105Y115_IOB_X1Y115_I),
.I4(CLBLL_L_X2Y126_SLICE_X0Y126_AO5),
.I5(CLBLL_L_X2Y130_SLICE_X0Y130_DO6),
.O5(CLBLM_R_X3Y128_SLICE_X3Y128_DO5),
.O6(CLBLM_R_X3Y128_SLICE_X3Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdcffdcffffffdc)
  ) CLBLM_R_X3Y128_SLICE_X3Y128_CLUT (
.I0(CLBLL_L_X2Y126_SLICE_X0Y126_AO6),
.I1(CLBLL_L_X2Y126_SLICE_X0Y126_CO6),
.I2(CLBLL_L_X4Y129_SLICE_X4Y129_AQ),
.I3(CLBLM_R_X3Y130_SLICE_X3Y130_CO6),
.I4(CLBLL_L_X4Y120_SLICE_X4Y120_DQ),
.I5(CLBLL_L_X4Y129_SLICE_X4Y129_BO6),
.O5(CLBLM_R_X3Y128_SLICE_X3Y128_CO5),
.O6(CLBLM_R_X3Y128_SLICE_X3Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffefffefe)
  ) CLBLM_R_X3Y128_SLICE_X3Y128_BLUT (
.I0(CLBLM_R_X3Y125_SLICE_X3Y125_DO6),
.I1(CLBLL_L_X4Y126_SLICE_X5Y126_CO6),
.I2(CLBLM_R_X3Y127_SLICE_X3Y127_BO6),
.I3(CLBLL_L_X2Y128_SLICE_X1Y128_DO6),
.I4(CLBLL_L_X2Y129_SLICE_X1Y129_DO6),
.I5(CLBLM_R_X3Y128_SLICE_X3Y128_CO6),
.O5(CLBLM_R_X3Y128_SLICE_X3Y128_BO5),
.O6(CLBLM_R_X3Y128_SLICE_X3Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0505370500003300)
  ) CLBLM_R_X3Y128_SLICE_X3Y128_ALUT (
.I0(CLBLL_L_X2Y130_SLICE_X0Y130_CO5),
.I1(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.I2(CLBLL_L_X2Y130_SLICE_X0Y130_AO6),
.I3(CLBLM_R_X3Y124_SLICE_X3Y124_BQ),
.I4(CLBLL_L_X2Y130_SLICE_X0Y130_BO6),
.I5(CLBLL_L_X2Y121_SLICE_X0Y121_BQ),
.O5(CLBLM_R_X3Y128_SLICE_X3Y128_AO5),
.O6(CLBLM_R_X3Y128_SLICE_X3Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y129_SLICE_X2Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y129_SLICE_X2Y129_AO6),
.Q(CLBLM_R_X3Y129_SLICE_X2Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000050)
  ) CLBLM_R_X3Y129_SLICE_X2Y129_DLUT (
.I0(CLBLL_L_X2Y128_SLICE_X0Y128_CO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y130_SLICE_X2Y130_BO6),
.I3(CLBLM_R_X3Y130_SLICE_X3Y130_AO5),
.I4(CLBLL_L_X2Y130_SLICE_X1Y130_CO6),
.I5(CLBLL_L_X2Y129_SLICE_X0Y129_CO6),
.O5(CLBLM_R_X3Y129_SLICE_X2Y129_DO5),
.O6(CLBLM_R_X3Y129_SLICE_X2Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X3Y129_SLICE_X2Y129_CLUT (
.I0(CLBLL_L_X4Y128_SLICE_X5Y128_CO6),
.I1(CLBLL_L_X2Y129_SLICE_X1Y129_CO6),
.I2(CLBLL_L_X4Y126_SLICE_X5Y126_AO6),
.I3(CLBLL_L_X4Y130_SLICE_X4Y130_CO6),
.I4(CLBLM_R_X3Y129_SLICE_X2Y129_DO6),
.I5(CLBLM_R_X3Y129_SLICE_X2Y129_BO6),
.O5(CLBLM_R_X3Y129_SLICE_X2Y129_CO5),
.O6(CLBLM_R_X3Y129_SLICE_X2Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X3Y129_SLICE_X2Y129_BLUT (
.I0(CLBLM_L_X8Y130_SLICE_X11Y130_DO6),
.I1(CLBLM_R_X3Y129_SLICE_X3Y129_BO6),
.I2(CLBLM_R_X3Y129_SLICE_X3Y129_CO6),
.I3(CLBLL_L_X2Y128_SLICE_X1Y128_CO6),
.I4(CLBLL_L_X2Y128_SLICE_X0Y128_DO6),
.I5(CLBLL_L_X2Y129_SLICE_X0Y129_DO6),
.O5(CLBLM_R_X3Y129_SLICE_X2Y129_BO5),
.O6(CLBLM_R_X3Y129_SLICE_X2Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff48c048c048c0)
  ) CLBLM_R_X3Y129_SLICE_X2Y129_ALUT (
.I0(CLBLM_R_X3Y123_SLICE_X2Y123_CQ),
.I1(CLBLM_R_X3Y132_SLICE_X2Y132_CO5),
.I2(CLBLM_R_X3Y129_SLICE_X2Y129_AQ),
.I3(CLBLM_R_X3Y132_SLICE_X2Y132_A5Q),
.I4(CLBLL_L_X4Y129_SLICE_X4Y129_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X3Y129_SLICE_X2Y129_AO5),
.O6(CLBLM_R_X3Y129_SLICE_X2Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf00cf00df55cf00)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_DLUT (
.I0(CLBLL_L_X2Y128_SLICE_X1Y128_AO5),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(CLBLM_R_X7Y129_SLICE_X8Y129_A5Q),
.I4(RIOB33_X105Y115_IOB_X1Y116_I),
.I5(CLBLL_L_X2Y130_SLICE_X0Y130_CO5),
.O5(CLBLM_R_X3Y129_SLICE_X3Y129_DO5),
.O6(CLBLM_R_X3Y129_SLICE_X3Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000020000000)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_CLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(CLBLL_L_X2Y130_SLICE_X0Y130_CO6),
.I2(CLBLL_L_X4Y129_SLICE_X5Y129_AQ),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X3Y129_SLICE_X3Y129_CO5),
.O6(CLBLM_R_X3Y129_SLICE_X3Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a3a0a0a0a0a0a0)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_BLUT (
.I0(CLBLL_L_X4Y124_SLICE_X4Y124_A5Q),
.I1(CLBLM_R_X7Y128_SLICE_X9Y128_BO5),
.I2(CLBLL_L_X2Y118_SLICE_X1Y118_CO6),
.I3(RIOB33_X105Y129_IOB_X1Y130_I),
.I4(CLBLL_L_X2Y130_SLICE_X1Y130_AO5),
.I5(RIOB33_X105Y135_IOB_X1Y135_I),
.O5(CLBLM_R_X3Y129_SLICE_X3Y129_BO5),
.O6(CLBLM_R_X3Y129_SLICE_X3Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbfffffffefff)
  ) CLBLM_R_X3Y129_SLICE_X3Y129_ALUT (
.I0(CLBLL_L_X2Y130_SLICE_X0Y130_CO5),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y129_SLICE_X3Y129_AO5),
.O6(CLBLM_R_X3Y129_SLICE_X3Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000800000000)
  ) CLBLM_R_X3Y130_SLICE_X2Y130_DLUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(CLBLL_L_X2Y128_SLICE_X0Y128_BO6),
.I2(CLBLL_L_X2Y130_SLICE_X1Y130_CO6),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(CLBLM_R_X3Y130_SLICE_X2Y130_BO5),
.I5(CLBLM_R_X3Y130_SLICE_X2Y130_BO6),
.O5(CLBLM_R_X3Y130_SLICE_X2Y130_DO5),
.O6(CLBLM_R_X3Y130_SLICE_X2Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff08080400)
  ) CLBLM_R_X3Y130_SLICE_X2Y130_CLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLL_L_X2Y130_SLICE_X0Y130_CO5),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(CLBLL_L_X2Y129_SLICE_X0Y129_CO6),
.O5(CLBLM_R_X3Y130_SLICE_X2Y130_CO5),
.O6(CLBLM_R_X3Y130_SLICE_X2Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff7ffff00020050)
  ) CLBLM_R_X3Y130_SLICE_X2Y130_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y130_SLICE_X2Y130_BO5),
.O6(CLBLM_R_X3Y130_SLICE_X2Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0afa0acc000000)
  ) CLBLM_R_X3Y130_SLICE_X2Y130_ALUT (
.I0(CLBLL_L_X4Y124_SLICE_X4Y124_CQ),
.I1(CLBLM_R_X3Y132_SLICE_X2Y132_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y131_SLICE_X2Y131_BQ),
.I4(CLBLM_R_X3Y131_SLICE_X2Y131_CO5),
.I5(1'b1),
.O5(CLBLM_R_X3Y130_SLICE_X2Y130_AO5),
.O6(CLBLM_R_X3Y130_SLICE_X2Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff75ff75ff30ff30)
  ) CLBLM_R_X3Y130_SLICE_X3Y130_DLUT (
.I0(CLBLM_R_X3Y130_SLICE_X3Y130_AO6),
.I1(CLBLL_L_X2Y130_SLICE_X1Y130_BO6),
.I2(LIOB33_X0Y67_IOB_X0Y68_I),
.I3(CLBLL_L_X4Y130_SLICE_X4Y130_DO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y123_SLICE_X2Y123_AQ),
.O5(CLBLM_R_X3Y130_SLICE_X3Y130_DO5),
.O6(CLBLM_R_X3Y130_SLICE_X3Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000010000000)
  ) CLBLM_R_X3Y130_SLICE_X3Y130_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.O5(CLBLM_R_X3Y130_SLICE_X3Y130_CO5),
.O6(CLBLM_R_X3Y130_SLICE_X3Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafefafefffffafe)
  ) CLBLM_R_X3Y130_SLICE_X3Y130_BLUT (
.I0(CLBLM_R_X3Y130_SLICE_X3Y130_DO6),
.I1(CLBLM_R_X3Y130_SLICE_X2Y130_DO6),
.I2(CLBLL_L_X4Y129_SLICE_X4Y129_DO6),
.I3(CLBLM_R_X3Y130_SLICE_X2Y130_CO6),
.I4(CLBLM_R_X7Y129_SLICE_X8Y129_DQ),
.I5(CLBLL_L_X4Y126_SLICE_X4Y126_BO6),
.O5(CLBLM_R_X3Y130_SLICE_X3Y130_BO5),
.O6(CLBLM_R_X3Y130_SLICE_X3Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfffffff21002000)
  ) CLBLM_R_X3Y130_SLICE_X3Y130_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLL_L_X2Y130_SLICE_X0Y130_CO5),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y130_SLICE_X3Y130_AO5),
.O6(CLBLM_R_X3Y130_SLICE_X3Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y131_SLICE_X2Y131_AO6),
.Q(CLBLM_R_X3Y131_SLICE_X2Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y131_SLICE_X2Y131_BO6),
.Q(CLBLM_R_X3Y131_SLICE_X2Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X2Y131_DO5),
.O6(CLBLM_R_X3Y131_SLICE_X2Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha000000080000000)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_CLUT (
.I0(CLBLM_R_X3Y129_SLICE_X2Y129_AQ),
.I1(CLBLM_R_X3Y131_SLICE_X2Y131_AQ),
.I2(CLBLM_R_X3Y132_SLICE_X2Y132_BQ),
.I3(CLBLM_R_X3Y132_SLICE_X2Y132_A5Q),
.I4(CLBLM_R_X3Y123_SLICE_X2Y123_CQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X2Y131_CO5),
.O6(CLBLM_R_X3Y131_SLICE_X2Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff02ff0800020008)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X3Y131_SLICE_X2Y131_BQ),
.I2(CLBLL_L_X2Y118_SLICE_X1Y118_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X3Y131_SLICE_X2Y131_CO5),
.I5(CLBLM_R_X7Y125_SLICE_X9Y125_A5Q),
.O5(CLBLM_R_X3Y131_SLICE_X2Y131_BO5),
.O6(CLBLM_R_X3Y131_SLICE_X2Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ce02cc00ec20)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y131_SLICE_X2Y131_AQ),
.I3(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.I4(CLBLL_L_X2Y118_SLICE_X1Y118_AQ),
.I5(CLBLM_R_X3Y131_SLICE_X2Y131_CO6),
.O5(CLBLM_R_X3Y131_SLICE_X2Y131_AO5),
.O6(CLBLM_R_X3Y131_SLICE_X2Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X3Y131_DO5),
.O6(CLBLM_R_X3Y131_SLICE_X3Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X3Y131_CO5),
.O6(CLBLM_R_X3Y131_SLICE_X3Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X3Y131_BO5),
.O6(CLBLM_R_X3Y131_SLICE_X3Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X3Y131_AO5),
.O6(CLBLM_R_X3Y131_SLICE_X3Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y132_SLICE_X2Y132_CO6),
.Q(CLBLM_R_X3Y132_SLICE_X2Y132_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y132_SLICE_X2Y132_AO6),
.Q(CLBLM_R_X3Y132_SLICE_X2Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y132_SLICE_X2Y132_BO6),
.Q(CLBLM_R_X3Y132_SLICE_X2Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa000000aa000000)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_DLUT (
.I0(CLBLM_R_X3Y123_SLICE_X2Y123_CQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X3Y132_SLICE_X2Y132_A5Q),
.I4(CLBLM_R_X3Y129_SLICE_X2Y129_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y132_SLICE_X2Y132_DO5),
.O6(CLBLM_R_X3Y132_SLICE_X2Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0b1a0a011110000)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X2Y118_SLICE_X1Y118_AQ),
.I2(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.I3(CLBLM_R_X3Y132_SLICE_X2Y132_A5Q),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y132_SLICE_X2Y132_CO5),
.O6(CLBLM_R_X3Y132_SLICE_X2Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff060000000600)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_BLUT (
.I0(CLBLM_R_X3Y132_SLICE_X2Y132_DO6),
.I1(CLBLM_R_X3Y132_SLICE_X2Y132_BQ),
.I2(CLBLL_L_X2Y118_SLICE_X1Y118_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y129_SLICE_X6Y129_BQ),
.O5(CLBLM_R_X3Y132_SLICE_X2Y132_BO5),
.O6(CLBLM_R_X3Y132_SLICE_X2Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888b888888b888)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_ALUT (
.I0(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y132_SLICE_X2Y132_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLL_L_X2Y118_SLICE_X1Y118_AQ),
.I5(CLBLL_L_X2Y132_SLICE_X1Y132_AO6),
.O5(CLBLM_R_X3Y132_SLICE_X2Y132_AO5),
.O6(CLBLM_R_X3Y132_SLICE_X2Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y132_SLICE_X3Y132_DO5),
.O6(CLBLM_R_X3Y132_SLICE_X3Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y132_SLICE_X3Y132_CO5),
.O6(CLBLM_R_X3Y132_SLICE_X3Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y132_SLICE_X3Y132_BO5),
.O6(CLBLM_R_X3Y132_SLICE_X3Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y132_SLICE_X3Y132_AO5),
.O6(CLBLM_R_X3Y132_SLICE_X3Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X6Y116_AO6),
.Q(CLBLM_R_X5Y116_SLICE_X6Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_DO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_CO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_BO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaa0ccccaaa0)
  ) CLBLM_R_X5Y116_SLICE_X6Y116_ALUT (
.I0(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I1(CLBLM_R_X5Y128_SLICE_X7Y128_BQ),
.I2(CLBLM_R_X5Y116_SLICE_X6Y116_AQ),
.I3(CLBLM_L_X8Y119_SLICE_X11Y119_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y116_SLICE_X6Y116_AO5),
.O6(CLBLM_R_X5Y116_SLICE_X6Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X7Y116_AO6),
.Q(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X7Y116_BO6),
.Q(CLBLM_R_X5Y116_SLICE_X7Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y116_SLICE_X7Y116_CO6),
.Q(CLBLM_R_X5Y116_SLICE_X7Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h200000002a000000)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_DLUT (
.I0(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_CQ),
.I2(CLBLL_L_X4Y117_SLICE_X5Y117_BQ),
.I3(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I4(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_DO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00f000c0)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_CLUT (
.I0(CLBLM_R_X5Y116_SLICE_X6Y116_AQ),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_BQ),
.I4(CLBLM_R_X5Y116_SLICE_X7Y116_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_CO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff330033ff300030)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y118_SLICE_X7Y118_DO6),
.I2(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y123_SLICE_X5Y123_AQ),
.I5(CLBLM_R_X5Y116_SLICE_X7Y116_BQ),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_BO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00ffcccc00f0)
  ) CLBLM_R_X5Y116_SLICE_X7Y116_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y117_SLICE_X8Y117_CQ),
.I2(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I3(CLBLM_R_X5Y118_SLICE_X7Y118_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y118_SLICE_X8Y118_AQ),
.O5(CLBLM_R_X5Y116_SLICE_X7Y116_AO5),
.O6(CLBLM_R_X5Y116_SLICE_X7Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y117_SLICE_X6Y117_DO6),
.Q(CLBLM_R_X5Y117_SLICE_X6Y117_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y117_SLICE_X6Y117_AO6),
.Q(CLBLM_R_X5Y117_SLICE_X6Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y117_SLICE_X6Y117_BO6),
.Q(CLBLM_R_X5Y117_SLICE_X6Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y117_SLICE_X6Y117_CO6),
.Q(CLBLM_R_X5Y117_SLICE_X6Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hddd88888000f000f)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y125_SLICE_X6Y125_A5Q),
.I2(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.I3(CLBLM_R_X5Y117_SLICE_X6Y117_A5Q),
.I4(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_DO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f0f3f303000303)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y117_SLICE_X9Y117_CO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.I4(RIOB33_X105Y141_IOB_X1Y142_I),
.I5(CLBLM_R_X5Y126_SLICE_X6Y126_BQ),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_CO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0f0caaaa0000)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_BLUT (
.I0(CLBLM_R_X3Y124_SLICE_X3Y124_CQ),
.I1(CLBLM_R_X5Y117_SLICE_X6Y117_BQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_R_X5Y117_SLICE_X6Y117_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_BO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00facccc00fa)
  ) CLBLM_R_X5Y117_SLICE_X6Y117_ALUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.I1(CLBLM_R_X5Y117_SLICE_X6Y117_BQ),
.I2(CLBLM_R_X5Y117_SLICE_X6Y117_AQ),
.I3(CLBLM_R_X5Y118_SLICE_X7Y118_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y117_SLICE_X6Y117_AO5),
.O6(CLBLM_R_X5Y117_SLICE_X6Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y117_SLICE_X7Y117_AO6),
.Q(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6f6f6f6ff6f6f6f6)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_DLUT (
.I0(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.I1(CLBLM_R_X5Y117_SLICE_X6Y117_A5Q),
.I2(CLBLM_L_X10Y119_SLICE_X13Y119_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_DO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000882200004411)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_CLUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I1(CLBLM_R_X7Y124_SLICE_X8Y124_B5Q),
.I2(1'b1),
.I3(CLBLM_R_X7Y118_SLICE_X8Y118_AQ),
.I4(CLBLM_R_X5Y117_SLICE_X7Y117_DO6),
.I5(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_CO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffb)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_BLUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I1(CLBLM_R_X5Y117_SLICE_X6Y117_DO5),
.I2(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I3(CLBLL_L_X4Y117_SLICE_X5Y117_AQ),
.I4(CLBLM_R_X5Y117_SLICE_X6Y117_AQ),
.I5(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_BO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0032323232)
  ) CLBLM_R_X5Y117_SLICE_X7Y117_ALUT (
.I0(CLBLM_R_X5Y117_SLICE_X6Y117_A5Q),
.I1(CLBLM_R_X5Y118_SLICE_X7Y118_DO6),
.I2(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I3(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y117_SLICE_X7Y117_AO5),
.O6(CLBLM_R_X5Y117_SLICE_X7Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y118_SLICE_X6Y118_CO6),
.Q(CLBLM_R_X5Y118_SLICE_X6Y118_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y118_SLICE_X6Y118_AO6),
.Q(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y118_SLICE_X6Y118_BO6),
.Q(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y118_SLICE_X6Y118_DO6),
.Q(CLBLM_R_X5Y118_SLICE_X6Y118_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00facccc0000)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_DLUT (
.I0(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.I1(CLBLM_R_X7Y120_SLICE_X8Y120_BQ),
.I2(CLBLM_R_X5Y118_SLICE_X6Y118_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_DO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2c0c0ffddffdd)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y119_SLICE_X6Y119_DQ),
.I3(CLBLM_L_X8Y123_SLICE_X11Y123_CQ),
.I4(CLBLM_R_X5Y118_SLICE_X6Y118_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_CO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000fc00fc)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.I2(CLBLM_R_X5Y117_SLICE_X7Y117_AQ),
.I3(CLBLM_R_X5Y118_SLICE_X7Y118_DO6),
.I4(CLBLM_R_X5Y123_SLICE_X7Y123_C5Q),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_BO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf808fa0a0000aaaa)
  ) CLBLM_R_X5Y118_SLICE_X6Y118_ALUT (
.I0(CLBLM_L_X8Y126_SLICE_X11Y126_B5Q),
.I1(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y119_SLICE_X11Y119_BQ),
.I4(RIOB33_X105Y141_IOB_X1Y142_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y118_SLICE_X6Y118_AO5),
.O6(CLBLM_R_X5Y118_SLICE_X6Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y119_SLICE_X6Y119_BO6),
.Q(CLBLM_R_X5Y118_SLICE_X7Y118_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y118_SLICE_X7Y118_AO6),
.Q(CLBLM_R_X5Y118_SLICE_X7Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaaaabaaaa)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_DLUT (
.I0(CLBLL_L_X2Y122_SLICE_X1Y122_CO6),
.I1(CLBLM_R_X3Y127_SLICE_X2Y127_DO6),
.I2(CLBLL_L_X2Y127_SLICE_X0Y127_CO6),
.I3(CLBLL_L_X4Y128_SLICE_X4Y128_AO6),
.I4(CLBLM_R_X5Y118_SLICE_X7Y118_BO5),
.I5(CLBLL_L_X4Y126_SLICE_X4Y126_DO6),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_DO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00fe00ff)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_CLUT (
.I0(CLBLL_L_X4Y128_SLICE_X4Y128_AO6),
.I1(CLBLM_R_X3Y127_SLICE_X2Y127_DO6),
.I2(CLBLL_L_X2Y127_SLICE_X0Y127_CO6),
.I3(CLBLM_R_X3Y124_SLICE_X3Y124_DO6),
.I4(CLBLM_R_X5Y118_SLICE_X7Y118_BO5),
.I5(CLBLL_L_X4Y126_SLICE_X4Y126_DO6),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_CO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5500550000000101)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_BLUT (
.I0(CLBLM_R_X3Y128_SLICE_X3Y128_BO6),
.I1(CLBLM_R_X3Y130_SLICE_X3Y130_BO6),
.I2(CLBLM_R_X3Y128_SLICE_X2Y128_AO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X3Y126_SLICE_X3Y126_AO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_BO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000055505550)
  ) CLBLM_R_X5Y118_SLICE_X7Y118_ALUT (
.I0(CLBLM_R_X5Y118_SLICE_X7Y118_DO6),
.I1(1'b1),
.I2(CLBLM_R_X5Y118_SLICE_X7Y118_AQ),
.I3(CLBLL_L_X4Y117_SLICE_X5Y117_AQ),
.I4(CLBLM_L_X10Y123_SLICE_X12Y123_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y118_SLICE_X7Y118_AO5),
.O6(CLBLM_R_X5Y118_SLICE_X7Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y119_SLICE_X6Y119_AO6),
.Q(CLBLM_R_X5Y119_SLICE_X6Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y119_SLICE_X6Y119_CO6),
.Q(CLBLM_R_X5Y119_SLICE_X6Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y119_SLICE_X6Y119_DO6),
.Q(CLBLM_R_X5Y119_SLICE_X6Y119_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddddd88d8d8d888)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y120_SLICE_X5Y120_AQ),
.I2(CLBLM_R_X5Y119_SLICE_X7Y119_DO6),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I5(CLBLM_R_X5Y119_SLICE_X6Y119_DQ),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_DO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfef0fef00e000e00)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_CLUT (
.I0(CLBLM_R_X5Y116_SLICE_X6Y116_AQ),
.I1(CLBLM_R_X5Y119_SLICE_X6Y119_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y123_SLICE_X3Y123_CQ),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_CO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaea5040f0c0f0c0)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y119_SLICE_X6Y119_DQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X8Y124_SLICE_X10Y124_BQ),
.I4(CLBLL_L_X4Y129_SLICE_X5Y129_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_BO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0d1d1c0c0e2e2)
  ) CLBLM_R_X5Y119_SLICE_X6Y119_ALUT (
.I0(CLBLM_R_X5Y120_SLICE_X6Y120_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y117_SLICE_X6Y117_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X8Y123_SLICE_X11Y123_DO6),
.O5(CLBLM_R_X5Y119_SLICE_X6Y119_AO5),
.O6(CLBLM_R_X5Y119_SLICE_X6Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y119_SLICE_X7Y119_AO6),
.Q(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y119_SLICE_X7Y119_BO6),
.Q(CLBLM_R_X5Y119_SLICE_X7Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y119_SLICE_X7Y119_CO6),
.Q(CLBLM_R_X5Y119_SLICE_X7Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcfcfc0c0c000c)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.I2(CLBLM_R_X3Y123_SLICE_X2Y123_DQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X3Y127_SLICE_X2Y127_DO6),
.I5(CLBLM_L_X8Y123_SLICE_X11Y123_DO6),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_DO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0faa00aa0caa00)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_CLUT (
.I0(CLBLL_L_X4Y126_SLICE_X4Y126_AQ),
.I1(CLBLM_R_X5Y119_SLICE_X7Y119_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I5(CLBLM_L_X8Y119_SLICE_X11Y119_AQ),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_CO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefefef00e0e0e00)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_BLUT (
.I0(CLBLM_R_X5Y118_SLICE_X6Y118_DQ),
.I1(CLBLM_R_X5Y119_SLICE_X7Y119_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLL_L_X2Y122_SLICE_X1Y122_A5Q),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_BO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafc30aaaafc30)
  ) CLBLM_R_X5Y119_SLICE_X7Y119_ALUT (
.I0(CLBLM_R_X5Y116_SLICE_X7Y116_AQ),
.I1(CLBLM_R_X5Y126_SLICE_X7Y126_CO5),
.I2(CLBLM_R_X5Y119_SLICE_X7Y119_AQ),
.I3(CLBLL_L_X4Y122_SLICE_X4Y122_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y119_SLICE_X7Y119_AO5),
.O6(CLBLM_R_X5Y119_SLICE_X7Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X6Y120_AO6),
.Q(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X6Y120_BO6),
.Q(CLBLM_R_X5Y120_SLICE_X6Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X6Y120_CO6),
.Q(CLBLM_R_X5Y120_SLICE_X6Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X6Y120_DO6),
.Q(CLBLM_R_X5Y120_SLICE_X6Y120_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haafaaafa00500050)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_DQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_DO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haabbaaee00110044)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X5Y121_SLICE_X6Y121_CO6),
.I5(CLBLM_R_X3Y120_SLICE_X3Y120_BQ),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_CO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f505f505f000)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.I4(CLBLM_R_X7Y121_SLICE_X8Y121_DO6),
.I5(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_BO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaaaaaffa0a0a0)
  ) CLBLM_R_X5Y120_SLICE_X6Y120_ALUT (
.I0(CLBLM_R_X5Y126_SLICE_X7Y126_CO6),
.I1(1'b1),
.I2(CLBLM_R_X5Y120_SLICE_X6Y120_AQ),
.I3(CLBLM_L_X10Y120_SLICE_X13Y120_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.O5(CLBLM_R_X5Y120_SLICE_X6Y120_AO5),
.O6(CLBLM_R_X5Y120_SLICE_X6Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X7Y120_AO5),
.Q(CLBLM_R_X5Y120_SLICE_X7Y120_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X7Y120_AO6),
.Q(CLBLM_R_X5Y120_SLICE_X7Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y120_SLICE_X7Y120_BO6),
.Q(CLBLM_R_X5Y120_SLICE_X7Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffb1b1ffffa0a0)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_DLUT (
.I0(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X5Y121_SLICE_X6Y121_CO6),
.I3(1'b1),
.I4(CLBLM_R_X3Y123_SLICE_X2Y123_DQ),
.I5(CLBLM_R_X3Y130_SLICE_X3Y130_BO6),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_DO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0066990000996600)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_CLUT (
.I0(CLBLM_R_X5Y121_SLICE_X7Y121_AQ),
.I1(CLBLM_L_X8Y123_SLICE_X11Y123_AQ),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.I5(CLBLL_L_X4Y121_SLICE_X4Y121_DQ),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_CO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hae04fe54ee44ee44)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y120_SLICE_X7Y120_BQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLL_L_X4Y125_SLICE_X4Y125_BQ),
.I4(CLBLM_R_X5Y118_SLICE_X7Y118_BO6),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_BO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00aaaa3333)
  ) CLBLM_R_X5Y120_SLICE_X7Y120_ALUT (
.I0(CLBLM_R_X5Y122_SLICE_X7Y122_BQ),
.I1(CLBLM_R_X3Y119_SLICE_X3Y119_CO6),
.I2(CLBLM_R_X7Y118_SLICE_X9Y118_AQ),
.I3(CLBLM_R_X5Y126_SLICE_X7Y126_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y120_SLICE_X7Y120_AO5),
.O6(CLBLM_R_X5Y120_SLICE_X7Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X6Y121_AO6),
.Q(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X6Y121_BO6),
.Q(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff7fffffffffff)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_DLUT (
.I0(CLBLM_R_X5Y119_SLICE_X6Y119_AQ),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_CQ),
.I2(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.I3(CLBLM_L_X8Y121_SLICE_X10Y121_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X3Y120_SLICE_X3Y120_BQ),
.O5(CLBLM_R_X5Y121_SLICE_X6Y121_DO5),
.O6(CLBLM_R_X5Y121_SLICE_X6Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa8888aaa0aaa0)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_CLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_R_X7Y121_SLICE_X9Y121_B5Q),
.I2(CLBLL_L_X4Y122_SLICE_X4Y122_DQ),
.I3(CLBLM_R_X7Y120_SLICE_X8Y120_BQ),
.I4(CLBLL_L_X4Y121_SLICE_X4Y121_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y121_SLICE_X6Y121_CO5),
.O6(CLBLM_R_X5Y121_SLICE_X6Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5c5c0c0c0c0c5c5)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y125_SLICE_X7Y125_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X5Y119_SLICE_X6Y119_AQ),
.I5(CLBLM_R_X5Y121_SLICE_X7Y121_BO5),
.O5(CLBLM_R_X5Y121_SLICE_X6Y121_BO5),
.O6(CLBLM_R_X5Y121_SLICE_X6Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5500ccccf5f0)
  ) CLBLM_R_X5Y121_SLICE_X6Y121_ALUT (
.I0(CLBLM_R_X5Y121_SLICE_X6Y121_DO6),
.I1(CLBLM_R_X11Y120_SLICE_X15Y120_AQ),
.I2(CLBLM_R_X5Y121_SLICE_X6Y121_AQ),
.I3(CLBLM_R_X5Y121_SLICE_X7Y121_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y121_SLICE_X6Y121_AO5),
.O6(CLBLM_R_X5Y121_SLICE_X6Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y121_SLICE_X7Y121_AO6),
.Q(CLBLM_R_X5Y121_SLICE_X7Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f300ffffff00)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_DLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLL_L_X2Y127_SLICE_X0Y127_CO6),
.I3(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.I4(CLBLM_R_X3Y123_SLICE_X2Y123_DQ),
.I5(CLBLM_R_X5Y121_SLICE_X7Y121_BO5),
.O5(CLBLM_R_X5Y121_SLICE_X7Y121_DO5),
.O6(CLBLM_R_X5Y121_SLICE_X7Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000008000000000)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_CLUT (
.I0(CLBLM_R_X3Y120_SLICE_X2Y120_CQ),
.I1(CLBLL_L_X4Y121_SLICE_X4Y121_DQ),
.I2(CLBLM_L_X8Y123_SLICE_X11Y123_AQ),
.I3(CLBLL_L_X4Y121_SLICE_X5Y121_DO6),
.I4(CLBLM_R_X5Y122_SLICE_X7Y122_DO6),
.I5(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.O5(CLBLM_R_X5Y121_SLICE_X7Y121_CO5),
.O6(CLBLM_R_X5Y121_SLICE_X7Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacacaca0f0f0fff)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_BLUT (
.I0(CLBLM_R_X7Y120_SLICE_X8Y120_AQ),
.I1(CLBLM_L_X8Y122_SLICE_X11Y122_AQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLL_L_X4Y123_SLICE_X5Y123_BQ),
.I4(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y121_SLICE_X7Y121_BO5),
.O6(CLBLM_R_X5Y121_SLICE_X7Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0c5c5caca)
  ) CLBLM_R_X5Y121_SLICE_X7Y121_ALUT (
.I0(CLBLM_L_X8Y121_SLICE_X10Y121_DO5),
.I1(CLBLM_R_X7Y121_SLICE_X9Y121_B5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X8Y123_SLICE_X11Y123_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y121_SLICE_X7Y121_AO5),
.O6(CLBLM_R_X5Y121_SLICE_X7Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X6Y122_AO6),
.Q(CLBLM_R_X5Y122_SLICE_X6Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X6Y122_BO6),
.Q(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X6Y122_CO6),
.Q(CLBLM_R_X5Y122_SLICE_X6Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000080000000)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_DLUT (
.I0(CLBLL_L_X4Y120_SLICE_X5Y120_BQ),
.I1(CLBLL_L_X4Y120_SLICE_X5Y120_AQ),
.I2(CLBLM_R_X5Y123_SLICE_X7Y123_BQ),
.I3(CLBLM_R_X3Y122_SLICE_X2Y122_CQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.O5(CLBLM_R_X5Y122_SLICE_X6Y122_DO5),
.O6(CLBLM_R_X5Y122_SLICE_X6Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccdd0011ccee0022)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_CLUT (
.I0(CLBLM_R_X5Y121_SLICE_X6Y121_CO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.I5(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.O5(CLBLM_R_X5Y122_SLICE_X6Y122_CO5),
.O6(CLBLM_R_X5Y122_SLICE_X6Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f303fc0c)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y122_SLICE_X9Y122_DO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y123_SLICE_X4Y123_BQ),
.I4(CLBLM_R_X7Y120_SLICE_X8Y120_DQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y122_SLICE_X6Y122_BO5),
.O6(CLBLM_R_X5Y122_SLICE_X6Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff7800000f780)
  ) CLBLM_R_X5Y122_SLICE_X6Y122_ALUT (
.I0(CLBLL_L_X4Y125_SLICE_X4Y125_BQ),
.I1(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.I2(CLBLM_R_X5Y122_SLICE_X6Y122_AQ),
.I3(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y121_SLICE_X8Y121_A5Q),
.O5(CLBLM_R_X5Y122_SLICE_X6Y122_AO5),
.O6(CLBLM_R_X5Y122_SLICE_X6Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X7Y122_AO6),
.Q(CLBLM_R_X5Y122_SLICE_X7Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y122_SLICE_X7Y122_BO6),
.Q(CLBLM_R_X5Y122_SLICE_X7Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffff0ffff)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.I4(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.I5(CLBLM_R_X5Y121_SLICE_X7Y121_AQ),
.O5(CLBLM_R_X5Y122_SLICE_X7Y122_DO5),
.O6(CLBLM_R_X5Y122_SLICE_X7Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcf9f90c0c0909)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_CLUT (
.I0(CLBLM_R_X7Y123_SLICE_X9Y123_DO5),
.I1(CLBLM_R_X3Y120_SLICE_X2Y120_BQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(1'b1),
.I4(CLBLL_L_X4Y124_SLICE_X4Y124_DQ),
.I5(CLBLL_L_X4Y123_SLICE_X5Y123_BQ),
.O5(CLBLM_R_X5Y122_SLICE_X7Y122_CO5),
.O6(CLBLM_R_X5Y122_SLICE_X7Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f606f606)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_BLUT (
.I0(CLBLM_L_X8Y124_SLICE_X10Y124_DO6),
.I1(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y121_SLICE_X7Y121_AQ),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y122_SLICE_X7Y122_BO5),
.O6(CLBLM_R_X5Y122_SLICE_X7Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000befa1450)
  ) CLBLM_R_X5Y122_SLICE_X7Y122_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y122_SLICE_X6Y122_DO6),
.I2(CLBLM_R_X5Y122_SLICE_X7Y122_AQ),
.I3(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I4(CLBLM_L_X10Y123_SLICE_X12Y123_BQ),
.I5(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.O5(CLBLM_R_X5Y122_SLICE_X7Y122_AO5),
.O6(CLBLM_R_X5Y122_SLICE_X7Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y123_SLICE_X6Y123_BO5),
.Q(CLBLM_R_X5Y123_SLICE_X6Y123_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y123_SLICE_X6Y123_AO6),
.Q(CLBLM_R_X5Y123_SLICE_X6Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y123_SLICE_X6Y123_BO6),
.Q(CLBLM_R_X5Y123_SLICE_X6Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y123_SLICE_X6Y123_CO6),
.Q(CLBLM_R_X5Y123_SLICE_X6Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800880000000000)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_DLUT (
.I0(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.I1(CLBLM_R_X5Y124_SLICE_X6Y124_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y120_SLICE_X5Y120_A5Q),
.O5(CLBLM_R_X5Y123_SLICE_X6Y123_DO5),
.O6(CLBLM_R_X5Y123_SLICE_X6Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0f5a0a0a0f5a0)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X5Y126_SLICE_X6Y126_DQ),
.I3(CLBLM_L_X8Y122_SLICE_X10Y122_A5Q),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y123_SLICE_X6Y123_CO5),
.O6(CLBLM_R_X5Y123_SLICE_X6Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd1111ce02ce02)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_BLUT (
.I0(RIOB33_X105Y119_IOB_X1Y119_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y123_SLICE_X6Y123_B5Q),
.I3(CLBLM_L_X8Y122_SLICE_X10Y122_A5Q),
.I4(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y123_SLICE_X6Y123_BO5),
.O6(CLBLM_R_X5Y123_SLICE_X6Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00007fff7fff)
  ) CLBLM_R_X5Y123_SLICE_X6Y123_ALUT (
.I0(CLBLM_L_X8Y126_SLICE_X11Y126_B5Q),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X5Y123_SLICE_X6Y123_AQ),
.I3(CLBLM_L_X8Y124_SLICE_X10Y124_B5Q),
.I4(CLBLL_L_X4Y121_SLICE_X5Y121_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y123_SLICE_X6Y123_AO5),
.O6(CLBLM_R_X5Y123_SLICE_X6Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y123_SLICE_X7Y123_CO5),
.Q(CLBLM_R_X5Y123_SLICE_X7Y123_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y123_SLICE_X7Y123_AO6),
.Q(CLBLM_R_X5Y123_SLICE_X7Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y123_SLICE_X7Y123_BO6),
.Q(CLBLM_R_X5Y123_SLICE_X7Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y123_SLICE_X7Y123_CO6),
.Q(CLBLM_R_X5Y123_SLICE_X7Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff7fff7fff)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_DLUT (
.I0(CLBLL_L_X4Y122_SLICE_X4Y122_BQ),
.I1(CLBLM_R_X5Y122_SLICE_X7Y122_BQ),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.I3(CLBLM_R_X7Y125_SLICE_X8Y125_BQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_BQ),
.O5(CLBLM_R_X5Y123_SLICE_X7Y123_DO5),
.O6(CLBLM_R_X5Y123_SLICE_X7Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hae04ae04dddd8888)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y123_SLICE_X7Y123_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X5Y127_SLICE_X7Y127_CQ),
.I4(CLBLL_L_X4Y124_SLICE_X4Y124_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y123_SLICE_X7Y123_CO5),
.O6(CLBLM_R_X5Y123_SLICE_X7Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcfff60f0c0f06)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X5Y123_SLICE_X7Y123_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.I4(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I5(CLBLM_R_X7Y125_SLICE_X8Y125_CQ),
.O5(CLBLM_R_X5Y123_SLICE_X7Y123_BO5),
.O6(CLBLM_R_X5Y123_SLICE_X7Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddd888d8ddd888d8)
  ) CLBLM_R_X5Y123_SLICE_X7Y123_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y122_SLICE_X9Y122_CQ),
.I2(CLBLM_R_X5Y123_SLICE_X7Y123_AQ),
.I3(CLBLM_R_X5Y126_SLICE_X7Y126_CO5),
.I4(CLBLM_R_X5Y119_SLICE_X6Y119_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y123_SLICE_X7Y123_AO5),
.O6(CLBLM_R_X5Y123_SLICE_X7Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X6Y124_DO6),
.Q(CLBLM_R_X5Y124_SLICE_X6Y124_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X6Y124_AO6),
.Q(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X6Y124_BO6),
.Q(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X6Y124_CO6),
.Q(CLBLM_R_X5Y124_SLICE_X6Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888dd88c0c00000)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y124_SLICE_X10Y124_B5Q),
.I2(CLBLM_L_X8Y126_SLICE_X11Y126_B5Q),
.I3(CLBLM_R_X3Y124_SLICE_X3Y124_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y124_SLICE_X6Y124_DO5),
.O6(CLBLM_R_X5Y124_SLICE_X6Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44aa00aa00)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y124_SLICE_X7Y124_C5Q),
.I2(1'b1),
.I3(CLBLM_R_X5Y129_SLICE_X6Y129_AQ),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y124_SLICE_X6Y124_CO5),
.O6(CLBLM_R_X5Y124_SLICE_X6Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f0f0ff00e4e4)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_BLUT (
.I0(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I1(CLBLM_R_X5Y124_SLICE_X6Y124_BQ),
.I2(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.I3(CLBLL_L_X4Y124_SLICE_X5Y124_DQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X5Y124_SLICE_X6Y124_BO5),
.O6(CLBLM_R_X5Y124_SLICE_X6Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888888b8888)
  ) CLBLM_R_X5Y124_SLICE_X6Y124_ALUT (
.I0(CLBLM_R_X5Y126_SLICE_X6Y126_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I3(CLBLM_R_X5Y123_SLICE_X6Y123_BQ),
.I4(RIOB33_X105Y119_IOB_X1Y119_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X5Y124_SLICE_X6Y124_AO5),
.O6(CLBLM_R_X5Y124_SLICE_X6Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X7Y124_CO5),
.Q(CLBLM_R_X5Y124_SLICE_X7Y124_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X7Y124_AO6),
.Q(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X7Y124_BO6),
.Q(CLBLM_R_X5Y124_SLICE_X7Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y124_SLICE_X7Y124_CO6),
.Q(CLBLM_R_X5Y124_SLICE_X7Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000300000000)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y123_SLICE_X7Y123_DO6),
.I2(CLBLM_R_X7Y126_SLICE_X8Y126_DO6),
.I3(CLBLM_R_X3Y124_SLICE_X3Y124_CQ),
.I4(CLBLM_R_X11Y126_SLICE_X14Y126_AQ),
.I5(CLBLM_R_X5Y123_SLICE_X6Y123_DO6),
.O5(CLBLM_R_X5Y124_SLICE_X7Y124_DO5),
.O6(CLBLM_R_X5Y124_SLICE_X7Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2e2e2ccfc0030)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_CLUT (
.I0(CLBLM_R_X7Y127_SLICE_X9Y127_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y122_SLICE_X11Y122_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X3Y123_SLICE_X2Y123_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y124_SLICE_X7Y124_CO5),
.O6(CLBLM_R_X5Y124_SLICE_X7Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefefcfcaaaa0000)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_BLUT (
.I0(CLBLM_L_X10Y123_SLICE_X12Y123_CQ),
.I1(CLBLM_R_X5Y124_SLICE_X7Y124_BQ),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y126_SLICE_X7Y126_CO6),
.O5(CLBLM_R_X5Y124_SLICE_X7Y124_BO5),
.O6(CLBLM_R_X5Y124_SLICE_X7Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aaaaff00fafa)
  ) CLBLM_R_X5Y124_SLICE_X7Y124_ALUT (
.I0(CLBLM_R_X5Y124_SLICE_X7Y124_DO6),
.I1(1'b1),
.I2(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.I3(CLBLM_R_X7Y127_SLICE_X9Y127_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y124_SLICE_X7Y124_AO5),
.O6(CLBLM_R_X5Y124_SLICE_X7Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X6Y125_CO5),
.Q(CLBLM_R_X5Y125_SLICE_X6Y125_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X6Y125_AO6),
.Q(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X6Y125_BO6),
.Q(CLBLM_R_X5Y125_SLICE_X6Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f2f3f0f2f2f0f0f)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_DLUT (
.I0(CLBLL_L_X4Y120_SLICE_X5Y120_BQ),
.I1(CLBLM_R_X3Y122_SLICE_X3Y122_CO6),
.I2(CLBLM_R_X7Y130_SLICE_X8Y130_CO6),
.I3(CLBLM_R_X5Y123_SLICE_X7Y123_BQ),
.I4(CLBLL_L_X4Y120_SLICE_X5Y120_AQ),
.I5(CLBLM_R_X3Y122_SLICE_X2Y122_CQ),
.O5(CLBLM_R_X5Y125_SLICE_X6Y125_DO5),
.O6(CLBLM_R_X5Y125_SLICE_X6Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccc0ccc0f0f0aaaa)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_CLUT (
.I0(CLBLL_L_X4Y123_SLICE_X4Y123_AQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_R_X11Y125_SLICE_X14Y125_BQ),
.I3(CLBLM_L_X8Y122_SLICE_X10Y122_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y125_SLICE_X6Y125_CO5),
.O6(CLBLM_R_X5Y125_SLICE_X6Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0f00cccc0f00)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y130_SLICE_X7Y130_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X8Y124_SLICE_X10Y124_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y125_SLICE_X6Y125_BO5),
.O6(CLBLM_R_X5Y125_SLICE_X6Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc000fcccc0f00)
  ) CLBLM_R_X5Y125_SLICE_X6Y125_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X8Y121_SLICE_X10Y121_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y125_SLICE_X6Y125_CO6),
.O5(CLBLM_R_X5Y125_SLICE_X6Y125_AO5),
.O6(CLBLM_R_X5Y125_SLICE_X6Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X7Y125_AO6),
.Q(CLBLM_R_X5Y125_SLICE_X7Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y125_SLICE_X7Y125_BO6),
.Q(CLBLM_R_X5Y125_SLICE_X7Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff03ff0fff33ffff)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y128_SLICE_X3Y128_BO6),
.I2(CLBLM_R_X3Y130_SLICE_X3Y130_BO6),
.I3(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.I4(CLBLL_L_X2Y127_SLICE_X0Y127_CO6),
.I5(CLBLM_R_X3Y127_SLICE_X2Y127_DO6),
.O5(CLBLM_R_X5Y125_SLICE_X7Y125_DO5),
.O6(CLBLM_R_X5Y125_SLICE_X7Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f01050f0f030f)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_CLUT (
.I0(CLBLM_R_X3Y128_SLICE_X2Y128_AO6),
.I1(CLBLM_R_X3Y126_SLICE_X3Y126_AO6),
.I2(CLBLM_R_X5Y125_SLICE_X6Y125_DO6),
.I3(CLBLL_L_X4Y126_SLICE_X4Y126_DO6),
.I4(CLBLM_R_X5Y125_SLICE_X7Y125_DO6),
.I5(CLBLL_L_X4Y128_SLICE_X4Y128_AO6),
.O5(CLBLM_R_X5Y125_SLICE_X7Y125_CO5),
.O6(CLBLM_R_X5Y125_SLICE_X7Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcffccf0f00000)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y125_SLICE_X7Y125_BQ),
.I2(CLBLM_R_X5Y124_SLICE_X7Y124_BQ),
.I3(CLBLM_R_X3Y120_SLICE_X2Y120_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y126_SLICE_X7Y126_CO6),
.O5(CLBLM_R_X5Y125_SLICE_X7Y125_BO5),
.O6(CLBLM_R_X5Y125_SLICE_X7Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5550ccccfff0)
  ) CLBLM_R_X5Y125_SLICE_X7Y125_ALUT (
.I0(CLBLL_L_X4Y125_SLICE_X4Y125_BQ),
.I1(CLBLM_L_X8Y130_SLICE_X10Y130_BQ),
.I2(CLBLM_R_X5Y125_SLICE_X7Y125_AQ),
.I3(CLBLM_R_X5Y123_SLICE_X7Y123_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.O5(CLBLM_R_X5Y125_SLICE_X7Y125_AO5),
.O6(CLBLM_R_X5Y125_SLICE_X7Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X6Y126_AO6),
.Q(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X6Y126_BO6),
.Q(CLBLM_R_X5Y126_SLICE_X6Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X6Y126_CO6),
.Q(CLBLM_R_X5Y126_SLICE_X6Y126_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X6Y126_DO6),
.Q(CLBLM_R_X5Y126_SLICE_X6Y126_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00ff55fa50)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X5Y126_SLICE_X6Y126_DQ),
.I3(CLBLM_L_X10Y128_SLICE_X12Y128_BQ),
.I4(CLBLM_R_X5Y123_SLICE_X7Y123_C5Q),
.I5(CLBLL_L_X2Y119_SLICE_X1Y119_BO6),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_DO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000fefe00005454)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y126_SLICE_X6Y126_CQ),
.I2(CLBLM_R_X7Y120_SLICE_X8Y120_DQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y126_SLICE_X7Y126_CO6),
.I5(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_CO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00ffaaaa00cc)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_BLUT (
.I0(CLBLM_R_X3Y124_SLICE_X2Y124_BQ),
.I1(CLBLM_R_X5Y126_SLICE_X6Y126_BQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y129_SLICE_X13Y129_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y127_SLICE_X10Y127_BQ),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_BO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa33f0aaaa00f0)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_ALUT (
.I0(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.I3(CLBLL_L_X4Y117_SLICE_X4Y117_AO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y126_SLICE_X4Y126_DO6),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_AO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X7Y126_AO5),
.Q(CLBLM_R_X5Y126_SLICE_X7Y126_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X7Y126_AO6),
.Q(CLBLM_R_X5Y126_SLICE_X7Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X7Y126_BO6),
.Q(CLBLM_R_X5Y126_SLICE_X7Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccddeeeeccddecec)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_DLUT (
.I0(CLBLM_R_X5Y130_SLICE_X7Y130_CO5),
.I1(CLBLM_R_X5Y125_SLICE_X7Y125_CO6),
.I2(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.I3(CLBLM_R_X7Y130_SLICE_X8Y130_CO6),
.I4(CLBLM_R_X5Y120_SLICE_X7Y120_AQ),
.I5(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_DO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h44404444ccc0cccc)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.I4(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_CO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfa0c0afcfa0c0a)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_BLUT (
.I0(CLBLL_L_X2Y122_SLICE_X1Y122_A5Q),
.I1(CLBLM_R_X5Y126_SLICE_X7Y126_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X2Y119_SLICE_X1Y119_BO6),
.I4(CLBLM_L_X10Y128_SLICE_X13Y128_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_BO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0fa0afa0a)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_ALUT (
.I0(CLBLM_R_X5Y128_SLICE_X7Y128_A5Q),
.I1(CLBLL_L_X4Y124_SLICE_X4Y124_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y127_SLICE_X10Y127_AQ),
.I4(RIOB33_X105Y127_IOB_X1Y127_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_AO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X6Y127_AO6),
.Q(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X6Y127_BO6),
.Q(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X6Y127_CO6),
.Q(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000200)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_DLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(CLBLM_R_X5Y126_SLICE_X6Y126_CQ),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_DO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ee44aa00ee44)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y128_SLICE_X7Y128_A5Q),
.I4(CLBLM_R_X5Y126_SLICE_X7Y126_CO5),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_CQ),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_CO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffacac0000acac)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_BLUT (
.I0(CLBLM_R_X5Y121_SLICE_X6Y121_BQ),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.I2(CLBLM_R_X5Y126_SLICE_X7Y126_CO5),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y119_SLICE_X5Y119_AQ),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_BO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fcfcff003030)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y126_SLICE_X7Y126_CO5),
.I2(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.I3(CLBLM_L_X10Y127_SLICE_X13Y127_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y122_SLICE_X6Y122_BQ),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_AO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X7Y127_BO5),
.Q(CLBLM_R_X5Y127_SLICE_X7Y127_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X7Y127_AO6),
.Q(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X7Y127_BO6),
.Q(CLBLM_R_X5Y127_SLICE_X7Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X7Y127_CO6),
.Q(CLBLM_R_X5Y127_SLICE_X7Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000400000)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_DLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(CLBLM_R_X7Y127_SLICE_X8Y127_BQ),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_DO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4e4f5f5a0a0)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y127_SLICE_X7Y127_CQ),
.I2(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y127_SLICE_X7Y127_B5Q),
.I5(CLBLL_L_X2Y119_SLICE_X1Y119_BO6),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_CO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0a0fc0cfc0c)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_BLUT (
.I0(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I1(CLBLL_L_X4Y124_SLICE_X4Y124_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y125_SLICE_X10Y125_DQ),
.I4(CLBLM_L_X10Y127_SLICE_X13Y127_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_BO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0000fc00)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_ALUT (
.I0(CLBLL_L_X4Y122_SLICE_X5Y122_AQ),
.I1(CLBLM_L_X8Y125_SLICE_X10Y125_DQ),
.I2(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_AO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X6Y128_CO6),
.Q(CLBLM_R_X5Y128_SLICE_X6Y128_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X6Y128_AO6),
.Q(CLBLM_R_X5Y128_SLICE_X6Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X6Y128_BO6),
.Q(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X6Y128_DO6),
.Q(CLBLM_R_X5Y128_SLICE_X6Y128_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbaba3030baba3030)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X2Y120_SLICE_X1Y120_BO6),
.I2(CLBLM_R_X5Y128_SLICE_X6Y128_DQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y127_SLICE_X7Y127_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X6Y128_DO5),
.O6(CLBLM_R_X5Y128_SLICE_X6Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbaa330050505050)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X2Y120_SLICE_X1Y120_BO6),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X5Y128_SLICE_X6Y128_A5Q),
.I4(CLBLM_R_X7Y128_SLICE_X9Y128_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X6Y128_CO5),
.O6(CLBLM_R_X5Y128_SLICE_X6Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hacafacaca0a0a0a0)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_BLUT (
.I0(CLBLL_L_X4Y119_SLICE_X5Y119_CQ),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y128_SLICE_X6Y128_BO5),
.O6(CLBLM_R_X5Y128_SLICE_X6Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff222300002223)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_ALUT (
.I0(CLBLM_L_X8Y129_SLICE_X11Y129_B5Q),
.I1(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I2(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.I3(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X2Y121_SLICE_X0Y121_A5Q),
.O5(CLBLM_R_X5Y128_SLICE_X6Y128_AO5),
.O6(CLBLM_R_X5Y128_SLICE_X6Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X7Y128_AO5),
.Q(CLBLM_R_X5Y128_SLICE_X7Y128_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X7Y128_BO5),
.Q(CLBLM_R_X5Y128_SLICE_X7Y128_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X7Y128_AO6),
.Q(CLBLM_R_X5Y128_SLICE_X7Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X7Y128_BO6),
.Q(CLBLM_R_X5Y128_SLICE_X7Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000022332200)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_DLUT (
.I0(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.I1(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.I2(1'b1),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_R_X7Y128_SLICE_X8Y128_CQ),
.I5(CLBLL_L_X2Y130_SLICE_X1Y130_AO6),
.O5(CLBLM_R_X5Y128_SLICE_X7Y128_DO5),
.O6(CLBLM_R_X5Y128_SLICE_X7Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000cc00f0)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y128_SLICE_X8Y128_BQ),
.I2(CLBLM_R_X5Y124_SLICE_X7Y124_BQ),
.I3(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLL_L_X2Y130_SLICE_X1Y130_AO6),
.O5(CLBLM_R_X5Y128_SLICE_X7Y128_CO5),
.O6(CLBLM_R_X5Y128_SLICE_X7Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00ccccff00)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y129_SLICE_X14Y129_AQ),
.I2(CLBLM_R_X3Y129_SLICE_X2Y129_AQ),
.I3(RIOB33_X105Y125_IOB_X1Y126_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X7Y128_BO5),
.O6(CLBLM_R_X5Y128_SLICE_X7Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0a0acacacaca)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_ALUT (
.I0(RIOB33_X105Y143_IOB_X1Y144_I),
.I1(CLBLM_L_X8Y128_SLICE_X11Y128_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLL_L_X2Y119_SLICE_X1Y119_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X7Y128_AO5),
.O6(CLBLM_R_X5Y128_SLICE_X7Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X6Y129_AO6),
.Q(CLBLM_R_X5Y129_SLICE_X6Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X6Y129_BO6),
.Q(CLBLM_R_X5Y129_SLICE_X6Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X6Y129_CO6),
.Q(CLBLM_R_X5Y129_SLICE_X6Y129_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y129_SLICE_X6Y129_DO5),
.O6(CLBLM_R_X5Y129_SLICE_X6Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5e4f5e4a0a0a0a0)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y129_SLICE_X6Y129_CQ),
.I2(CLBLM_R_X5Y123_SLICE_X7Y123_AQ),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_D5Q),
.I4(1'b1),
.I5(CLBLL_L_X2Y119_SLICE_X1Y119_BO6),
.O5(CLBLM_R_X5Y129_SLICE_X6Y129_CO5),
.O6(CLBLM_R_X5Y129_SLICE_X6Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5050cccc5050)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_BLUT (
.I0(CLBLM_R_X7Y131_SLICE_X9Y131_BO5),
.I1(CLBLM_L_X10Y129_SLICE_X13Y129_AQ),
.I2(CLBLM_R_X5Y129_SLICE_X6Y129_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y129_SLICE_X6Y129_BO5),
.O6(CLBLM_R_X5Y129_SLICE_X6Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f0f5f005000500)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_ALUT (
.I0(CLBLM_R_X7Y131_SLICE_X9Y131_BO5),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y129_SLICE_X8Y129_BQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y119_SLICE_X6Y119_CQ),
.O5(CLBLM_R_X5Y129_SLICE_X6Y129_AO5),
.O6(CLBLM_R_X5Y129_SLICE_X6Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X7Y129_AO6),
.Q(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y129_SLICE_X7Y129_DO5),
.O6(CLBLM_R_X5Y129_SLICE_X7Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y129_SLICE_X7Y129_CO5),
.O6(CLBLM_R_X5Y129_SLICE_X7Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0aa0a0a00a20a0a0)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_BLUT (
.I0(CLBLM_R_X5Y128_SLICE_X6Y128_CO5),
.I1(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I2(CLBLM_L_X8Y129_SLICE_X11Y129_B5Q),
.I3(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.I4(CLBLM_R_X5Y130_SLICE_X7Y130_CO5),
.I5(CLBLM_L_X8Y131_SLICE_X10Y131_DO6),
.O5(CLBLM_R_X5Y129_SLICE_X7Y129_BO5),
.O6(CLBLM_R_X5Y129_SLICE_X7Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0c0c0cacfc0c0)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_ALUT (
.I0(CLBLM_R_X7Y130_SLICE_X8Y130_CO6),
.I1(CLBLM_R_X5Y118_SLICE_X6Y118_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_BO6),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.O5(CLBLM_R_X5Y129_SLICE_X7Y129_AO5),
.O6(CLBLM_R_X5Y129_SLICE_X7Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X6Y130_AO6),
.Q(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X6Y130_BO6),
.Q(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_DO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000055005500)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_CLUT (
.I0(CLBLM_R_X5Y130_SLICE_X7Y130_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X7Y129_SLICE_X9Y129_CQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y130_SLICE_X7Y130_BQ),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_CO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fe000ef0f40004)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_BLUT (
.I0(CLBLM_L_X8Y131_SLICE_X10Y131_DO6),
.I1(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X3Y132_SLICE_X2Y132_AQ),
.I5(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_BO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcf00cffffc00fc)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y130_SLICE_X8Y130_CO6),
.I2(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y120_SLICE_X6Y120_BQ),
.I5(CLBLM_R_X5Y130_SLICE_X6Y130_CO6),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_AO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X7Y130_AO6),
.Q(CLBLM_R_X5Y130_SLICE_X7Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X7Y130_BO6),
.Q(CLBLM_R_X5Y130_SLICE_X7Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000040000)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_DLUT (
.I0(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.I1(CLBLM_R_X7Y129_SLICE_X9Y129_CQ),
.I2(CLBLM_R_X5Y130_SLICE_X7Y130_BQ),
.I3(CLBLM_L_X8Y129_SLICE_X11Y129_B5Q),
.I4(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.I5(CLBLM_R_X5Y130_SLICE_X7Y130_AQ),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_DO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5554555500030000)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_CLUT (
.I0(CLBLM_R_X7Y130_SLICE_X8Y130_CO6),
.I1(CLBLM_R_X5Y130_SLICE_X7Y130_AQ),
.I2(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.I3(CLBLM_R_X5Y130_SLICE_X7Y130_BQ),
.I4(CLBLM_R_X7Y129_SLICE_X9Y129_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_CO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf303fc0cf000f000)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y129_SLICE_X9Y129_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y128_SLICE_X8Y128_BQ),
.I4(CLBLM_R_X5Y130_SLICE_X7Y130_BQ),
.I5(CLBLM_R_X5Y130_SLICE_X7Y130_CO6),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_BO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50be14aa00aa00)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y129_SLICE_X9Y129_CQ),
.I2(CLBLM_R_X5Y130_SLICE_X7Y130_AQ),
.I3(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.I4(CLBLM_R_X5Y130_SLICE_X7Y130_BQ),
.I5(CLBLM_R_X5Y130_SLICE_X7Y130_CO6),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_AO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_DO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_CO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_BO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0002fffd11111111)
  ) CLBLM_R_X7Y115_SLICE_X8Y115_ALUT (
.I0(CLBLL_L_X4Y117_SLICE_X5Y117_BQ),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_CQ),
.I2(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I3(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I4(CLBLM_R_X5Y119_SLICE_X6Y119_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X8Y115_AO5),
.O6(CLBLM_R_X7Y115_SLICE_X8Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_DO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_CO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0022ffdd0000ffff)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_BLUT (
.I0(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I1(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y116_SLICE_X7Y116_CQ),
.I4(CLBLM_L_X10Y119_SLICE_X12Y119_CQ),
.I5(CLBLL_L_X4Y117_SLICE_X5Y117_BQ),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_BO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f4b0f0f55005500)
  ) CLBLM_R_X7Y115_SLICE_X9Y115_ALUT (
.I0(CLBLL_L_X4Y117_SLICE_X5Y117_BQ),
.I1(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I2(CLBLM_R_X5Y116_SLICE_X6Y116_AQ),
.I3(CLBLM_R_X5Y116_SLICE_X7Y116_CQ),
.I4(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y115_SLICE_X9Y115_AO5),
.O6(CLBLM_R_X7Y115_SLICE_X9Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y116_SLICE_X8Y116_AO6),
.Q(CLBLM_R_X7Y116_SLICE_X8Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000505000f0505)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_DLUT (
.I0(CLBLM_R_X7Y118_SLICE_X8Y118_C5Q),
.I1(1'b1),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_AQ),
.I3(CLBLM_R_X7Y119_SLICE_X8Y119_CQ),
.I4(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I5(CLBLM_L_X8Y118_SLICE_X11Y118_CO6),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_DO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h05050909000f000f)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_CLUT (
.I0(CLBLM_R_X5Y116_SLICE_X6Y116_AQ),
.I1(CLBLM_R_X7Y115_SLICE_X8Y115_AO5),
.I2(CLBLM_R_X7Y117_SLICE_X8Y117_DQ),
.I3(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.I4(CLBLM_R_X7Y116_SLICE_X8Y116_BO5),
.I5(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_CO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h333333630fff0fff)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_BLUT (
.I0(CLBLL_L_X4Y117_SLICE_X5Y117_BQ),
.I1(CLBLM_L_X8Y119_SLICE_X11Y119_BQ),
.I2(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I3(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I4(CLBLM_R_X5Y116_SLICE_X7Y116_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_BO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5555cccc0055)
  ) CLBLM_R_X7Y116_SLICE_X8Y116_ALUT (
.I0(CLBLM_R_X7Y116_SLICE_X8Y116_DO6),
.I1(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.I2(1'b1),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.O5(CLBLM_R_X7Y116_SLICE_X8Y116_AO5),
.O6(CLBLM_R_X7Y116_SLICE_X8Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y116_SLICE_X9Y116_AO6),
.Q(CLBLM_R_X7Y116_SLICE_X9Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y116_SLICE_X9Y116_BO6),
.Q(CLBLM_R_X7Y116_SLICE_X9Y116_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5500550000005555)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_DLUT (
.I0(CLBLM_R_X7Y116_SLICE_X9Y116_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X7Y116_SLICE_X8Y116_BO6),
.I4(CLBLM_R_X7Y124_SLICE_X8Y124_B5Q),
.I5(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_DO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0f00f66f066)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_CLUT (
.I0(CLBLM_R_X7Y115_SLICE_X8Y115_AO6),
.I1(CLBLM_R_X7Y117_SLICE_X9Y117_AO6),
.I2(CLBLM_L_X10Y120_SLICE_X13Y120_A5Q),
.I3(CLBLM_R_X3Y124_SLICE_X3Y124_DO6),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.I5(CLBLM_R_X3Y126_SLICE_X2Y126_BO6),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_CO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf505f505f101f101)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_BLUT (
.I0(CLBLM_R_X7Y116_SLICE_X9Y116_DO6),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y119_SLICE_X10Y119_BQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_BO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0050505050)
  ) CLBLM_R_X7Y116_SLICE_X9Y116_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(CLBLM_R_X7Y116_SLICE_X9Y116_AQ),
.I3(CLBLM_R_X7Y118_SLICE_X8Y118_C5Q),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y116_SLICE_X9Y116_AO5),
.O6(CLBLM_R_X7Y116_SLICE_X9Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X8Y117_AO6),
.Q(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X8Y117_BO6),
.Q(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X8Y117_CO6),
.Q(CLBLM_R_X7Y117_SLICE_X8Y117_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y117_SLICE_X8Y117_DO6),
.Q(CLBLM_R_X7Y117_SLICE_X8Y117_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbabbbab11011101)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y116_SLICE_X8Y116_CO6),
.I2(RIOB33_X105Y141_IOB_X1Y142_I),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y122_SLICE_X3Y122_AQ),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_DO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaaafaf05000505)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X7Y117_SLICE_X9Y117_BO6),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.I4(RIOB33_X105Y141_IOB_X1Y142_I),
.I5(CLBLM_R_X7Y123_SLICE_X9Y123_A5Q),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_CO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0aca0a3a0a0a0a0)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_BLUT (
.I0(CLBLM_L_X10Y118_SLICE_X12Y118_AQ),
.I1(CLBLM_L_X8Y117_SLICE_X10Y117_CO5),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_BQ),
.I4(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_BO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff100010ff100010)
  ) CLBLM_R_X7Y117_SLICE_X8Y117_ALUT (
.I0(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y116_SLICE_X9Y116_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y117_SLICE_X8Y117_AO5),
.O6(CLBLM_R_X7Y117_SLICE_X8Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000020028008)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_DLUT (
.I0(CLBLM_R_X5Y117_SLICE_X7Y117_CO6),
.I1(CLBLM_R_X7Y118_SLICE_X9Y118_DO6),
.I2(CLBLM_R_X5Y116_SLICE_X7Y116_BQ),
.I3(CLBLM_L_X10Y120_SLICE_X13Y120_A5Q),
.I4(CLBLM_L_X10Y121_SLICE_X12Y121_CQ),
.I5(CLBLM_L_X8Y117_SLICE_X11Y117_CO6),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_DO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00080a02050d0f07)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_CLUT (
.I0(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I1(CLBLM_R_X7Y115_SLICE_X9Y115_AO5),
.I2(CLBLM_R_X5Y117_SLICE_X6Y117_CQ),
.I3(CLBLM_R_X7Y117_SLICE_X9Y117_AO5),
.I4(CLBLM_R_X7Y118_SLICE_X8Y118_DQ),
.I5(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_CO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033030322110303)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_BLUT (
.I0(CLBLM_L_X8Y117_SLICE_X10Y117_DO6),
.I1(CLBLM_R_X7Y117_SLICE_X8Y117_CQ),
.I2(CLBLL_L_X4Y120_SLICE_X4Y120_C5Q),
.I3(CLBLM_L_X10Y119_SLICE_X12Y119_CQ),
.I4(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I5(CLBLM_R_X7Y117_SLICE_X9Y117_AO5),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_BO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555955f0fff0ff)
  ) CLBLM_R_X7Y117_SLICE_X9Y117_ALUT (
.I0(CLBLM_R_X7Y118_SLICE_X8Y118_DQ),
.I1(CLBLM_R_X5Y116_SLICE_X7Y116_CQ),
.I2(CLBLM_L_X10Y117_SLICE_X12Y117_AQ),
.I3(CLBLM_R_X7Y117_SLICE_X8Y117_BQ),
.I4(CLBLL_L_X4Y117_SLICE_X5Y117_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y117_SLICE_X9Y117_AO5),
.O6(CLBLM_R_X7Y117_SLICE_X9Y117_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y118_SLICE_X8Y118_CO5),
.Q(CLBLM_R_X7Y118_SLICE_X8Y118_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y118_SLICE_X8Y118_AO6),
.Q(CLBLM_R_X7Y118_SLICE_X8Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y118_SLICE_X8Y118_BO6),
.Q(CLBLM_R_X7Y118_SLICE_X8Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y118_SLICE_X8Y118_CO6),
.Q(CLBLM_R_X7Y118_SLICE_X8Y118_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y118_SLICE_X8Y118_DO6),
.Q(CLBLM_R_X7Y118_SLICE_X8Y118_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55fa50aa00aa00)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X7Y118_SLICE_X8Y118_DQ),
.I3(CLBLM_R_X5Y118_SLICE_X7Y118_A5Q),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_DQ),
.I5(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.O5(CLBLM_R_X7Y118_SLICE_X8Y118_DO5),
.O6(CLBLM_R_X7Y118_SLICE_X8Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500e4e4e4e4)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y118_SLICE_X7Y118_A5Q),
.I2(CLBLM_R_X7Y116_SLICE_X8Y116_AQ),
.I3(CLBLM_R_X5Y120_SLICE_X7Y120_CO6),
.I4(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y118_SLICE_X8Y118_CO5),
.O6(CLBLM_R_X7Y118_SLICE_X8Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ffe0ef000f404)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_BLUT (
.I0(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I1(CLBLM_R_X7Y118_SLICE_X8Y118_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y119_SLICE_X7Y119_BQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLL_L_X4Y118_SLICE_X4Y118_AQ),
.O5(CLBLM_R_X7Y118_SLICE_X8Y118_BO5),
.O6(CLBLM_R_X7Y118_SLICE_X8Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0a0a3a3a0a0)
  ) CLBLM_R_X7Y118_SLICE_X8Y118_ALUT (
.I0(CLBLM_R_X7Y129_SLICE_X8Y129_DQ),
.I1(CLBLM_R_X7Y118_SLICE_X9Y118_DO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X3Y125_SLICE_X2Y125_BO6),
.I5(CLBLM_R_X7Y118_SLICE_X8Y118_AQ),
.O5(CLBLM_R_X7Y118_SLICE_X8Y118_AO5),
.O6(CLBLM_R_X7Y118_SLICE_X8Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y118_SLICE_X9Y118_AO6),
.Q(CLBLM_R_X7Y118_SLICE_X9Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa005100aaff51ff)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_DLUT (
.I0(CLBLM_L_X8Y118_SLICE_X11Y118_BQ),
.I1(CLBLM_L_X8Y118_SLICE_X11Y118_DO6),
.I2(CLBLM_R_X5Y117_SLICE_X7Y117_BO6),
.I3(CLBLM_R_X3Y119_SLICE_X3Y119_BO5),
.I4(CLBLM_R_X5Y118_SLICE_X7Y118_AQ),
.I5(CLBLM_L_X10Y121_SLICE_X12Y121_CQ),
.O5(CLBLM_R_X7Y118_SLICE_X9Y118_DO5),
.O6(CLBLM_R_X7Y118_SLICE_X9Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffdffffffff)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_CLUT (
.I0(CLBLM_R_X3Y126_SLICE_X3Y126_AO6),
.I1(CLBLM_R_X7Y128_SLICE_X9Y128_BO6),
.I2(CLBLL_L_X4Y126_SLICE_X4Y126_DO6),
.I3(CLBLM_R_X3Y128_SLICE_X2Y128_AO6),
.I4(CLBLL_L_X4Y128_SLICE_X4Y128_AO6),
.I5(CLBLM_R_X5Y118_SLICE_X7Y118_BO6),
.O5(CLBLM_R_X7Y118_SLICE_X9Y118_CO5),
.O6(CLBLM_R_X7Y118_SLICE_X9Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00003333fffffffa)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_BLUT (
.I0(CLBLL_L_X2Y127_SLICE_X0Y127_CO6),
.I1(CLBLM_R_X7Y128_SLICE_X9Y128_BO6),
.I2(CLBLL_L_X4Y128_SLICE_X4Y128_AO6),
.I3(CLBLL_L_X4Y126_SLICE_X4Y126_DO6),
.I4(CLBLM_R_X3Y127_SLICE_X2Y127_DO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y118_SLICE_X9Y118_BO5),
.O6(CLBLM_R_X7Y118_SLICE_X9Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafc00aaaafc00)
  ) CLBLM_R_X7Y118_SLICE_X9Y118_ALUT (
.I0(CLBLM_R_X7Y125_SLICE_X9Y125_DQ),
.I1(CLBLM_L_X8Y116_SLICE_X10Y116_BQ),
.I2(CLBLM_R_X7Y118_SLICE_X9Y118_AQ),
.I3(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y118_SLICE_X9Y118_AO5),
.O6(CLBLM_R_X7Y118_SLICE_X9Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X8Y119_AO6),
.Q(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X8Y119_BO6),
.Q(CLBLM_R_X7Y119_SLICE_X8Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X8Y119_CO6),
.Q(CLBLM_R_X7Y119_SLICE_X8Y119_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X8Y119_DO6),
.Q(CLBLM_R_X7Y119_SLICE_X8Y119_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaafc00fc00)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_DLUT (
.I0(CLBLM_R_X5Y124_SLICE_X7Y124_AQ),
.I1(CLBLM_R_X7Y119_SLICE_X8Y119_CQ),
.I2(CLBLM_R_X7Y119_SLICE_X8Y119_DQ),
.I3(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_DO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0a0af8f80808)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_CLUT (
.I0(CLBLM_R_X5Y118_SLICE_X7Y118_CO6),
.I1(CLBLM_R_X7Y119_SLICE_X8Y119_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X7Y125_SLICE_X8Y125_DQ),
.I5(CLBLM_L_X10Y119_SLICE_X12Y119_DQ),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_CO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf055f044f000f000)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X7Y119_SLICE_X8Y119_BQ),
.I2(CLBLM_R_X5Y119_SLICE_X6Y119_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y116_SLICE_X9Y116_BQ),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_BO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfaccfaccfacc00)
  ) CLBLM_R_X7Y119_SLICE_X8Y119_ALUT (
.I0(CLBLM_R_X7Y123_SLICE_X8Y123_B5Q),
.I1(CLBLM_R_X7Y119_SLICE_X8Y119_BQ),
.I2(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.O5(CLBLM_R_X7Y119_SLICE_X8Y119_AO5),
.O6(CLBLM_R_X7Y119_SLICE_X8Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X9Y119_AO6),
.Q(CLBLM_R_X7Y119_SLICE_X9Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y119_SLICE_X9Y119_BO6),
.Q(CLBLM_R_X7Y119_SLICE_X9Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001100000011)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_DLUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I1(CLBLM_L_X8Y118_SLICE_X10Y118_CQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y119_SLICE_X5Y119_BQ),
.I4(CLBLM_R_X3Y119_SLICE_X3Y119_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_DO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddfffc00000000)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_CLUT (
.I0(CLBLM_L_X8Y118_SLICE_X10Y118_BQ),
.I1(CLBLM_L_X10Y122_SLICE_X12Y122_AQ),
.I2(CLBLL_L_X2Y127_SLICE_X0Y127_CO6),
.I3(CLBLM_R_X7Y128_SLICE_X9Y128_BO6),
.I4(CLBLM_R_X7Y119_SLICE_X9Y119_DO6),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_CO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0afaca0a0a0a0)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_BLUT (
.I0(CLBLM_L_X8Y118_SLICE_X10Y118_CQ),
.I1(CLBLM_R_X7Y119_SLICE_X9Y119_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y119_SLICE_X7Y119_DO6),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_BO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f1f4f401010404)
  ) CLBLM_R_X7Y119_SLICE_X9Y119_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y124_SLICE_X13Y124_DQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X5Y119_SLICE_X6Y119_BO5),
.I5(CLBLL_L_X4Y119_SLICE_X5Y119_BQ),
.O5(CLBLM_R_X7Y119_SLICE_X9Y119_AO5),
.O6(CLBLM_R_X7Y119_SLICE_X9Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y120_SLICE_X8Y120_AO6),
.Q(CLBLM_R_X7Y120_SLICE_X8Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y120_SLICE_X8Y120_BO6),
.Q(CLBLM_R_X7Y120_SLICE_X8Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y120_SLICE_X8Y120_CO6),
.Q(CLBLM_R_X7Y120_SLICE_X8Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y120_SLICE_X8Y120_DO6),
.Q(CLBLM_R_X7Y120_SLICE_X8Y120_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0a3aca3ac)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_DLUT (
.I0(CLBLM_R_X7Y118_SLICE_X8Y118_BQ),
.I1(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y122_SLICE_X8Y122_CO6),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_DO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5e4a0a0a0e4)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y120_SLICE_X8Y120_CQ),
.I2(CLBLM_R_X7Y128_SLICE_X8Y128_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I5(CLBLM_R_X7Y119_SLICE_X8Y119_BQ),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_CO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ffa0afc0cf808)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_BLUT (
.I0(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I1(CLBLM_R_X7Y120_SLICE_X8Y120_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y128_SLICE_X11Y128_BQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X7Y122_SLICE_X8Y122_CO6),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_BO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fcfcff00a8a8)
  ) CLBLM_R_X7Y120_SLICE_X8Y120_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X7Y122_SLICE_X9Y122_DO6),
.I2(CLBLM_R_X7Y120_SLICE_X8Y120_AQ),
.I3(CLBLM_R_X7Y120_SLICE_X8Y120_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.O5(CLBLM_R_X7Y120_SLICE_X8Y120_AO5),
.O6(CLBLM_R_X7Y120_SLICE_X8Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0000ffcc0033ff)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y127_SLICE_X2Y127_DO6),
.I2(1'b1),
.I3(CLBLM_R_X11Y122_SLICE_X14Y122_BQ),
.I4(CLBLM_R_X5Y119_SLICE_X7Y119_BQ),
.I5(CLBLM_R_X7Y128_SLICE_X9Y128_BO6),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_DO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffffffefffe)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I2(CLBLM_R_X3Y123_SLICE_X2Y123_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_CO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffa2ff22)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_BLUT (
.I0(CLBLL_L_X4Y126_SLICE_X4Y126_DO6),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLL_L_X4Y118_SLICE_X5Y118_AQ),
.I3(CLBLM_L_X8Y121_SLICE_X11Y121_DO5),
.I4(CLBLM_R_X5Y124_SLICE_X6Y124_CQ),
.I5(CLBLM_R_X7Y120_SLICE_X9Y120_CO6),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_BO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ecfceccc)
  ) CLBLM_R_X7Y120_SLICE_X9Y120_ALUT (
.I0(CLBLM_L_X8Y122_SLICE_X11Y122_AQ),
.I1(CLBLM_L_X8Y121_SLICE_X11Y121_DO5),
.I2(CLBLM_R_X3Y126_SLICE_X3Y126_AO6),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X7Y120_SLICE_X8Y120_AQ),
.I5(CLBLM_R_X7Y120_SLICE_X9Y120_CO6),
.O5(CLBLM_R_X7Y120_SLICE_X9Y120_AO5),
.O6(CLBLM_R_X7Y120_SLICE_X9Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y121_SLICE_X10Y121_AO6),
.Q(CLBLM_R_X7Y121_SLICE_X8Y121_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X8Y121_AO6),
.Q(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X8Y121_BO6),
.Q(CLBLM_R_X7Y121_SLICE_X8Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f000fb00f044)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_DLUT (
.I0(CLBLM_L_X8Y124_SLICE_X10Y124_AQ),
.I1(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.I2(CLBLL_L_X4Y122_SLICE_X5Y122_DQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X7Y127_SLICE_X8Y127_CQ),
.I5(CLBLM_R_X7Y124_SLICE_X8Y124_CO5),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_DO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f2f0f0dfffd)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_CLUT (
.I0(CLBLM_L_X8Y124_SLICE_X10Y124_AQ),
.I1(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X7Y124_SLICE_X8Y124_CO5),
.I4(CLBLM_L_X8Y122_SLICE_X11Y122_AQ),
.I5(CLBLM_R_X5Y120_SLICE_X6Y120_DQ),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_CO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000c0cff000303)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y125_SLICE_X8Y125_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X11Y122_SLICE_X14Y122_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y121_SLICE_X8Y121_CO6),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_BO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0c0aaaaffcc)
  ) CLBLM_R_X7Y121_SLICE_X8Y121_ALUT (
.I0(CLBLM_R_X3Y126_SLICE_X2Y126_A5Q),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y121_SLICE_X8Y121_CO6),
.O5(CLBLM_R_X7Y121_SLICE_X8Y121_AO5),
.O6(CLBLM_R_X7Y121_SLICE_X8Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X9Y121_BO5),
.Q(CLBLM_R_X7Y121_SLICE_X9Y121_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X9Y121_AO6),
.Q(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y121_SLICE_X9Y121_BO6),
.Q(CLBLM_R_X7Y121_SLICE_X9Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00c000cf00c000)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y121_SLICE_X6Y121_CO5),
.I2(CLBLM_R_X3Y123_SLICE_X2Y123_DQ),
.I3(CLBLM_L_X8Y118_SLICE_X10Y118_AO5),
.I4(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.I5(CLBLM_R_X5Y118_SLICE_X7Y118_BO6),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_DO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_CLUT (
.I0(CLBLM_L_X8Y119_SLICE_X10Y119_BQ),
.I1(CLBLM_R_X5Y120_SLICE_X6Y120_DQ),
.I2(CLBLM_R_X5Y123_SLICE_X7Y123_CQ),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_B5Q),
.I4(CLBLM_R_X7Y116_SLICE_X9Y116_AQ),
.I5(CLBLM_L_X8Y123_SLICE_X11Y123_C5Q),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_CO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacacacfa0af000)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_BLUT (
.I0(CLBLM_R_X5Y123_SLICE_X6Y123_CQ),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_A5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y121_SLICE_X14Y121_AQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_BO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d88888d8d8)
  ) CLBLM_R_X7Y121_SLICE_X9Y121_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y123_SLICE_X8Y123_B5Q),
.I2(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.O5(CLBLM_R_X7Y121_SLICE_X9Y121_AO5),
.O6(CLBLM_R_X7Y121_SLICE_X9Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X8Y122_AO6),
.Q(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X8Y122_BO6),
.Q(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f000f004b000f)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_DLUT (
.I0(CLBLM_L_X8Y124_SLICE_X10Y124_AQ),
.I1(CLBLL_L_X4Y124_SLICE_X4Y124_DQ),
.I2(CLBLM_L_X8Y121_SLICE_X11Y121_CQ),
.I3(CLBLM_R_X3Y122_SLICE_X2Y122_A5Q),
.I4(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.I5(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_DO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf077f088f0fff000)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_CLUT (
.I0(CLBLM_L_X8Y124_SLICE_X10Y124_AQ),
.I1(CLBLM_R_X7Y124_SLICE_X8Y124_CO6),
.I2(CLBLM_R_X5Y124_SLICE_X6Y124_CQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X5Y123_SLICE_X7Y123_CQ),
.I5(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_CO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5050cccca0a0)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_BLUT (
.I0(CLBLM_R_X7Y123_SLICE_X8Y123_DO6),
.I1(CLBLM_R_X5Y125_SLICE_X6Y125_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y119_SLICE_X9Y119_CO6),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_BO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888dd888888dd8)
  ) CLBLM_R_X7Y122_SLICE_X8Y122_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y122_SLICE_X15Y122_AQ),
.I2(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I3(CLBLM_R_X5Y122_SLICE_X6Y122_DO6),
.I4(CLBLM_R_X7Y119_SLICE_X8Y119_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y122_SLICE_X8Y122_AO5),
.O6(CLBLM_R_X7Y122_SLICE_X8Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X9Y122_AO6),
.Q(CLBLM_R_X7Y122_SLICE_X9Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X9Y122_BO6),
.Q(CLBLM_R_X7Y122_SLICE_X9Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y122_SLICE_X9Y122_CO6),
.Q(CLBLM_R_X7Y122_SLICE_X9Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f000f070f080)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_DLUT (
.I0(CLBLM_L_X8Y124_SLICE_X10Y124_AQ),
.I1(CLBLM_R_X7Y124_SLICE_X8Y124_CO6),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X10Y126_SLICE_X12Y126_CQ),
.I4(CLBLM_L_X8Y123_SLICE_X11Y123_C5Q),
.I5(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_DO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0b1a0b1a0)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y122_SLICE_X10Y122_BO6),
.I2(CLBLM_R_X5Y128_SLICE_X7Y128_B5Q),
.I3(CLBLM_L_X10Y122_SLICE_X12Y122_AQ),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_CO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00044f0f00000)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y123_SLICE_X10Y123_BQ),
.I2(CLBLM_R_X7Y121_SLICE_X9Y121_AQ),
.I3(CLBLM_L_X8Y122_SLICE_X10Y122_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y122_SLICE_X12Y122_AQ),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_BO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00facccc0000)
  ) CLBLM_R_X7Y122_SLICE_X9Y122_ALUT (
.I0(CLBLM_R_X7Y117_SLICE_X8Y117_CQ),
.I1(CLBLM_L_X8Y123_SLICE_X10Y123_BQ),
.I2(CLBLM_R_X7Y122_SLICE_X9Y122_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.O5(CLBLM_R_X7Y122_SLICE_X9Y122_AO5),
.O6(CLBLM_R_X7Y122_SLICE_X9Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X8Y123_BO5),
.Q(CLBLM_R_X7Y123_SLICE_X8Y123_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X8Y123_AO6),
.Q(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X8Y123_BO6),
.Q(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3cc3c3c3c33c3c)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y124_SLICE_X6Y124_A5Q),
.I2(CLBLM_R_X11Y126_SLICE_X14Y126_AQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y127_SLICE_X11Y127_CQ),
.I5(CLBLM_R_X7Y122_SLICE_X8Y122_BQ),
.O5(CLBLM_R_X7Y123_SLICE_X8Y123_DO5),
.O6(CLBLM_R_X7Y123_SLICE_X8Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0c0f0c0f0c0)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_CLUT (
.I0(CLBLM_L_X8Y120_SLICE_X10Y120_AQ),
.I1(CLBLL_L_X4Y122_SLICE_X4Y122_DQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X7Y123_SLICE_X9Y123_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y123_SLICE_X8Y123_CO5),
.O6(CLBLM_R_X7Y123_SLICE_X8Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf202f202fff50f05)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_BLUT (
.I0(RIOB33_X105Y119_IOB_X1Y119_I),
.I1(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y123_SLICE_X6Y123_BQ),
.I4(CLBLM_R_X3Y121_SLICE_X2Y121_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y123_SLICE_X8Y123_BO5),
.O6(CLBLM_R_X7Y123_SLICE_X8Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00c0aaaa00c0)
  ) CLBLM_R_X7Y123_SLICE_X8Y123_ALUT (
.I0(CLBLM_R_X5Y122_SLICE_X6Y122_CQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.I3(CLBLM_R_X5Y124_SLICE_X7Y124_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y123_SLICE_X8Y123_AO5),
.O6(CLBLM_R_X7Y123_SLICE_X8Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X9Y123_AO5),
.Q(CLBLM_R_X7Y123_SLICE_X9Y123_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X9Y123_AO6),
.Q(CLBLM_R_X7Y123_SLICE_X9Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X9Y123_BO6),
.Q(CLBLM_R_X7Y123_SLICE_X9Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y123_SLICE_X9Y123_CO6),
.Q(CLBLM_R_X7Y123_SLICE_X9Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff04fbfffff5f5)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_DLUT (
.I0(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.I1(CLBLL_L_X4Y124_SLICE_X4Y124_DQ),
.I2(CLBLM_L_X8Y124_SLICE_X10Y124_AQ),
.I3(CLBLM_R_X7Y123_SLICE_X9Y123_AQ),
.I4(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y123_SLICE_X9Y123_DO5),
.O6(CLBLM_R_X7Y123_SLICE_X9Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffe4e4ffffe4a0)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y123_SLICE_X9Y123_CQ),
.I2(CLBLL_L_X4Y119_SLICE_X4Y119_BQ),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I4(CLBLM_R_X7Y121_SLICE_X9Y121_DO6),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X7Y123_SLICE_X9Y123_CO5),
.O6(CLBLM_R_X7Y123_SLICE_X9Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0aca0afafacac)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_BLUT (
.I0(CLBLM_L_X10Y120_SLICE_X13Y120_CQ),
.I1(CLBLM_R_X7Y123_SLICE_X9Y123_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y120_SLICE_X14Y120_DO6),
.I4(CLBLL_L_X4Y120_SLICE_X5Y120_BQ),
.I5(CLBLM_R_X7Y123_SLICE_X9Y123_A5Q),
.O5(CLBLM_R_X7Y123_SLICE_X9Y123_BO5),
.O6(CLBLM_R_X7Y123_SLICE_X9Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff002222aaaaf0f0)
  ) CLBLM_R_X7Y123_SLICE_X9Y123_ALUT (
.I0(CLBLM_R_X7Y123_SLICE_X9Y123_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLL_L_X4Y121_SLICE_X5Y121_AQ),
.I3(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y123_SLICE_X9Y123_AO5),
.O6(CLBLM_R_X7Y123_SLICE_X9Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X8Y124_BO5),
.Q(CLBLM_R_X7Y124_SLICE_X8Y124_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X8Y124_AO6),
.Q(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X8Y124_BO6),
.Q(CLBLM_R_X7Y124_SLICE_X8Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff02c402ff00cc00)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_DLUT (
.I0(CLBLM_L_X8Y124_SLICE_X10Y124_AQ),
.I1(CLBLM_R_X7Y129_SLICE_X9Y129_DQ),
.I2(CLBLM_R_X7Y124_SLICE_X8Y124_CO5),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLL_L_X4Y122_SLICE_X4Y122_DQ),
.I5(CLBLM_L_X8Y124_SLICE_X11Y124_AQ),
.O5(CLBLM_R_X7Y124_SLICE_X8Y124_DO5),
.O6(CLBLM_R_X7Y124_SLICE_X8Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00550055aaffaaff)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_CLUT (
.I0(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X4Y124_SLICE_X4Y124_DQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y124_SLICE_X8Y124_CO5),
.O6(CLBLM_R_X7Y124_SLICE_X8Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0f0ccccff00)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_BLUT (
.I0(CLBLM_L_X8Y128_SLICE_X10Y128_AQ),
.I1(CLBLM_R_X3Y125_SLICE_X3Y125_BQ),
.I2(CLBLM_L_X10Y124_SLICE_X13Y124_A5Q),
.I3(CLBLM_R_X7Y121_SLICE_X8Y121_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y124_SLICE_X8Y124_BO5),
.O6(CLBLM_R_X7Y124_SLICE_X8Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa33aa00aa30aa00)
  ) CLBLM_R_X7Y124_SLICE_X8Y124_ALUT (
.I0(CLBLM_R_X3Y124_SLICE_X2Y124_B5Q),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I5(CLBLM_R_X7Y116_SLICE_X8Y116_AQ),
.O5(CLBLM_R_X7Y124_SLICE_X8Y124_AO5),
.O6(CLBLM_R_X7Y124_SLICE_X8Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y124_SLICE_X9Y124_AO6),
.Q(CLBLM_R_X7Y124_SLICE_X9Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffeeffee)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_DLUT (
.I0(CLBLM_R_X11Y124_SLICE_X14Y124_AQ),
.I1(CLBLM_L_X8Y121_SLICE_X11Y121_CQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y129_SLICE_X9Y129_DQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y120_SLICE_X2Y120_BQ),
.O5(CLBLM_R_X7Y124_SLICE_X9Y124_DO5),
.O6(CLBLM_R_X7Y124_SLICE_X9Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000fffffffe)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_CLUT (
.I0(CLBLM_R_X7Y121_SLICE_X9Y121_CO6),
.I1(CLBLM_R_X7Y124_SLICE_X9Y124_AQ),
.I2(CLBLM_R_X7Y123_SLICE_X9Y123_AQ),
.I3(CLBLM_R_X7Y127_SLICE_X8Y127_CQ),
.I4(CLBLM_R_X7Y124_SLICE_X9Y124_DO6),
.I5(CLBLM_R_X11Y125_SLICE_X14Y125_CQ),
.O5(CLBLM_R_X7Y124_SLICE_X9Y124_CO5),
.O6(CLBLM_R_X7Y124_SLICE_X9Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc0c0c00770077)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_BLUT (
.I0(CLBLM_R_X3Y123_SLICE_X3Y123_AQ),
.I1(CLBLM_R_X3Y128_SLICE_X2Y128_AO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.I4(CLBLM_L_X10Y123_SLICE_X13Y123_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y124_SLICE_X9Y124_BO5),
.O6(CLBLM_R_X7Y124_SLICE_X9Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0f00aaaa0f00)
  ) CLBLM_R_X7Y124_SLICE_X9Y124_ALUT (
.I0(CLBLM_R_X7Y120_SLICE_X8Y120_DQ),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y124_SLICE_X9Y124_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y124_SLICE_X9Y124_AO5),
.O6(CLBLM_R_X7Y124_SLICE_X9Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X8Y125_AO6),
.Q(CLBLM_R_X7Y125_SLICE_X8Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X8Y125_BO6),
.Q(CLBLM_R_X7Y125_SLICE_X8Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X8Y125_CO6),
.Q(CLBLM_R_X7Y125_SLICE_X8Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X8Y125_DO6),
.Q(CLBLM_R_X7Y125_SLICE_X8Y125_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfa00ccccfafa)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_DLUT (
.I0(CLBLM_R_X7Y122_SLICE_X8Y122_AQ),
.I1(CLBLM_R_X7Y127_SLICE_X8Y127_CQ),
.I2(CLBLM_R_X7Y125_SLICE_X8Y125_DQ),
.I3(CLBLM_R_X11Y120_SLICE_X14Y120_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y123_SLICE_X9Y123_A5Q),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_DO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc05050a0a)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_CLUT (
.I0(CLBLM_R_X7Y123_SLICE_X8Y123_CO5),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_AQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(1'b1),
.I4(CLBLM_L_X8Y127_SLICE_X11Y127_DQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_CO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00033f0f03300)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y126_SLICE_X8Y126_AQ),
.I3(CLBLL_L_X4Y122_SLICE_X4Y122_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y124_SLICE_X8Y124_DO6),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_BO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccaaccaaccaa)
  ) CLBLM_R_X7Y125_SLICE_X8Y125_ALUT (
.I0(CLBLL_L_X4Y120_SLICE_X5Y120_AQ),
.I1(CLBLM_R_X11Y125_SLICE_X14Y125_CQ),
.I2(CLBLM_R_X7Y125_SLICE_X8Y125_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.I5(CLBLL_L_X4Y125_SLICE_X4Y125_BQ),
.O5(CLBLM_R_X7Y125_SLICE_X8Y125_AO5),
.O6(CLBLM_R_X7Y125_SLICE_X8Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y125_SLICE_X10Y125_BO6),
.Q(CLBLM_R_X7Y125_SLICE_X9Y125_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X9Y127_DO6),
.Q(CLBLM_R_X7Y125_SLICE_X9Y125_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X9Y125_AO6),
.Q(CLBLM_R_X7Y125_SLICE_X9Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X9Y125_BO6),
.Q(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X9Y125_CO6),
.Q(CLBLM_R_X7Y125_SLICE_X9Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y125_SLICE_X9Y125_DO6),
.Q(CLBLM_R_X7Y125_SLICE_X9Y125_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa3333aaaa3030)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_DLUT (
.I0(CLBLM_L_X8Y123_SLICE_X10Y123_CQ),
.I1(CLBLM_L_X10Y129_SLICE_X13Y129_DO6),
.I2(CLBLM_R_X7Y125_SLICE_X9Y125_DQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y127_SLICE_X12Y127_CQ),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_DO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00fcaaaa00fc)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_CLUT (
.I0(CLBLM_R_X7Y123_SLICE_X8Y123_AQ),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_CQ),
.I2(CLBLM_L_X10Y125_SLICE_X12Y125_CQ),
.I3(CLBLM_L_X10Y129_SLICE_X13Y129_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_CO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000e0eff00eeee)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_BLUT (
.I0(CLBLM_R_X3Y123_SLICE_X3Y123_AQ),
.I1(CLBLM_R_X7Y125_SLICE_X9Y125_BQ),
.I2(CLBLM_L_X8Y121_SLICE_X11Y121_BQ),
.I3(CLBLM_L_X10Y126_SLICE_X12Y126_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y125_SLICE_X4Y125_BQ),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_BO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffaeaffff5040)
  ) CLBLM_R_X7Y125_SLICE_X9Y125_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X7Y125_SLICE_X9Y125_AQ),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I4(CLBLM_R_X7Y120_SLICE_X9Y120_BO6),
.I5(CLBLM_R_X5Y126_SLICE_X7Y126_AQ),
.O5(CLBLM_R_X7Y125_SLICE_X9Y125_AO5),
.O6(CLBLM_R_X7Y125_SLICE_X9Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X8Y126_AO6),
.Q(CLBLM_R_X7Y126_SLICE_X8Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X8Y126_BO6),
.Q(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X8Y126_CO6),
.Q(CLBLM_R_X7Y126_SLICE_X8Y126_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffbffffffffff)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y128_SLICE_X11Y128_DQ),
.I2(CLBLM_R_X7Y120_SLICE_X8Y120_DQ),
.I3(CLBLM_L_X8Y127_SLICE_X11Y127_CQ),
.I4(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.I5(CLBLM_L_X8Y126_SLICE_X10Y126_AO5),
.O5(CLBLM_R_X7Y126_SLICE_X8Y126_DO5),
.O6(CLBLM_R_X7Y126_SLICE_X8Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0f0aaaacccc)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_CLUT (
.I0(CLBLM_L_X8Y123_SLICE_X11Y123_AQ),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_CQ),
.I2(CLBLM_R_X11Y126_SLICE_X14Y126_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y126_SLICE_X7Y126_CO5),
.O5(CLBLM_R_X7Y126_SLICE_X8Y126_CO5),
.O6(CLBLM_R_X7Y126_SLICE_X8Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaf0f0cccc)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_BLUT (
.I0(CLBLM_R_X7Y124_SLICE_X8Y124_B5Q),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.I2(CLBLM_L_X8Y123_SLICE_X11Y123_AQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y126_SLICE_X7Y126_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y126_SLICE_X8Y126_BO5),
.O6(CLBLM_R_X7Y126_SLICE_X8Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf5cca0ccf5cca0)
  ) CLBLM_R_X7Y126_SLICE_X8Y126_ALUT (
.I0(CLBLM_L_X10Y129_SLICE_X13Y129_DO6),
.I1(CLBLM_L_X8Y126_SLICE_X11Y126_DQ),
.I2(CLBLM_R_X7Y126_SLICE_X8Y126_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X8Y126_AO5),
.O6(CLBLM_R_X7Y126_SLICE_X8Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X9Y126_BO5),
.Q(CLBLM_R_X7Y126_SLICE_X9Y126_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X9Y126_CO5),
.Q(CLBLM_R_X7Y126_SLICE_X9Y126_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X9Y126_DO5),
.Q(CLBLM_R_X7Y126_SLICE_X9Y126_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X9Y126_AO6),
.Q(CLBLM_R_X7Y126_SLICE_X9Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X9Y126_BO6),
.Q(CLBLM_R_X7Y126_SLICE_X9Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X9Y126_CO6),
.Q(CLBLM_R_X7Y126_SLICE_X9Y126_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y126_SLICE_X9Y126_DO6),
.Q(CLBLM_R_X7Y126_SLICE_X9Y126_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf505f000fcfc0c0c)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLL_L_X4Y122_SLICE_X4Y122_A5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y121_SLICE_X10Y121_BQ),
.I4(CLBLM_L_X10Y127_SLICE_X12Y127_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X9Y126_DO5),
.O6(CLBLM_R_X7Y126_SLICE_X9Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf4f40404cfc0cfc0)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y126_SLICE_X9Y126_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y128_SLICE_X4Y128_AO6),
.I4(CLBLM_L_X10Y125_SLICE_X12Y125_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X9Y126_CO5),
.O6(CLBLM_R_X7Y126_SLICE_X9Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee4444fa50fa50)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y129_SLICE_X12Y129_BQ),
.I2(CLBLM_R_X7Y130_SLICE_X9Y130_AQ),
.I3(CLBLM_L_X10Y124_SLICE_X13Y124_DQ),
.I4(CLBLM_R_X7Y116_SLICE_X9Y116_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y126_SLICE_X9Y126_BO5),
.O6(CLBLM_R_X7Y126_SLICE_X9Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h888888dd88dd8888)
  ) CLBLM_R_X7Y126_SLICE_X9Y126_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y129_SLICE_X9Y129_BQ),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X7Y125_SLICE_X8Y125_CQ),
.I5(CLBLM_R_X7Y127_SLICE_X9Y127_DO5),
.O5(CLBLM_R_X7Y126_SLICE_X9Y126_AO5),
.O6(CLBLM_R_X7Y126_SLICE_X9Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X8Y127_AO6),
.Q(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X8Y127_BO6),
.Q(CLBLM_R_X7Y127_SLICE_X8Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X8Y127_CO6),
.Q(CLBLM_R_X7Y127_SLICE_X8Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X8Y127_DO6),
.Q(CLBLM_R_X7Y127_SLICE_X8Y127_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aafcaafc)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_DLUT (
.I0(CLBLM_R_X7Y130_SLICE_X9Y130_AQ),
.I1(CLBLM_R_X3Y124_SLICE_X2Y124_B5Q),
.I2(CLBLM_R_X7Y127_SLICE_X8Y127_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLL_L_X2Y119_SLICE_X1Y119_BO6),
.O5(CLBLM_R_X7Y127_SLICE_X8Y127_DO5),
.O6(CLBLM_R_X7Y127_SLICE_X8Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0044444444)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y127_SLICE_X8Y127_CQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y128_SLICE_X8Y128_CQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y127_SLICE_X8Y127_CO5),
.O6(CLBLM_R_X7Y127_SLICE_X8Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff0ccf000f0cc)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y127_SLICE_X8Y127_BQ),
.I2(CLBLM_R_X7Y125_SLICE_X8Y125_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y126_SLICE_X7Y126_CO5),
.I5(CLBLM_L_X8Y121_SLICE_X10Y121_BQ),
.O5(CLBLM_R_X7Y127_SLICE_X8Y127_BO5),
.O6(CLBLM_R_X7Y127_SLICE_X8Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc55cc50cc55cc50)
  ) CLBLM_R_X7Y127_SLICE_X8Y127_ALUT (
.I0(CLBLM_L_X10Y129_SLICE_X13Y129_DO6),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.I2(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y119_SLICE_X9Y119_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y127_SLICE_X8Y127_AO5),
.O6(CLBLM_R_X7Y127_SLICE_X8Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X9Y127_AO6),
.Q(CLBLM_R_X7Y127_SLICE_X9Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X9Y127_BO6),
.Q(CLBLM_R_X7Y127_SLICE_X9Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y127_SLICE_X9Y127_CO6),
.Q(CLBLM_R_X7Y127_SLICE_X9Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5e4a0a0ffcc0000)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y122_SLICE_X11Y122_AQ),
.I2(CLBLM_R_X7Y126_SLICE_X9Y126_B5Q),
.I3(CLBLM_R_X7Y127_SLICE_X9Y127_AQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y127_SLICE_X9Y127_DO5),
.O6(CLBLM_R_X7Y127_SLICE_X9Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haeff0455aeaa0400)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y127_SLICE_X9Y127_CQ),
.I2(CLBLM_R_X7Y130_SLICE_X8Y130_CO6),
.I3(CLBLM_R_X5Y130_SLICE_X7Y130_DO6),
.I4(CLBLM_R_X7Y127_SLICE_X8Y127_DQ),
.I5(CLBLM_L_X8Y128_SLICE_X11Y128_BQ),
.O5(CLBLM_R_X7Y127_SLICE_X9Y127_CO5),
.O6(CLBLM_R_X7Y127_SLICE_X9Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffd0f0f0f0d)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_BLUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y129_SLICE_X12Y129_CO6),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_R_X5Y118_SLICE_X6Y118_B5Q),
.O5(CLBLM_R_X7Y127_SLICE_X9Y127_BO5),
.O6(CLBLM_R_X7Y127_SLICE_X9Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefedcdcfeeedccc)
  ) CLBLM_R_X7Y127_SLICE_X9Y127_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y120_SLICE_X9Y120_AO6),
.I2(CLBLM_R_X7Y127_SLICE_X9Y127_AQ),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I4(CLBLM_R_X7Y127_SLICE_X8Y127_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X7Y127_SLICE_X9Y127_AO5),
.O6(CLBLM_R_X7Y127_SLICE_X9Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X8Y128_AO6),
.Q(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X8Y128_BO6),
.Q(CLBLM_R_X7Y128_SLICE_X8Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X8Y128_CO6),
.Q(CLBLM_R_X7Y128_SLICE_X8Y128_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X8Y128_DO6),
.Q(CLBLM_R_X7Y128_SLICE_X8Y128_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfeccfe00320032)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_DLUT (
.I0(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y128_SLICE_X8Y128_DQ),
.I3(CLBLM_R_X5Y126_SLICE_X7Y126_CO5),
.I4(1'b1),
.I5(CLBLM_L_X8Y126_SLICE_X10Y126_AQ),
.O5(CLBLM_R_X7Y128_SLICE_X8Y128_DO5),
.O6(CLBLM_R_X7Y128_SLICE_X8Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaee5044faee5044)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y128_SLICE_X8Y128_CQ),
.I2(CLBLM_R_X7Y125_SLICE_X8Y125_BQ),
.I3(CLBLM_R_X5Y126_SLICE_X7Y126_CO5),
.I4(CLBLM_L_X8Y129_SLICE_X11Y129_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y128_SLICE_X8Y128_CO5),
.O6(CLBLM_R_X7Y128_SLICE_X8Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ccccf0f0aaaa)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_BLUT (
.I0(CLBLM_L_X8Y128_SLICE_X11Y128_DQ),
.I1(CLBLM_R_X7Y128_SLICE_X8Y128_BQ),
.I2(CLBLM_R_X5Y125_SLICE_X6Y125_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y126_SLICE_X7Y126_CO5),
.O5(CLBLM_R_X7Y128_SLICE_X8Y128_BO5),
.O6(CLBLM_R_X7Y128_SLICE_X8Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffc00fcff300030)
  ) CLBLM_R_X7Y128_SLICE_X8Y128_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y126_SLICE_X7Y126_CO5),
.I2(CLBLM_R_X7Y128_SLICE_X8Y128_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y126_SLICE_X13Y126_CQ),
.I5(CLBLM_L_X8Y127_SLICE_X11Y127_CQ),
.O5(CLBLM_R_X7Y128_SLICE_X8Y128_AO5),
.O6(CLBLM_R_X7Y128_SLICE_X8Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y128_SLICE_X9Y128_AO6),
.Q(CLBLM_R_X7Y128_SLICE_X9Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333f3f37373f3f)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_DLUT (
.I0(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.I1(CLBLM_R_X5Y130_SLICE_X7Y130_CO5),
.I2(CLBLM_R_X7Y131_SLICE_X9Y131_DO6),
.I3(1'b1),
.I4(CLBLM_R_X5Y120_SLICE_X7Y120_AQ),
.I5(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.O5(CLBLM_R_X7Y128_SLICE_X9Y128_DO5),
.O6(CLBLM_R_X7Y128_SLICE_X9Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbb050f4444faf0)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_CLUT (
.I0(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I1(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.I2(CLBLM_L_X8Y129_SLICE_X11Y129_B5Q),
.I3(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.I4(CLBLM_R_X5Y120_SLICE_X7Y120_AQ),
.I5(CLBLM_R_X5Y118_SLICE_X7Y118_BO6),
.O5(CLBLM_R_X7Y128_SLICE_X9Y128_CO5),
.O6(CLBLM_R_X7Y128_SLICE_X9Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000ccfcfcfcf)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(RIOB33_X105Y135_IOB_X1Y135_I),
.I4(CLBLM_L_X10Y129_SLICE_X12Y129_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y128_SLICE_X9Y128_BO5),
.O6(CLBLM_R_X7Y128_SLICE_X9Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff002222ff00e2e2)
  ) CLBLM_R_X7Y128_SLICE_X9Y128_ALUT (
.I0(CLBLM_L_X8Y127_SLICE_X11Y127_AQ),
.I1(CLBLM_R_X5Y130_SLICE_X7Y130_DO6),
.I2(CLBLM_R_X7Y128_SLICE_X9Y128_AQ),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_D5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y130_SLICE_X8Y130_CO6),
.O5(CLBLM_R_X7Y128_SLICE_X9Y128_AO5),
.O6(CLBLM_R_X7Y128_SLICE_X9Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X8Y129_AO5),
.Q(CLBLM_R_X7Y129_SLICE_X8Y129_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X8Y129_AO6),
.Q(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X8Y129_BO6),
.Q(CLBLM_R_X7Y129_SLICE_X8Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X8Y129_CO6),
.Q(CLBLM_R_X7Y129_SLICE_X8Y129_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X8Y129_DO6),
.Q(CLBLM_R_X7Y129_SLICE_X8Y129_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe54fe54ba10ba10)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y129_SLICE_X13Y129_DO6),
.I2(CLBLM_R_X7Y129_SLICE_X8Y129_DQ),
.I3(CLBLM_R_X5Y128_SLICE_X6Y128_AQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y127_SLICE_X11Y127_DQ),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_DO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafc0caaaafc0c)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_CLUT (
.I0(CLBLM_R_X7Y129_SLICE_X8Y129_BQ),
.I1(CLBLM_R_X7Y129_SLICE_X8Y129_CQ),
.I2(CLBLM_L_X10Y129_SLICE_X13Y129_DO6),
.I3(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_CO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcfcfcfcfc0c0)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y126_SLICE_X9Y126_C5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X7Y131_SLICE_X9Y131_BO5),
.I5(CLBLM_R_X7Y129_SLICE_X9Y129_CQ),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_BO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heaeaeaeafff00f00)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_ALUT (
.I0(CLBLM_R_X7Y130_SLICE_X8Y130_DO6),
.I1(CLBLM_L_X8Y122_SLICE_X10Y122_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y126_SLICE_X4Y126_DO6),
.I4(CLBLM_R_X7Y117_SLICE_X8Y117_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_AO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X9Y129_AO6),
.Q(CLBLM_R_X7Y129_SLICE_X9Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X9Y129_BO6),
.Q(CLBLM_R_X7Y129_SLICE_X9Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X9Y129_CO6),
.Q(CLBLM_R_X7Y129_SLICE_X9Y129_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y129_SLICE_X9Y129_DO6),
.Q(CLBLM_R_X7Y129_SLICE_X9Y129_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888d8d88888d8d8)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y129_SLICE_X9Y129_CQ),
.I2(CLBLM_R_X7Y129_SLICE_X9Y129_DQ),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_DO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc55005500)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_CLUT (
.I0(CLBLM_R_X7Y131_SLICE_X9Y131_BO5),
.I1(CLBLM_R_X3Y126_SLICE_X2Y126_AQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y129_SLICE_X9Y129_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_CO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fcfc00000c0c)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y129_SLICE_X6Y129_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X7Y131_SLICE_X9Y131_BO5),
.I5(CLBLM_R_X11Y126_SLICE_X14Y126_DQ),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_BO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0ff40550cff0455)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y131_SLICE_X9Y131_BO6),
.I2(CLBLM_R_X7Y129_SLICE_X9Y129_AQ),
.I3(CLBLM_R_X7Y131_SLICE_X8Y131_CO6),
.I4(CLBLM_R_X7Y129_SLICE_X9Y129_DQ),
.I5(CLBLM_L_X8Y129_SLICE_X10Y129_BO6),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_AO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X8Y130_AO6),
.Q(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X8Y130_BO6),
.Q(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000031313322)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_DLUT (
.I0(CLBLM_L_X8Y127_SLICE_X10Y127_AQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_R_X5Y130_SLICE_X7Y130_DO6),
.I3(CLBLM_R_X7Y130_SLICE_X8Y130_CO5),
.I4(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y130_SLICE_X8Y130_DO5),
.O6(CLBLM_R_X7Y130_SLICE_X8Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010100000200)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_CLUT (
.I0(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I1(CLBLM_L_X8Y129_SLICE_X11Y129_B5Q),
.I2(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.I3(CLBLM_R_X5Y130_SLICE_X7Y130_CO5),
.I4(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y130_SLICE_X8Y130_CO5),
.O6(CLBLM_R_X7Y130_SLICE_X8Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fff0ff505f404)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_BLUT (
.I0(CLBLM_R_X5Y130_SLICE_X7Y130_DO6),
.I1(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.I4(CLBLM_L_X8Y127_SLICE_X10Y127_AQ),
.I5(CLBLM_R_X7Y130_SLICE_X8Y130_CO6),
.O5(CLBLM_R_X7Y130_SLICE_X8Y130_BO5),
.O6(CLBLM_R_X7Y130_SLICE_X8Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff004444ff00e4e4)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_ALUT (
.I0(CLBLM_R_X5Y130_SLICE_X7Y130_DO6),
.I1(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.I2(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.I3(CLBLL_L_X4Y124_SLICE_X4Y124_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y130_SLICE_X8Y130_CO6),
.O5(CLBLM_R_X7Y130_SLICE_X8Y130_AO5),
.O6(CLBLM_R_X7Y130_SLICE_X8Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X9Y130_AO6),
.Q(CLBLM_R_X7Y130_SLICE_X9Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff23ff00ff00ff)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_DLUT (
.I0(CLBLM_R_X7Y130_SLICE_X9Y130_CO5),
.I1(CLBLM_R_X7Y128_SLICE_X9Y128_CO6),
.I2(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_AQ),
.I4(CLBLM_R_X7Y131_SLICE_X9Y131_BO5),
.I5(CLBLM_R_X5Y129_SLICE_X6Y129_BQ),
.O5(CLBLM_R_X7Y130_SLICE_X9Y130_DO5),
.O6(CLBLM_R_X7Y130_SLICE_X9Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33337777ffffffcc)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_CLUT (
.I0(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I1(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y129_SLICE_X11Y129_B5Q),
.I4(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y130_SLICE_X9Y130_CO5),
.O6(CLBLM_R_X7Y130_SLICE_X9Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7878ffff02020202)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_BLUT (
.I0(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.I1(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.I2(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y131_SLICE_X10Y131_DO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y130_SLICE_X9Y130_BO5),
.O6(CLBLM_R_X7Y130_SLICE_X9Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccf0f0aaff)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_ALUT (
.I0(CLBLM_R_X7Y130_SLICE_X9Y130_BO5),
.I1(CLBLM_L_X10Y128_SLICE_X12Y128_AQ),
.I2(CLBLM_R_X7Y124_SLICE_X9Y124_BO5),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_DO6),
.I4(CLBLM_R_X7Y130_SLICE_X8Y130_CO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y130_SLICE_X9Y130_AO5),
.O6(CLBLM_R_X7Y130_SLICE_X9Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X8Y131_AO6),
.Q(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_DO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555050555550505)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_L_X8Y131_SLICE_X10Y131_DO6),
.I3(1'b1),
.I4(CLBLM_R_X7Y131_SLICE_X8Y131_BO5),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_CO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd3d303d34647f647)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_BLUT (
.I0(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.I1(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.I2(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I3(CLBLM_L_X8Y129_SLICE_X11Y129_B5Q),
.I4(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_BO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdccd1001dcdc1010)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_ALUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I3(CLBLM_R_X7Y131_SLICE_X8Y131_BO6),
.I4(CLBLM_L_X8Y127_SLICE_X10Y127_BQ),
.I5(CLBLM_L_X8Y131_SLICE_X10Y131_DO6),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_AO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X9Y131_AO6),
.Q(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0088008800880088)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_DLUT (
.I0(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I1(CLBLM_L_X8Y129_SLICE_X11Y129_B5Q),
.I2(1'b1),
.I3(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_DO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffffff00fffdff)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_CLUT (
.I0(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I1(CLBLM_L_X8Y129_SLICE_X11Y129_B5Q),
.I2(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.I3(CLBLM_R_X5Y130_SLICE_X7Y130_CO5),
.I4(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.I5(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_CO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h555555540000cccf)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_BLUT (
.I0(CLBLM_L_X8Y131_SLICE_X10Y131_DO6),
.I1(CLBLM_L_X8Y129_SLICE_X11Y129_B5Q),
.I2(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.I3(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.I4(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_BO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc444f5554c445f55)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_ALUT (
.I0(CLBLM_R_X7Y131_SLICE_X8Y131_CO6),
.I1(CLBLM_R_X5Y127_SLICE_X7Y127_BQ),
.I2(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I3(CLBLM_R_X7Y131_SLICE_X9Y131_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y131_SLICE_X11Y131_BO6),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_AO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y119_SLICE_X14Y119_AO6),
.Q(CLBLM_R_X11Y119_SLICE_X14Y119_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y119_SLICE_X14Y119_BO6),
.Q(CLBLM_R_X11Y119_SLICE_X14Y119_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X14Y119_DO5),
.O6(CLBLM_R_X11Y119_SLICE_X14Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X14Y119_CO5),
.O6(CLBLM_R_X11Y119_SLICE_X14Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f0f0ee00)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_BLUT (
.I0(CLBLM_R_X7Y117_SLICE_X8Y117_DQ),
.I1(CLBLM_R_X11Y119_SLICE_X14Y119_BQ),
.I2(CLBLM_R_X11Y119_SLICE_X14Y119_AQ),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X11Y119_SLICE_X14Y119_BO5),
.O6(CLBLM_R_X11Y119_SLICE_X14Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000c0aac0aa)
  ) CLBLM_R_X11Y119_SLICE_X14Y119_ALUT (
.I0(CLBLM_R_X11Y123_SLICE_X14Y123_CQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X11Y119_SLICE_X14Y119_AQ),
.I3(CLBLM_L_X8Y123_SLICE_X10Y123_DO6),
.I4(CLBLM_L_X10Y122_SLICE_X12Y122_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y119_SLICE_X14Y119_AO5),
.O6(CLBLM_R_X11Y119_SLICE_X14Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X15Y119_DO5),
.O6(CLBLM_R_X11Y119_SLICE_X15Y119_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X15Y119_CO5),
.O6(CLBLM_R_X11Y119_SLICE_X15Y119_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y119_SLICE_X15Y119_BO5),
.O6(CLBLM_R_X11Y119_SLICE_X15Y119_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffeeeeeeee)
  ) CLBLM_R_X11Y119_SLICE_X15Y119_ALUT (
.I0(CLBLM_L_X10Y124_SLICE_X13Y124_BQ),
.I1(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y120_SLICE_X12Y120_CQ),
.O5(CLBLM_R_X11Y119_SLICE_X15Y119_AO5),
.O6(CLBLM_R_X11Y119_SLICE_X15Y119_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y120_SLICE_X14Y120_AO6),
.Q(CLBLM_R_X11Y120_SLICE_X14Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y120_SLICE_X14Y120_BO6),
.Q(CLBLM_R_X11Y120_SLICE_X14Y120_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y120_SLICE_X14Y120_CO6),
.Q(CLBLM_R_X11Y120_SLICE_X14Y120_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f7f3f3f7f)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_DLUT (
.I0(CLBLM_L_X10Y121_SLICE_X13Y121_DO6),
.I1(CLBLM_L_X8Y123_SLICE_X10Y123_DO6),
.I2(CLBLM_R_X11Y120_SLICE_X15Y120_BO5),
.I3(CLBLM_R_X11Y120_SLICE_X15Y120_DO6),
.I4(CLBLM_R_X7Y120_SLICE_X9Y120_DO6),
.I5(CLBLM_L_X8Y120_SLICE_X11Y120_AO6),
.O5(CLBLM_R_X11Y120_SLICE_X14Y120_DO5),
.O6(CLBLM_R_X11Y120_SLICE_X14Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000feaa5400)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y120_SLICE_X14Y120_CQ),
.I2(CLBLM_R_X5Y120_SLICE_X7Y120_DO6),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I4(CLBLM_L_X10Y122_SLICE_X13Y122_CQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X11Y120_SLICE_X14Y120_CO5),
.O6(CLBLM_R_X11Y120_SLICE_X14Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8f8fff008080f00)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X11Y120_SLICE_X14Y120_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y121_SLICE_X14Y121_AQ),
.I4(CLBLM_L_X8Y123_SLICE_X10Y123_DO6),
.I5(CLBLM_R_X11Y123_SLICE_X14Y123_AQ),
.O5(CLBLM_R_X11Y120_SLICE_X14Y120_BO5),
.O6(CLBLM_R_X11Y120_SLICE_X14Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff002800000028)
  ) CLBLM_R_X11Y120_SLICE_X14Y120_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X11Y120_SLICE_X15Y120_CO5),
.I2(CLBLM_R_X11Y120_SLICE_X14Y120_AQ),
.I3(CLBLM_R_X5Y127_SLICE_X7Y127_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y124_SLICE_X10Y124_AQ),
.O5(CLBLM_R_X11Y120_SLICE_X14Y120_AO5),
.O6(CLBLM_R_X11Y120_SLICE_X14Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y120_SLICE_X15Y120_AO6),
.Q(CLBLM_R_X11Y120_SLICE_X15Y120_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3c3c3c3c3c3c1c1)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_DLUT (
.I0(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I1(CLBLM_R_X11Y119_SLICE_X14Y119_AQ),
.I2(CLBLM_R_X11Y123_SLICE_X14Y123_CQ),
.I3(1'b1),
.I4(CLBLM_R_X11Y121_SLICE_X15Y121_DO6),
.I5(CLBLM_R_X11Y119_SLICE_X15Y119_AO6),
.O5(CLBLM_R_X11Y120_SLICE_X15Y120_DO5),
.O6(CLBLM_R_X11Y120_SLICE_X15Y120_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00080808040c0c0c)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_CLUT (
.I0(CLBLM_R_X11Y120_SLICE_X14Y120_AQ),
.I1(CLBLM_R_X11Y123_SLICE_X15Y123_AQ),
.I2(CLBLM_L_X8Y123_SLICE_X10Y123_DO6),
.I3(CLBLM_R_X11Y120_SLICE_X15Y120_AQ),
.I4(CLBLM_R_X11Y121_SLICE_X15Y121_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y120_SLICE_X15Y120_CO5),
.O6(CLBLM_R_X11Y120_SLICE_X15Y120_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h02000000a0000000)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_BLUT (
.I0(CLBLM_R_X11Y121_SLICE_X15Y121_AQ),
.I1(CLBLM_L_X8Y123_SLICE_X10Y123_DO6),
.I2(CLBLM_R_X11Y120_SLICE_X15Y120_AQ),
.I3(CLBLM_R_X11Y123_SLICE_X15Y123_AQ),
.I4(CLBLM_R_X11Y120_SLICE_X14Y120_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y120_SLICE_X15Y120_BO5),
.O6(CLBLM_R_X11Y120_SLICE_X15Y120_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f2f0f003020000)
  ) CLBLM_R_X11Y120_SLICE_X15Y120_ALUT (
.I0(CLBLM_R_X11Y120_SLICE_X15Y120_AQ),
.I1(CLBLM_R_X5Y127_SLICE_X7Y127_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y120_SLICE_X15Y120_BO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X11Y122_SLICE_X14Y122_CQ),
.O5(CLBLM_R_X11Y120_SLICE_X15Y120_AO5),
.O6(CLBLM_R_X11Y120_SLICE_X15Y120_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y121_SLICE_X14Y121_AO6),
.Q(CLBLM_R_X11Y121_SLICE_X14Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y121_SLICE_X14Y121_BO6),
.Q(CLBLM_R_X11Y121_SLICE_X14Y121_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y121_SLICE_X14Y121_CO6),
.Q(CLBLM_R_X11Y121_SLICE_X14Y121_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_DLUT (
.I0(CLBLM_R_X11Y121_SLICE_X14Y121_BQ),
.I1(CLBLM_R_X11Y121_SLICE_X14Y121_CQ),
.I2(CLBLM_L_X12Y121_SLICE_X16Y121_AQ),
.I3(CLBLM_R_X11Y120_SLICE_X14Y120_BQ),
.I4(CLBLM_R_X11Y123_SLICE_X14Y123_BQ),
.I5(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.O5(CLBLM_R_X11Y121_SLICE_X14Y121_DO5),
.O6(CLBLM_R_X11Y121_SLICE_X14Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44aa00fa50fa50)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y121_SLICE_X14Y121_CQ),
.I2(CLBLM_L_X12Y121_SLICE_X16Y121_AQ),
.I3(CLBLM_L_X8Y121_SLICE_X10Y121_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X8Y123_SLICE_X10Y123_DO6),
.O5(CLBLM_R_X11Y121_SLICE_X14Y121_CO5),
.O6(CLBLM_R_X11Y121_SLICE_X14Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4a0a0f5a0f5a0)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y121_SLICE_X8Y121_AQ),
.I3(CLBLM_R_X11Y123_SLICE_X14Y123_BQ),
.I4(CLBLM_R_X11Y121_SLICE_X14Y121_BQ),
.I5(CLBLM_L_X8Y123_SLICE_X10Y123_DO6),
.O5(CLBLM_R_X11Y121_SLICE_X14Y121_BO5),
.O6(CLBLM_R_X11Y121_SLICE_X14Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf000aaaacccc)
  ) CLBLM_R_X11Y121_SLICE_X14Y121_ALUT (
.I0(CLBLL_L_X4Y124_SLICE_X4Y124_DQ),
.I1(CLBLM_L_X8Y121_SLICE_X11Y121_AQ),
.I2(CLBLM_R_X11Y121_SLICE_X14Y121_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y123_SLICE_X10Y123_DO6),
.O5(CLBLM_R_X11Y121_SLICE_X14Y121_AO5),
.O6(CLBLM_R_X11Y121_SLICE_X14Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y121_SLICE_X15Y121_AO6),
.Q(CLBLM_R_X11Y121_SLICE_X15Y121_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffeeffee)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_DLUT (
.I0(CLBLM_R_X11Y121_SLICE_X14Y121_AQ),
.I1(CLBLM_L_X10Y121_SLICE_X12Y121_BQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y122_SLICE_X15Y122_AQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y122_SLICE_X15Y122_BQ),
.O5(CLBLM_R_X11Y121_SLICE_X15Y121_DO5),
.O6(CLBLM_R_X11Y121_SLICE_X15Y121_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30fcfcfc303030)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y120_SLICE_X15Y120_BO5),
.I2(CLBLM_R_X7Y120_SLICE_X9Y120_DO6),
.I3(CLBLM_R_X11Y123_SLICE_X14Y123_CQ),
.I4(CLBLM_R_X11Y119_SLICE_X14Y119_AQ),
.I5(CLBLM_R_X11Y121_SLICE_X15Y121_BO6),
.O5(CLBLM_R_X11Y121_SLICE_X15Y121_CO5),
.O6(CLBLM_R_X11Y121_SLICE_X15Y121_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0e0f)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_BLUT (
.I0(CLBLM_R_X11Y121_SLICE_X15Y121_DO6),
.I1(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.I2(CLBLM_R_X11Y123_SLICE_X14Y123_CQ),
.I3(CLBLM_R_X11Y121_SLICE_X14Y121_DO6),
.I4(CLBLM_L_X10Y120_SLICE_X12Y120_CQ),
.I5(CLBLM_L_X10Y124_SLICE_X13Y124_BQ),
.O5(CLBLM_R_X11Y121_SLICE_X15Y121_BO5),
.O6(CLBLM_R_X11Y121_SLICE_X15Y121_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000480048)
  ) CLBLM_R_X11Y121_SLICE_X15Y121_ALUT (
.I0(CLBLM_R_X11Y120_SLICE_X15Y120_CO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X11Y121_SLICE_X15Y121_AQ),
.I3(CLBLM_R_X5Y127_SLICE_X7Y127_BQ),
.I4(CLBLM_R_X11Y126_SLICE_X14Y126_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y121_SLICE_X15Y121_AO5),
.O6(CLBLM_R_X11Y121_SLICE_X15Y121_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y122_SLICE_X14Y122_AO6),
.Q(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y122_SLICE_X14Y122_BO6),
.Q(CLBLM_R_X11Y122_SLICE_X14Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y122_SLICE_X14Y122_CO6),
.Q(CLBLM_R_X11Y122_SLICE_X14Y122_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y122_SLICE_X14Y122_DO6),
.Q(CLBLM_R_X11Y122_SLICE_X14Y122_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefedcdcfeeedccc)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y122_SLICE_X11Y122_BO6),
.I2(CLBLM_R_X11Y122_SLICE_X14Y122_DQ),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I4(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X11Y122_SLICE_X14Y122_DO5),
.O6(CLBLM_R_X11Y122_SLICE_X14Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcccecc03000200)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_CLUT (
.I0(CLBLM_L_X10Y119_SLICE_X12Y119_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I4(CLBLM_R_X11Y122_SLICE_X14Y122_CQ),
.I5(CLBLM_R_X11Y124_SLICE_X14Y124_BQ),
.O5(CLBLM_R_X11Y122_SLICE_X14Y122_CO5),
.O6(CLBLM_R_X11Y122_SLICE_X14Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefefef00e0e0e00)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_BLUT (
.I0(CLBLM_R_X11Y122_SLICE_X14Y122_CQ),
.I1(CLBLM_R_X11Y122_SLICE_X14Y122_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I5(CLBLM_R_X11Y124_SLICE_X14Y124_A5Q),
.O5(CLBLM_R_X11Y122_SLICE_X14Y122_BO5),
.O6(CLBLM_R_X11Y122_SLICE_X14Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff00e0e0)
  ) CLBLM_R_X11Y122_SLICE_X14Y122_ALUT (
.I0(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.I3(CLBLM_L_X8Y122_SLICE_X11Y122_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y122_SLICE_X11Y122_BO6),
.O5(CLBLM_R_X11Y122_SLICE_X14Y122_AO5),
.O6(CLBLM_R_X11Y122_SLICE_X14Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y122_SLICE_X15Y122_AO6),
.Q(CLBLM_R_X11Y122_SLICE_X15Y122_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y122_SLICE_X15Y122_BO6),
.Q(CLBLM_R_X11Y122_SLICE_X15Y122_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y122_SLICE_X15Y122_DO5),
.O6(CLBLM_R_X11Y122_SLICE_X15Y122_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y122_SLICE_X15Y122_CO5),
.O6(CLBLM_R_X11Y122_SLICE_X15Y122_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff008f8fff008080)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X11Y122_SLICE_X15Y122_BQ),
.I2(CLBLM_L_X8Y123_SLICE_X10Y123_DO6),
.I3(CLBLM_R_X7Y126_SLICE_X9Y126_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y124_SLICE_X13Y124_BQ),
.O5(CLBLM_R_X11Y122_SLICE_X15Y122_BO5),
.O6(CLBLM_R_X11Y122_SLICE_X15Y122_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaccaa00aacc)
  ) CLBLM_R_X11Y122_SLICE_X15Y122_ALUT (
.I0(CLBLM_R_X11Y126_SLICE_X15Y126_AQ),
.I1(CLBLM_R_X11Y122_SLICE_X15Y122_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y123_SLICE_X10Y123_DO6),
.I5(CLBLM_R_X11Y122_SLICE_X15Y122_AQ),
.O5(CLBLM_R_X11Y122_SLICE_X15Y122_AO5),
.O6(CLBLM_R_X11Y122_SLICE_X15Y122_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y123_SLICE_X14Y123_AO6),
.Q(CLBLM_R_X11Y123_SLICE_X14Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y123_SLICE_X14Y123_BO6),
.Q(CLBLM_R_X11Y123_SLICE_X14Y123_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y123_SLICE_X14Y123_CO6),
.Q(CLBLM_R_X11Y123_SLICE_X14Y123_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y123_SLICE_X14Y123_DO6),
.Q(CLBLM_R_X11Y123_SLICE_X14Y123_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5c5c5c5c0c0c0c0)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X11Y123_SLICE_X14Y123_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_CQ),
.O5(CLBLM_R_X11Y123_SLICE_X14Y123_DO5),
.O6(CLBLM_R_X11Y123_SLICE_X14Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf808ff0ff808f000)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X11Y123_SLICE_X14Y123_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y125_SLICE_X11Y125_AQ),
.I4(CLBLM_L_X8Y123_SLICE_X10Y123_DO6),
.I5(CLBLM_R_X11Y121_SLICE_X14Y121_BQ),
.O5(CLBLM_R_X11Y123_SLICE_X14Y123_CO5),
.O6(CLBLM_R_X11Y123_SLICE_X14Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfaf0fa0c0a000a)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_BLUT (
.I0(CLBLM_R_X11Y120_SLICE_X14Y120_BQ),
.I1(CLBLM_R_X11Y123_SLICE_X14Y123_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y123_SLICE_X10Y123_DO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X10Y126_SLICE_X13Y126_BQ),
.O5(CLBLM_R_X11Y123_SLICE_X14Y123_BO5),
.O6(CLBLM_R_X11Y123_SLICE_X14Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaccccaaaaccf0)
  ) CLBLM_R_X11Y123_SLICE_X14Y123_ALUT (
.I0(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.I1(CLBLM_R_X11Y119_SLICE_X14Y119_BQ),
.I2(CLBLM_R_X11Y123_SLICE_X14Y123_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.O5(CLBLM_R_X11Y123_SLICE_X14Y123_AO5),
.O6(CLBLM_R_X11Y123_SLICE_X14Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y123_SLICE_X15Y123_AO6),
.Q(CLBLM_R_X11Y123_SLICE_X15Y123_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y123_SLICE_X15Y123_DO5),
.O6(CLBLM_R_X11Y123_SLICE_X15Y123_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y123_SLICE_X15Y123_CO5),
.O6(CLBLM_R_X11Y123_SLICE_X15Y123_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y123_SLICE_X15Y123_BO5),
.O6(CLBLM_R_X11Y123_SLICE_X15Y123_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa2a2a2ff828282)
  ) CLBLM_R_X11Y123_SLICE_X15Y123_ALUT (
.I0(CLBLM_R_X11Y126_SLICE_X14Y126_AO5),
.I1(CLBLM_L_X8Y123_SLICE_X10Y123_DO6),
.I2(CLBLM_R_X11Y123_SLICE_X15Y123_AQ),
.I3(CLBLM_R_X11Y127_SLICE_X14Y127_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y120_SLICE_X15Y120_BO5),
.O5(CLBLM_R_X11Y123_SLICE_X15Y123_AO5),
.O6(CLBLM_R_X11Y123_SLICE_X15Y123_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X14Y124_AO5),
.Q(CLBLM_R_X11Y124_SLICE_X14Y124_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X14Y124_AO6),
.Q(CLBLM_R_X11Y124_SLICE_X14Y124_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X14Y124_BO6),
.Q(CLBLM_R_X11Y124_SLICE_X14Y124_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y124_SLICE_X14Y124_CO6),
.Q(CLBLM_R_X11Y124_SLICE_X14Y124_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000fcfc0000ffaa)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_DLUT (
.I0(CLBLM_R_X11Y122_SLICE_X14Y122_AQ),
.I1(CLBLM_R_X7Y119_SLICE_X9Y119_BQ),
.I2(CLBLM_R_X11Y124_SLICE_X14Y124_BQ),
.I3(CLBLM_R_X11Y120_SLICE_X14Y120_CQ),
.I4(CLBLM_R_X7Y123_SLICE_X8Y123_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y124_SLICE_X14Y124_DO5),
.O6(CLBLM_R_X11Y124_SLICE_X14Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefefeaa54545400)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y124_SLICE_X14Y124_CQ),
.I2(CLBLM_R_X5Y121_SLICE_X7Y121_DO6),
.I3(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X12Y126_SLICE_X16Y126_AQ),
.O5(CLBLM_R_X11Y124_SLICE_X14Y124_CO5),
.O6(CLBLM_R_X11Y124_SLICE_X14Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffccf0f0aa88)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X11Y124_SLICE_X14Y124_BQ),
.I2(CLBLM_R_X3Y124_SLICE_X3Y124_C5Q),
.I3(CLBLM_L_X8Y124_SLICE_X11Y124_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.O5(CLBLM_R_X11Y124_SLICE_X14Y124_BO5),
.O6(CLBLM_R_X11Y124_SLICE_X14Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00c0c0f0f0aaaa)
  ) CLBLM_R_X11Y124_SLICE_X14Y124_ALUT (
.I0(CLBLM_R_X3Y123_SLICE_X3Y123_BQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X11Y124_SLICE_X14Y124_AQ),
.I3(CLBLM_L_X8Y119_SLICE_X10Y119_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y124_SLICE_X14Y124_AO5),
.O6(CLBLM_R_X11Y124_SLICE_X14Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y124_SLICE_X15Y124_DO5),
.O6(CLBLM_R_X11Y124_SLICE_X15Y124_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y124_SLICE_X15Y124_CO5),
.O6(CLBLM_R_X11Y124_SLICE_X15Y124_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y124_SLICE_X15Y124_BO5),
.O6(CLBLM_R_X11Y124_SLICE_X15Y124_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y124_SLICE_X15Y124_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y124_SLICE_X15Y124_AO5),
.O6(CLBLM_R_X11Y124_SLICE_X15Y124_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y125_SLICE_X14Y125_AO6),
.Q(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y125_SLICE_X14Y125_BO6),
.Q(CLBLM_R_X11Y125_SLICE_X14Y125_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y125_SLICE_X14Y125_CO6),
.Q(CLBLM_R_X11Y125_SLICE_X14Y125_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y125_SLICE_X14Y125_DO5),
.O6(CLBLM_R_X11Y125_SLICE_X14Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf404f404f404f404)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X11Y125_SLICE_X14Y125_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y126_SLICE_X14Y126_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y125_SLICE_X14Y125_CO5),
.O6(CLBLM_R_X11Y125_SLICE_X14Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafacacafa0aca0)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_BLUT (
.I0(CLBLM_L_X10Y124_SLICE_X13Y124_CQ),
.I1(CLBLM_R_X11Y125_SLICE_X14Y125_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X8Y124_SLICE_X10Y124_DO6),
.I5(CLBLM_R_X5Y124_SLICE_X6Y124_AQ),
.O5(CLBLM_R_X11Y125_SLICE_X14Y125_BO5),
.O6(CLBLM_R_X11Y125_SLICE_X14Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff0fa0000f0fa)
  ) CLBLM_R_X11Y125_SLICE_X14Y125_ALUT (
.I0(RIOB33_X105Y141_IOB_X1Y142_I),
.I1(1'b1),
.I2(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.I3(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y125_SLICE_X11Y125_BQ),
.O5(CLBLM_R_X11Y125_SLICE_X14Y125_AO5),
.O6(CLBLM_R_X11Y125_SLICE_X14Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y125_SLICE_X15Y125_DO5),
.O6(CLBLM_R_X11Y125_SLICE_X15Y125_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y125_SLICE_X15Y125_CO5),
.O6(CLBLM_R_X11Y125_SLICE_X15Y125_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y125_SLICE_X15Y125_BO5),
.O6(CLBLM_R_X11Y125_SLICE_X15Y125_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y125_SLICE_X15Y125_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y125_SLICE_X15Y125_AO5),
.O6(CLBLM_R_X11Y125_SLICE_X15Y125_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y126_SLICE_X14Y126_AO6),
.Q(CLBLM_R_X11Y126_SLICE_X14Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y126_SLICE_X14Y126_BO6),
.Q(CLBLM_R_X11Y126_SLICE_X14Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y126_SLICE_X14Y126_CO6),
.Q(CLBLM_R_X11Y126_SLICE_X14Y126_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y126_SLICE_X14Y126_DO6),
.Q(CLBLM_R_X11Y126_SLICE_X14Y126_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd11fd31cc00ec20)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_DLUT (
.I0(CLBLM_R_X11Y126_SLICE_X15Y126_DO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y126_SLICE_X14Y126_DQ),
.I3(CLBLM_R_X11Y123_SLICE_X14Y123_DQ),
.I4(CLBLM_L_X10Y128_SLICE_X13Y128_CO6),
.I5(CLBLM_L_X10Y128_SLICE_X12Y128_BQ),
.O5(CLBLM_R_X11Y126_SLICE_X14Y126_DO5),
.O6(CLBLM_R_X11Y126_SLICE_X14Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ffbe00be)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_CLUT (
.I0(CLBLM_R_X11Y130_SLICE_X14Y130_BO5),
.I1(CLBLM_R_X11Y126_SLICE_X14Y126_CQ),
.I2(CLBLM_R_X11Y128_SLICE_X15Y128_CO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y126_SLICE_X12Y126_CQ),
.I5(CLBLM_R_X11Y127_SLICE_X15Y127_BO5),
.O5(CLBLM_R_X11Y126_SLICE_X14Y126_CO5),
.O6(CLBLM_R_X11Y126_SLICE_X14Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000abeeabee)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_BLUT (
.I0(CLBLM_L_X10Y128_SLICE_X13Y128_CO6),
.I1(CLBLM_R_X11Y126_SLICE_X14Y126_BQ),
.I2(CLBLM_R_X11Y128_SLICE_X14Y128_AO6),
.I3(CLBLM_L_X10Y125_SLICE_X13Y125_DO5),
.I4(CLBLL_L_X2Y120_SLICE_X1Y120_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y126_SLICE_X14Y126_BO5),
.O6(CLBLM_R_X11Y126_SLICE_X14Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0c0c000000f0)
  ) CLBLM_R_X11Y126_SLICE_X14Y126_ALUT (
.I0(CLBLM_L_X10Y127_SLICE_X13Y127_DQ),
.I1(CLBLM_L_X8Y128_SLICE_X11Y128_DQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X5Y127_SLICE_X7Y127_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y126_SLICE_X14Y126_AO5),
.O6(CLBLM_R_X11Y126_SLICE_X14Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y126_SLICE_X15Y126_AO6),
.Q(CLBLM_R_X11Y126_SLICE_X15Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y126_SLICE_X15Y126_BO6),
.Q(CLBLM_R_X11Y126_SLICE_X15Y126_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y126_SLICE_X15Y126_CO6),
.Q(CLBLM_R_X11Y126_SLICE_X15Y126_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7577777700880088)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_DLUT (
.I0(CLBLM_L_X10Y125_SLICE_X13Y125_DO5),
.I1(CLBLM_L_X8Y129_SLICE_X11Y129_BQ),
.I2(CLBLM_R_X11Y127_SLICE_X15Y127_CO6),
.I3(CLBLM_R_X11Y126_SLICE_X15Y126_BQ),
.I4(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y126_SLICE_X15Y126_DO5),
.O6(CLBLM_R_X11Y126_SLICE_X15Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haeae0404ffaa5500)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y126_SLICE_X15Y126_CQ),
.I2(CLBLM_L_X10Y128_SLICE_X13Y128_CO6),
.I3(CLBLM_L_X10Y128_SLICE_X13Y128_BQ),
.I4(CLBLM_R_X5Y125_SLICE_X7Y125_BQ),
.I5(CLBLM_R_X11Y126_SLICE_X15Y126_DO5),
.O5(CLBLM_R_X11Y126_SLICE_X15Y126_CO5),
.O6(CLBLM_R_X11Y126_SLICE_X15Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000202ff000d0d)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_BLUT (
.I0(CLBLM_R_X11Y126_SLICE_X15Y126_DO6),
.I1(CLBLM_R_X11Y129_SLICE_X15Y129_AO6),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLL_L_X4Y125_SLICE_X5Y125_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y126_SLICE_X15Y126_BQ),
.O5(CLBLM_R_X11Y126_SLICE_X15Y126_BO5),
.O6(CLBLM_R_X11Y126_SLICE_X15Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f033333300)
  ) CLBLM_R_X11Y126_SLICE_X15Y126_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y127_SLICE_X15Y127_BO5),
.I2(CLBLM_R_X7Y124_SLICE_X8Y124_AQ),
.I3(CLBLM_R_X11Y128_SLICE_X15Y128_BO6),
.I4(CLBLM_R_X11Y130_SLICE_X14Y130_BO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y126_SLICE_X15Y126_AO5),
.O6(CLBLM_R_X11Y126_SLICE_X15Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y127_SLICE_X14Y127_AO6),
.Q(CLBLM_R_X11Y127_SLICE_X14Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff0f4f5f5f)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_DLUT (
.I0(CLBLM_L_X10Y128_SLICE_X12Y128_AQ),
.I1(CLBLM_L_X8Y129_SLICE_X11Y129_BQ),
.I2(CLBLM_L_X10Y127_SLICE_X13Y127_DQ),
.I3(CLBLM_R_X11Y128_SLICE_X15Y128_AQ),
.I4(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.I5(CLBLM_R_X11Y126_SLICE_X15Y126_BQ),
.O5(CLBLM_R_X11Y127_SLICE_X14Y127_DO5),
.O6(CLBLM_R_X11Y127_SLICE_X14Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fc50fcf0fca0cc)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_CLUT (
.I0(CLBLM_L_X10Y124_SLICE_X13Y124_A5Q),
.I1(CLBLM_R_X11Y127_SLICE_X14Y127_BO5),
.I2(CLBLM_R_X11Y127_SLICE_X14Y127_AQ),
.I3(CLBLM_R_X11Y130_SLICE_X14Y130_AQ),
.I4(CLBLM_R_X11Y127_SLICE_X14Y127_DO6),
.I5(CLBLM_R_X11Y127_SLICE_X14Y127_BO6),
.O5(CLBLM_R_X11Y127_SLICE_X14Y127_CO5),
.O6(CLBLM_R_X11Y127_SLICE_X14Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaf113305000500)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_BLUT (
.I0(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.I1(CLBLM_R_X11Y126_SLICE_X15Y126_BQ),
.I2(CLBLM_L_X10Y128_SLICE_X12Y128_AQ),
.I3(CLBLM_R_X11Y128_SLICE_X15Y128_AQ),
.I4(CLBLM_R_X11Y126_SLICE_X14Y126_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y127_SLICE_X14Y127_BO5),
.O6(CLBLM_R_X11Y127_SLICE_X14Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfcfcfc0c0c0)
  ) CLBLM_R_X11Y127_SLICE_X14Y127_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y127_SLICE_X15Y127_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y123_SLICE_X5Y123_CO6),
.I4(CLBLM_L_X10Y128_SLICE_X13Y128_CO6),
.I5(CLBLM_R_X11Y127_SLICE_X14Y127_CO6),
.O5(CLBLM_R_X11Y127_SLICE_X14Y127_AO5),
.O6(CLBLM_R_X11Y127_SLICE_X14Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y127_SLICE_X15Y127_AO6),
.Q(CLBLM_R_X11Y127_SLICE_X15Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333cccc33333c6c)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_DLUT (
.I0(CLBLM_L_X12Y127_SLICE_X17Y127_BO6),
.I1(CLBLM_R_X11Y127_SLICE_X15Y127_AQ),
.I2(CLBLM_L_X10Y127_SLICE_X13Y127_BQ),
.I3(CLBLM_L_X12Y127_SLICE_X16Y127_CO6),
.I4(CLBLM_L_X10Y129_SLICE_X13Y129_CO6),
.I5(CLBLM_R_X11Y128_SLICE_X14Y128_AO5),
.O5(CLBLM_R_X11Y127_SLICE_X15Y127_DO5),
.O6(CLBLM_R_X11Y127_SLICE_X15Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00bb008800bb0088)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_CLUT (
.I0(CLBLM_L_X12Y127_SLICE_X17Y127_BO6),
.I1(CLBLM_R_X11Y127_SLICE_X15Y127_AQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y128_SLICE_X14Y128_AO5),
.I4(CLBLM_L_X12Y127_SLICE_X16Y127_CO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y127_SLICE_X15Y127_CO5),
.O6(CLBLM_R_X11Y127_SLICE_X15Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h330033110f0f0f0e)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_BLUT (
.I0(CLBLM_R_X11Y128_SLICE_X15Y128_AQ),
.I1(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.I2(CLBLM_R_X11Y127_SLICE_X15Y127_CO6),
.I3(CLBLM_R_X11Y126_SLICE_X15Y126_BQ),
.I4(CLBLM_L_X10Y128_SLICE_X12Y128_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y127_SLICE_X15Y127_BO5),
.O6(CLBLM_R_X11Y127_SLICE_X15Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5c5c5c0c5c5c5c0)
  ) CLBLM_R_X11Y127_SLICE_X15Y127_ALUT (
.I0(CLBLM_R_X11Y127_SLICE_X15Y127_BO5),
.I1(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y127_SLICE_X15Y127_DO6),
.I4(CLBLM_R_X11Y130_SLICE_X14Y130_BO5),
.I5(1'b1),
.O5(CLBLM_R_X11Y127_SLICE_X15Y127_AO5),
.O6(CLBLM_R_X11Y127_SLICE_X15Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X10Y128_SLICE_X13Y128_BQ),
.Q(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.R(CLBLM_L_X8Y131_SLICE_X11Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000a0002000a000)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_DLUT (
.I0(CLBLM_L_X12Y127_SLICE_X16Y127_AQ),
.I1(CLBLM_R_X11Y128_SLICE_X15Y128_AQ),
.I2(CLBLM_R_X11Y129_SLICE_X14Y129_BQ),
.I3(CLBLM_R_X11Y129_SLICE_X14Y129_AQ),
.I4(CLBLM_L_X10Y128_SLICE_X12Y128_AQ),
.I5(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.O5(CLBLM_R_X11Y128_SLICE_X14Y128_DO5),
.O6(CLBLM_R_X11Y128_SLICE_X14Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0005a0002004a000)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_CLUT (
.I0(CLBLM_L_X12Y127_SLICE_X16Y127_AQ),
.I1(CLBLM_R_X11Y128_SLICE_X15Y128_AQ),
.I2(CLBLM_R_X11Y129_SLICE_X14Y129_BQ),
.I3(CLBLM_R_X11Y129_SLICE_X14Y129_AQ),
.I4(CLBLM_L_X10Y128_SLICE_X12Y128_AQ),
.I5(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.O5(CLBLM_R_X11Y128_SLICE_X14Y128_CO5),
.O6(CLBLM_R_X11Y128_SLICE_X14Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff51aeffff55aa)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_BLUT (
.I0(CLBLM_L_X10Y129_SLICE_X13Y129_CO6),
.I1(CLBLM_L_X10Y128_SLICE_X12Y128_CQ),
.I2(CLBLM_R_X11Y128_SLICE_X14Y128_AO5),
.I3(CLBLM_L_X10Y128_SLICE_X13Y128_AQ),
.I4(CLBLM_R_X11Y130_SLICE_X14Y130_BO5),
.I5(CLBLM_R_X11Y128_SLICE_X14Y128_CO6),
.O5(CLBLM_R_X11Y128_SLICE_X14Y128_BO5),
.O6(CLBLM_R_X11Y128_SLICE_X14Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f0f33773777)
  ) CLBLM_R_X11Y128_SLICE_X14Y128_ALUT (
.I0(CLBLM_R_X11Y129_SLICE_X15Y129_AO5),
.I1(CLBLM_L_X10Y125_SLICE_X13Y125_DO5),
.I2(CLBLM_L_X10Y128_SLICE_X12Y128_AQ),
.I3(CLBLM_R_X11Y126_SLICE_X14Y126_BQ),
.I4(CLBLM_R_X11Y128_SLICE_X15Y128_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y128_SLICE_X14Y128_AO5),
.O6(CLBLM_R_X11Y128_SLICE_X14Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y128_SLICE_X15Y128_AO6),
.Q(CLBLM_R_X11Y128_SLICE_X15Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000020200000200)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_DLUT (
.I0(CLBLM_L_X10Y128_SLICE_X12Y128_AQ),
.I1(CLBLM_R_X11Y129_SLICE_X14Y129_AQ),
.I2(CLBLM_L_X12Y127_SLICE_X16Y127_AQ),
.I3(CLBLM_R_X11Y128_SLICE_X15Y128_AQ),
.I4(CLBLM_R_X11Y129_SLICE_X14Y129_BQ),
.I5(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.O5(CLBLM_R_X11Y128_SLICE_X15Y128_DO5),
.O6(CLBLM_R_X11Y128_SLICE_X15Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0f0faf2f2)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_CLUT (
.I0(CLBLM_L_X10Y128_SLICE_X13Y128_BQ),
.I1(CLBLM_R_X11Y129_SLICE_X15Y129_CO6),
.I2(CLBLM_L_X10Y129_SLICE_X13Y129_CO6),
.I3(CLBLM_R_X11Y129_SLICE_X15Y129_DO6),
.I4(CLBLM_R_X11Y126_SLICE_X15Y126_AQ),
.I5(CLBLM_R_X11Y128_SLICE_X14Y128_AO5),
.O5(CLBLM_R_X11Y128_SLICE_X15Y128_CO5),
.O6(CLBLM_R_X11Y128_SLICE_X15Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a1e5a5a1e1e)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_BLUT (
.I0(CLBLM_L_X10Y129_SLICE_X13Y129_CO6),
.I1(CLBLM_L_X10Y126_SLICE_X13Y126_AQ),
.I2(CLBLM_R_X11Y126_SLICE_X15Y126_AQ),
.I3(CLBLM_R_X11Y129_SLICE_X15Y129_DO6),
.I4(CLBLM_R_X11Y128_SLICE_X14Y128_AO5),
.I5(CLBLM_R_X11Y129_SLICE_X15Y129_CO6),
.O5(CLBLM_R_X11Y128_SLICE_X15Y128_BO5),
.O6(CLBLM_R_X11Y128_SLICE_X15Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5fe050ef0f00000)
  ) CLBLM_R_X11Y128_SLICE_X15Y128_ALUT (
.I0(CLBLM_R_X11Y128_SLICE_X15Y128_AQ),
.I1(CLBLM_L_X10Y128_SLICE_X13Y128_CO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y129_SLICE_X15Y129_BO6),
.I4(CLBLM_R_X11Y123_SLICE_X15Y123_AQ),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_R_X11Y128_SLICE_X15Y128_AO5),
.O6(CLBLM_R_X11Y128_SLICE_X15Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y129_SLICE_X14Y129_AO6),
.Q(CLBLM_R_X11Y129_SLICE_X14Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y129_SLICE_X14Y129_BO6),
.Q(CLBLM_R_X11Y129_SLICE_X14Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555aaa65555aa6a)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_DLUT (
.I0(CLBLM_R_X11Y129_SLICE_X14Y129_BQ),
.I1(CLBLM_R_X11Y126_SLICE_X14Y126_DQ),
.I2(CLBLM_L_X12Y127_SLICE_X16Y127_AQ),
.I3(CLBLM_R_X11Y128_SLICE_X14Y128_AO5),
.I4(CLBLM_L_X10Y129_SLICE_X13Y129_CO6),
.I5(CLBLM_L_X10Y129_SLICE_X13Y129_BO5),
.O5(CLBLM_R_X11Y129_SLICE_X14Y129_DO5),
.O6(CLBLM_R_X11Y129_SLICE_X14Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffef0000dfff)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_CLUT (
.I0(CLBLM_R_X11Y129_SLICE_X14Y129_BQ),
.I1(CLBLM_R_X11Y128_SLICE_X14Y128_AO5),
.I2(CLBLM_L_X10Y126_SLICE_X13Y126_BQ),
.I3(CLBLM_L_X12Y127_SLICE_X16Y127_AQ),
.I4(CLBLM_L_X10Y129_SLICE_X13Y129_CO6),
.I5(CLBLM_L_X10Y129_SLICE_X13Y129_BO5),
.O5(CLBLM_R_X11Y129_SLICE_X14Y129_CO5),
.O6(CLBLM_R_X11Y129_SLICE_X14Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f40504f5f40504)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_BLUT (
.I0(CLBLM_R_X11Y127_SLICE_X15Y127_BO5),
.I1(CLBLM_R_X11Y130_SLICE_X14Y130_BO5),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y129_SLICE_X14Y129_DO6),
.I4(CLBLM_L_X10Y125_SLICE_X13Y125_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y129_SLICE_X14Y129_BO5),
.O6(CLBLM_R_X11Y129_SLICE_X14Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff005454ff004545)
  ) CLBLM_R_X11Y129_SLICE_X14Y129_ALUT (
.I0(CLBLM_R_X11Y127_SLICE_X15Y127_BO5),
.I1(CLBLM_R_X11Y130_SLICE_X14Y130_BO5),
.I2(CLBLM_R_X11Y129_SLICE_X14Y129_AQ),
.I3(CLBLM_L_X8Y129_SLICE_X11Y129_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y129_SLICE_X14Y129_CO6),
.O5(CLBLM_R_X11Y129_SLICE_X14Y129_AO5),
.O6(CLBLM_R_X11Y129_SLICE_X14Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfffffffffffffff)
  ) CLBLM_R_X11Y129_SLICE_X15Y129_DLUT (
.I0(CLBLM_R_X11Y129_SLICE_X14Y129_AQ),
.I1(CLBLM_L_X10Y129_SLICE_X13Y129_BO5),
.I2(CLBLM_L_X12Y126_SLICE_X16Y126_BQ),
.I3(CLBLM_L_X10Y128_SLICE_X13Y128_AQ),
.I4(CLBLM_L_X12Y127_SLICE_X16Y127_AQ),
.I5(CLBLM_R_X11Y129_SLICE_X14Y129_BQ),
.O5(CLBLM_R_X11Y129_SLICE_X15Y129_DO5),
.O6(CLBLM_R_X11Y129_SLICE_X15Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffeff)
  ) CLBLM_R_X11Y129_SLICE_X15Y129_CLUT (
.I0(CLBLM_R_X11Y129_SLICE_X14Y129_AQ),
.I1(CLBLM_L_X12Y127_SLICE_X16Y127_AQ),
.I2(CLBLM_L_X12Y126_SLICE_X16Y126_BQ),
.I3(CLBLM_L_X10Y129_SLICE_X13Y129_BO5),
.I4(CLBLM_L_X10Y128_SLICE_X13Y128_AQ),
.I5(CLBLM_R_X11Y129_SLICE_X14Y129_BQ),
.O5(CLBLM_R_X11Y129_SLICE_X15Y129_CO5),
.O6(CLBLM_R_X11Y129_SLICE_X15Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8060f0f080608060)
  ) CLBLM_R_X11Y129_SLICE_X15Y129_BLUT (
.I0(CLBLM_R_X11Y128_SLICE_X15Y128_AQ),
.I1(CLBLM_L_X10Y128_SLICE_X12Y128_AQ),
.I2(CLBLM_R_X11Y127_SLICE_X15Y127_CO5),
.I3(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.I4(CLBLM_R_X11Y130_SLICE_X14Y130_AQ),
.I5(CLBLM_R_X11Y129_SLICE_X15Y129_AO5),
.O5(CLBLM_R_X11Y129_SLICE_X15Y129_BO5),
.O6(CLBLM_R_X11Y129_SLICE_X15Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000400044004400)
  ) CLBLM_R_X11Y129_SLICE_X15Y129_ALUT (
.I0(CLBLM_L_X8Y129_SLICE_X11Y129_BQ),
.I1(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.I2(CLBLM_R_X11Y127_SLICE_X15Y127_CO5),
.I3(CLBLM_R_X11Y126_SLICE_X15Y126_BQ),
.I4(CLBLM_R_X11Y130_SLICE_X14Y130_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y129_SLICE_X15Y129_AO5),
.O6(CLBLM_R_X11Y129_SLICE_X15Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y130_SLICE_X14Y130_AO6),
.Q(CLBLM_R_X11Y130_SLICE_X14Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y130_SLICE_X14Y130_DO5),
.O6(CLBLM_R_X11Y130_SLICE_X14Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y130_SLICE_X14Y130_CO5),
.O6(CLBLM_R_X11Y130_SLICE_X14Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h303000058ac5aaf0)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_BLUT (
.I0(CLBLM_R_X11Y128_SLICE_X15Y128_AQ),
.I1(CLBLM_L_X8Y129_SLICE_X11Y129_BQ),
.I2(CLBLM_L_X10Y129_SLICE_X12Y129_AQ),
.I3(CLBLM_L_X10Y128_SLICE_X12Y128_AQ),
.I4(CLBLM_R_X11Y126_SLICE_X15Y126_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y130_SLICE_X14Y130_BO5),
.O6(CLBLM_R_X11Y130_SLICE_X14Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfafaccccaafa)
  ) CLBLM_R_X11Y130_SLICE_X14Y130_ALUT (
.I0(CLBLM_R_X11Y129_SLICE_X15Y129_AO6),
.I1(CLBLM_R_X7Y126_SLICE_X8Y126_BQ),
.I2(CLBLM_R_X11Y130_SLICE_X14Y130_AQ),
.I3(CLBLM_R_X11Y130_SLICE_X14Y130_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y127_SLICE_X15Y127_BO5),
.O5(CLBLM_R_X11Y130_SLICE_X14Y130_AO5),
.O6(CLBLM_R_X11Y130_SLICE_X14Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y130_SLICE_X15Y130_DO5),
.O6(CLBLM_R_X11Y130_SLICE_X15Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y130_SLICE_X15Y130_CO5),
.O6(CLBLM_R_X11Y130_SLICE_X15Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y130_SLICE_X15Y130_BO5),
.O6(CLBLM_R_X11Y130_SLICE_X15Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y130_SLICE_X15Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y130_SLICE_X15Y130_AO5),
.O6(CLBLM_R_X11Y130_SLICE_X15Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_DO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_CO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_BO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_AO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y131_SLICE_X15Y131_AO6),
.Q(CLBLM_R_X11Y131_SLICE_X15Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_DO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_CO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_BO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfb51fa50fb51fa50)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.I2(CLBLM_R_X11Y131_SLICE_X15Y131_AQ),
.I3(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.I4(RIOB33_X105Y141_IOB_X1Y142_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_AO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y151_SLICE_X14Y151_DO5),
.O6(CLBLM_R_X11Y151_SLICE_X14Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y151_SLICE_X14Y151_CO5),
.O6(CLBLM_R_X11Y151_SLICE_X14Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y151_SLICE_X14Y151_BO5),
.O6(CLBLM_R_X11Y151_SLICE_X14Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0f)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X11Y124_SLICE_X14Y124_A5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y151_SLICE_X14Y151_AO5),
.O6(CLBLM_R_X11Y151_SLICE_X14Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y151_SLICE_X15Y151_DO5),
.O6(CLBLM_R_X11Y151_SLICE_X15Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y151_SLICE_X15Y151_CO5),
.O6(CLBLM_R_X11Y151_SLICE_X15Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y151_SLICE_X15Y151_BO5),
.O6(CLBLM_R_X11Y151_SLICE_X15Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y151_SLICE_X15Y151_AO5),
.O6(CLBLM_R_X11Y151_SLICE_X15Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y127_SLICE_X18Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y127_SLICE_X18Y127_AO6),
.Q(CLBLM_R_X13Y127_SLICE_X18Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y127_SLICE_X18Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y127_SLICE_X18Y127_DO5),
.O6(CLBLM_R_X13Y127_SLICE_X18Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y127_SLICE_X18Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y127_SLICE_X18Y127_CO5),
.O6(CLBLM_R_X13Y127_SLICE_X18Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y127_SLICE_X18Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y127_SLICE_X18Y127_BO5),
.O6(CLBLM_R_X13Y127_SLICE_X18Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f3f003030300)
  ) CLBLM_R_X13Y127_SLICE_X18Y127_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y127_SLICE_X15Y127_BO5),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y127_SLICE_X17Y127_AO6),
.I4(CLBLM_R_X11Y130_SLICE_X14Y130_BO5),
.I5(CLBLM_R_X11Y120_SLICE_X14Y120_CQ),
.O5(CLBLM_R_X13Y127_SLICE_X18Y127_AO5),
.O6(CLBLM_R_X13Y127_SLICE_X18Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y127_SLICE_X19Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y127_SLICE_X19Y127_DO5),
.O6(CLBLM_R_X13Y127_SLICE_X19Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y127_SLICE_X19Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y127_SLICE_X19Y127_CO5),
.O6(CLBLM_R_X13Y127_SLICE_X19Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y127_SLICE_X19Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y127_SLICE_X19Y127_BO5),
.O6(CLBLM_R_X13Y127_SLICE_X19Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y127_SLICE_X19Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y127_SLICE_X19Y127_AO5),
.O6(CLBLM_R_X13Y127_SLICE_X19Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y140_SLICE_X162Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y140_SLICE_X162Y140_DO5),
.O6(CLBLM_R_X103Y140_SLICE_X162Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y140_SLICE_X162Y140_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y140_SLICE_X162Y140_CO5),
.O6(CLBLM_R_X103Y140_SLICE_X162Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y140_SLICE_X162Y140_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y140_SLICE_X162Y140_BO5),
.O6(CLBLM_R_X103Y140_SLICE_X162Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y140_SLICE_X162Y140_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y140_SLICE_X162Y140_AO5),
.O6(CLBLM_R_X103Y140_SLICE_X162Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y140_SLICE_X163Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y140_SLICE_X163Y140_DO5),
.O6(CLBLM_R_X103Y140_SLICE_X163Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y140_SLICE_X163Y140_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y140_SLICE_X163Y140_CO5),
.O6(CLBLM_R_X103Y140_SLICE_X163Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y140_SLICE_X163Y140_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y140_SLICE_X163Y140_BO5),
.O6(CLBLM_R_X103Y140_SLICE_X163Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0000088008800)
  ) CLBLM_R_X103Y140_SLICE_X163Y140_ALUT (
.I0(RIOB33_X105Y141_IOB_X1Y141_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(RIOB33_X105Y137_IOB_X1Y138_I),
.I3(RIOB33_X105Y139_IOB_X1Y140_I),
.I4(RIOB33_X105Y139_IOB_X1Y139_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y140_SLICE_X163Y140_AO5),
.O6(CLBLM_R_X103Y140_SLICE_X163Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_DO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_CO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_BO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_AO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_DO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_CO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_BO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fffff0f0ffff)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_AO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y171_SLICE_X162Y171_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y171_SLICE_X162Y171_DO5),
.O6(CLBLM_R_X103Y171_SLICE_X162Y171_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y171_SLICE_X162Y171_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y171_SLICE_X162Y171_CO5),
.O6(CLBLM_R_X103Y171_SLICE_X162Y171_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y171_SLICE_X162Y171_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y171_SLICE_X162Y171_BO5),
.O6(CLBLM_R_X103Y171_SLICE_X162Y171_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y171_SLICE_X162Y171_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y171_SLICE_X162Y171_AO5),
.O6(CLBLM_R_X103Y171_SLICE_X162Y171_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y171_SLICE_X163Y171_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y171_SLICE_X163Y171_DO5),
.O6(CLBLM_R_X103Y171_SLICE_X163Y171_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y171_SLICE_X163Y171_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y171_SLICE_X163Y171_CO5),
.O6(CLBLM_R_X103Y171_SLICE_X163Y171_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddddddf5f5f5f5)
  ) CLBLM_R_X103Y171_SLICE_X163Y171_BLUT (
.I0(RIOB33_X105Y143_IOB_X1Y143_I),
.I1(CLBLM_L_X12Y126_SLICE_X16Y126_AQ),
.I2(CLBLM_L_X8Y126_SLICE_X10Y126_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y171_SLICE_X163Y171_BO5),
.O6(CLBLM_R_X103Y171_SLICE_X163Y171_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaffffff00ffff)
  ) CLBLM_R_X103Y171_SLICE_X163Y171_ALUT (
.I0(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y171_SLICE_X163Y171_AO5),
.O6(CLBLM_R_X103Y171_SLICE_X163Y171_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y173_SLICE_X162Y173_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y173_SLICE_X162Y173_DO5),
.O6(CLBLM_R_X103Y173_SLICE_X162Y173_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y173_SLICE_X162Y173_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y173_SLICE_X162Y173_CO5),
.O6(CLBLM_R_X103Y173_SLICE_X162Y173_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y173_SLICE_X162Y173_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y173_SLICE_X162Y173_BO5),
.O6(CLBLM_R_X103Y173_SLICE_X162Y173_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y173_SLICE_X162Y173_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y173_SLICE_X162Y173_AO5),
.O6(CLBLM_R_X103Y173_SLICE_X162Y173_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y173_SLICE_X163Y173_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y173_SLICE_X163Y173_DO5),
.O6(CLBLM_R_X103Y173_SLICE_X163Y173_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y173_SLICE_X163Y173_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y173_SLICE_X163Y173_CO5),
.O6(CLBLM_R_X103Y173_SLICE_X163Y173_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y173_SLICE_X163Y173_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y173_SLICE_X163Y173_BO5),
.O6(CLBLM_R_X103Y173_SLICE_X163Y173_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaffffff00ffff)
  ) CLBLM_R_X103Y173_SLICE_X163Y173_ALUT (
.I0(CLBLM_L_X12Y121_SLICE_X16Y121_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X11Y131_SLICE_X15Y131_AQ),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y173_SLICE_X163Y173_AO5),
.O6(CLBLM_R_X103Y173_SLICE_X163Y173_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y175_SLICE_X162Y175_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y175_SLICE_X162Y175_DO5),
.O6(CLBLM_R_X103Y175_SLICE_X162Y175_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y175_SLICE_X162Y175_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y175_SLICE_X162Y175_CO5),
.O6(CLBLM_R_X103Y175_SLICE_X162Y175_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y175_SLICE_X162Y175_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y175_SLICE_X162Y175_BO5),
.O6(CLBLM_R_X103Y175_SLICE_X162Y175_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y175_SLICE_X162Y175_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y175_SLICE_X162Y175_AO5),
.O6(CLBLM_R_X103Y175_SLICE_X162Y175_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y175_SLICE_X163Y175_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y175_SLICE_X163Y175_DO5),
.O6(CLBLM_R_X103Y175_SLICE_X163Y175_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y175_SLICE_X163Y175_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y175_SLICE_X163Y175_CO5),
.O6(CLBLM_R_X103Y175_SLICE_X163Y175_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y175_SLICE_X163Y175_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y175_SLICE_X163Y175_BO5),
.O6(CLBLM_R_X103Y175_SLICE_X163Y175_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffccffcc)
  ) CLBLM_R_X103Y175_SLICE_X163Y175_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y127_IOB_X1Y128_I),
.I2(1'b1),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(1'b1),
.I5(RIOB33_X105Y129_IOB_X1Y130_I),
.O5(CLBLM_R_X103Y175_SLICE_X163Y175_AO5),
.O6(CLBLM_R_X103Y175_SLICE_X163Y175_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_DO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_CO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_BO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_AO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_DO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_CO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_BO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0f0fff0fff0f)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y143_IOB_X1Y143_I),
.I3(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.I4(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_AO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(LIOB33_X0Y77_IOB_X0Y78_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y51_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y51_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y51_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y52_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y52_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y53_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y53_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y53_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y54_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y54_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y55_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y55_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y56_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y56_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y57_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y57_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y57_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y58_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y58_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y59_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y59_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y60_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y60_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y61_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y61_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y62_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y62_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y63_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y63_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y64_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y64_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y64_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y65_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y65_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y65_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y66_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y66_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y66_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y67_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y67_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y67_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y68_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y68_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y68_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y69_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y69_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y69_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y70_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y70_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y70_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y71_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y71_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y71_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y72_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y72_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y72_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y73_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y73_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y73_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y74_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y74_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y74_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y75_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y75_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y75_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y76_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y76_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y76_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y77_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y77_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y77_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y78_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y78_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y78_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y79_IOB_X0Y79_IBUF (
.I(LIOB33_X0Y79_IOB_X0Y79_IPAD),
.O(LIOB33_X0Y79_IOB_X0Y79_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y79_IOB_X0Y80_OBUF (
.I(CLBLL_L_X2Y117_SLICE_X0Y117_AO6),
.O(LIOB33_X0Y79_IOB_X0Y80_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y101_OBUF (
.I(CLBLL_L_X2Y118_SLICE_X0Y118_AO5),
.O(LIOB33_X0Y101_IOB_X0Y101_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y102_OBUF (
.I(CLBLL_L_X2Y117_SLICE_X0Y117_BO6),
.O(LIOB33_X0Y101_IOB_X0Y102_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y103_OBUF (
.I(CLBLL_L_X2Y125_SLICE_X1Y125_CO6),
.O(LIOB33_X0Y103_IOB_X0Y103_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y104_OBUF (
.I(CLBLL_L_X2Y117_SLICE_X0Y117_AO5),
.O(LIOB33_X0Y103_IOB_X0Y104_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y105_OBUF (
.I(CLBLL_L_X2Y117_SLICE_X0Y117_CO6),
.O(LIOB33_X0Y105_IOB_X0Y105_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y106_OBUF (
.I(CLBLL_L_X2Y117_SLICE_X0Y117_CO5),
.O(LIOB33_X0Y105_IOB_X0Y106_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y107_OBUF (
.I(CLBLL_L_X2Y115_SLICE_X0Y115_AO5),
.O(LIOB33_X0Y107_IOB_X0Y107_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y108_OBUF (
.I(CLBLL_L_X2Y117_SLICE_X0Y117_BO5),
.O(LIOB33_X0Y107_IOB_X0Y108_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y109_OBUF (
.I(CLBLL_L_X2Y118_SLICE_X1Y118_CO5),
.O(LIOB33_X0Y109_IOB_X0Y109_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y110_OBUF (
.I(CLBLL_L_X2Y115_SLICE_X0Y115_AO6),
.O(LIOB33_X0Y109_IOB_X0Y110_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y111_OBUF (
.I(1'b0),
.O(LIOB33_X0Y111_IOB_X0Y111_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y112_OBUF (
.I(CLBLM_L_X10Y121_SLICE_X13Y121_B5Q),
.O(LIOB33_X0Y111_IOB_X0Y112_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y113_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_I),
.O(LIOB33_X0Y113_IOB_X0Y113_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y114_OBUF (
.I(CLBLL_L_X4Y118_SLICE_X5Y118_CQ),
.O(LIOB33_X0Y113_IOB_X0Y114_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y115_OBUF (
.I(CLBLM_L_X10Y121_SLICE_X13Y121_BQ),
.O(LIOB33_X0Y115_IOB_X0Y115_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y116_OBUF (
.I(CLBLM_R_X5Y128_SLICE_X7Y128_BQ),
.O(LIOB33_X0Y115_IOB_X0Y116_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y117_OBUF (
.I(CLBLL_L_X2Y122_SLICE_X1Y122_AQ),
.O(LIOB33_X0Y117_IOB_X0Y117_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y118_OBUF (
.I(CLBLL_L_X4Y122_SLICE_X5Y122_CQ),
.O(LIOB33_X0Y117_IOB_X0Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUF (
.I(CLBLM_L_X8Y122_SLICE_X10Y122_AQ),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUF (
.I(CLBLM_L_X10Y120_SLICE_X13Y120_AQ),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUF (
.I(CLBLM_R_X5Y128_SLICE_X7Y128_B5Q),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUF (
.I(CLBLM_R_X5Y126_SLICE_X7Y126_AQ),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUF (
.I(CLBLL_L_X4Y118_SLICE_X5Y118_C5Q),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(CLBLL_L_X4Y122_SLICE_X5Y122_C5Q),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y125_OBUF (
.I(CLBLM_L_X8Y123_SLICE_X10Y123_C5Q),
.O(LIOB33_X0Y125_IOB_X0Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y126_OBUF (
.I(CLBLM_R_X3Y125_SLICE_X2Y125_AQ),
.O(LIOB33_X0Y125_IOB_X0Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y127_OBUF (
.I(CLBLL_L_X4Y126_SLICE_X4Y126_AQ),
.O(LIOB33_X0Y127_IOB_X0Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y128_OBUF (
.I(CLBLL_L_X2Y118_SLICE_X1Y118_B5Q),
.O(LIOB33_X0Y127_IOB_X0Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y129_OBUF (
.I(CLBLM_R_X3Y123_SLICE_X3Y123_CQ),
.O(LIOB33_X0Y129_IOB_X0Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y130_OBUF (
.I(CLBLL_L_X52Y126_SLICE_X78Y126_AO6),
.O(LIOB33_X0Y129_IOB_X0Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y131_OBUF (
.I(CLBLM_R_X5Y118_SLICE_X6Y118_AO5),
.O(LIOB33_X0Y131_IOB_X0Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y132_OBUF (
.I(CLBLM_R_X5Y118_SLICE_X6Y118_AQ),
.O(LIOB33_X0Y131_IOB_X0Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y133_OBUF (
.I(CLBLM_R_X3Y132_SLICE_X2Y132_A5Q),
.O(LIOB33_X0Y133_IOB_X0Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y134_OBUF (
.I(CLBLM_R_X3Y123_SLICE_X2Y123_CQ),
.O(LIOB33_X0Y133_IOB_X0Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y135_OBUF (
.I(CLBLM_R_X3Y129_SLICE_X2Y129_AQ),
.O(LIOB33_X0Y135_IOB_X0Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUF (
.I(CLBLM_R_X3Y132_SLICE_X2Y132_BQ),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUF (
.I(CLBLM_R_X3Y131_SLICE_X2Y131_AQ),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUF (
.I(CLBLM_R_X3Y131_SLICE_X2Y131_BQ),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUF (
.I(CLBLM_R_X3Y132_SLICE_X2Y132_AQ),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUF (
.I(CLBLL_L_X2Y125_SLICE_X1Y125_AQ),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y141_OBUF (
.I(CLBLL_L_X2Y126_SLICE_X1Y126_AQ),
.O(LIOB33_X0Y141_IOB_X0Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y142_OBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_I),
.O(LIOB33_X0Y141_IOB_X0Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y143_IOB_X0Y143_OBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_I),
.O(LIOB33_X0Y143_IOB_X0Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y145_OBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_I),
.O(LIOB33_X0Y145_IOB_X0Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y146_OBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_I),
.O(LIOB33_X0Y145_IOB_X0Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y147_OBUF (
.I(LIOB33_X0Y71_IOB_X0Y71_I),
.O(LIOB33_X0Y147_IOB_X0Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y148_OBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_I),
.O(LIOB33_X0Y147_IOB_X0Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y151_OBUF (
.I(LIOB33_X0Y65_IOB_X0Y65_I),
.O(LIOB33_X0Y151_IOB_X0Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y152_OBUF (
.I(LIOB33_X0Y65_IOB_X0Y66_I),
.O(LIOB33_X0Y151_IOB_X0Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y153_OBUF (
.I(LIOB33_X0Y67_IOB_X0Y67_I),
.O(LIOB33_X0Y153_IOB_X0Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y154_OBUF (
.I(LIOB33_X0Y67_IOB_X0Y68_I),
.O(LIOB33_X0Y153_IOB_X0Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y155_OBUF (
.I(LIOB33_X0Y69_IOB_X0Y70_I),
.O(LIOB33_X0Y155_IOB_X0Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y156_OBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_I),
.O(LIOB33_X0Y155_IOB_X0Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y157_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_I),
.O(LIOB33_X0Y157_IOB_X0Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y158_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_I),
.O(LIOB33_X0Y157_IOB_X0Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y159_OBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_I),
.O(LIOB33_X0Y159_IOB_X0Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y160_OBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_I),
.O(LIOB33_X0Y159_IOB_X0Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y161_OBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_I),
.O(LIOB33_X0Y161_IOB_X0Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y162_OBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_I),
.O(LIOB33_X0Y161_IOB_X0Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y163_OBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_I),
.O(LIOB33_X0Y163_IOB_X0Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y164_OBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_I),
.O(LIOB33_X0Y163_IOB_X0Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y165_OBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_I),
.O(LIOB33_X0Y165_IOB_X0Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y166_OBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_I),
.O(LIOB33_X0Y165_IOB_X0Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y167_OBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_I),
.O(LIOB33_X0Y167_IOB_X0Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y168_OBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_I),
.O(LIOB33_X0Y167_IOB_X0Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y169_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_I),
.O(LIOB33_X0Y169_IOB_X0Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y170_OBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.O(LIOB33_X0Y169_IOB_X0Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y171_OBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.O(LIOB33_X0Y171_IOB_X0Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y172_OBUF (
.I(CLBLM_R_X103Y140_SLICE_X163Y140_AO6),
.O(LIOB33_X0Y171_IOB_X0Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y173_OBUF (
.I(CLBLM_R_X103Y140_SLICE_X163Y140_AO5),
.O(LIOB33_X0Y173_IOB_X0Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y174_OBUF (
.I(CLBLM_R_X11Y151_SLICE_X14Y151_AO6),
.O(LIOB33_X0Y173_IOB_X0Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y175_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_I),
.O(LIOB33_X0Y175_IOB_X0Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y176_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_I),
.O(LIOB33_X0Y175_IOB_X0Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y177_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_I),
.O(LIOB33_X0Y177_IOB_X0Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y178_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_I),
.O(LIOB33_X0Y177_IOB_X0Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y179_OBUF (
.I(RIOB33_X105Y131_IOB_X1Y131_I),
.O(LIOB33_X0Y179_IOB_X0Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y180_OBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_I),
.O(LIOB33_X0Y179_IOB_X0Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y181_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_I),
.O(LIOB33_X0Y181_IOB_X0Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y182_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_I),
.O(LIOB33_X0Y181_IOB_X0Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y183_OBUF (
.I(RIOB33_X105Y135_IOB_X1Y135_I),
.O(LIOB33_X0Y183_IOB_X0Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y184_OBUF (
.I(RIOB33_X105Y135_IOB_X1Y136_I),
.O(LIOB33_X0Y183_IOB_X0Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y185_OBUF (
.I(RIOB33_X105Y137_IOB_X1Y137_I),
.O(LIOB33_X0Y185_IOB_X0Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y186_OBUF (
.I(RIOB33_X105Y143_IOB_X1Y143_I),
.O(LIOB33_X0Y185_IOB_X0Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y187_OBUF (
.I(RIOB33_X105Y143_IOB_X1Y144_I),
.O(LIOB33_X0Y187_IOB_X0Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y188_OBUF (
.I(RIOB33_X105Y145_IOB_X1Y145_I),
.O(LIOB33_X0Y187_IOB_X0Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y189_OBUF (
.I(RIOB33_X105Y145_IOB_X1Y146_I),
.O(LIOB33_X0Y189_IOB_X0Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y190_OBUF (
.I(RIOB33_X105Y147_IOB_X1Y147_I),
.O(LIOB33_X0Y189_IOB_X0Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y191_OBUF (
.I(RIOB33_X105Y147_IOB_X1Y148_I),
.O(LIOB33_X0Y191_IOB_X0Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y192_OBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_I),
.O(LIOB33_X0Y191_IOB_X0Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y193_OBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_I),
.O(LIOB33_X0Y193_IOB_X0Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y194_OBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_I),
.O(LIOB33_X0Y193_IOB_X0Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y195_OBUF (
.I(LIOB33_X0Y63_IOB_X0Y64_I),
.O(LIOB33_X0Y195_IOB_X0Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y196_OBUF (
.I(LIOB33_X0Y69_IOB_X0Y69_I),
.O(LIOB33_X0Y195_IOB_X0Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y197_OBUF (
.I(LIOB33_X0Y71_IOB_X0Y72_I),
.O(LIOB33_X0Y197_IOB_X0Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y198_OBUF (
.I(LIOB33_X0Y73_IOB_X0Y73_I),
.O(LIOB33_X0Y197_IOB_X0Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y50_IOB_X0Y50_IBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_IPAD),
.O(LIOB33_SING_X0Y50_IOB_X0Y50_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y100_IOB_X0Y100_OBUF (
.I(CLBLL_L_X2Y118_SLICE_X0Y118_AO6),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_OBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_I),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y150_IOB_X0Y150_OBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_I),
.O(LIOB33_SING_X0Y150_IOB_X0Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y199_IOB_X0Y199_OBUF (
.I(LIOB33_X0Y73_IOB_X0Y74_I),
.O(LIOB33_SING_X0Y199_IOB_X0Y199_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y101_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y102_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y103_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y104_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y105_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y105_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y106_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y107_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y108_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y109_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y110_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y111_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y112_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y113_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y114_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y115_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y116_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y117_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y118_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y118_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y119_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y119_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y120_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y121_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y122_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y123_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y124_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y124_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y125_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y126_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y127_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y128_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y129_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y129_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y130_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y130_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y131_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y131_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y131_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y132_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y132_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y133_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y133_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y134_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y134_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y135_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y135_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y135_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y136_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y136_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y136_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y137_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y137_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y137_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y138_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y138_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y138_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y139_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y139_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y139_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y140_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y140_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y140_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y141_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y141_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y141_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y142_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y142_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y142_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y143_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y143_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y143_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y144_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y144_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y144_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y145_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y145_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y145_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y146_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y146_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y146_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y147_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y147_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y147_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y148_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y148_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y151_OBUF (
.I(LIOB33_X0Y75_IOB_X0Y76_I),
.O(RIOB33_X105Y151_IOB_X1Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y152_OBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O(RIOB33_X105Y151_IOB_X1Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y153_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_I),
.O(RIOB33_X105Y153_IOB_X1Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y154_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_I),
.O(RIOB33_X105Y153_IOB_X1Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y155_OBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_I),
.O(RIOB33_X105Y155_IOB_X1Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y156_OBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_I),
.O(RIOB33_X105Y155_IOB_X1Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y157_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_I),
.O(RIOB33_X105Y157_IOB_X1Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y158_OBUF (
.I(CLBLL_L_X36Y124_SLICE_X54Y124_AO6),
.O(RIOB33_X105Y157_IOB_X1Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y159_OBUF (
.I(CLBLM_R_X11Y124_SLICE_X14Y124_DO6),
.O(RIOB33_X105Y159_IOB_X1Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y160_OBUF (
.I(CLBLM_R_X11Y124_SLICE_X14Y124_DO5),
.O(RIOB33_X105Y159_IOB_X1Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y161_OBUF (
.I(CLBLM_L_X10Y126_SLICE_X12Y126_DO6),
.O(RIOB33_X105Y161_IOB_X1Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y162_OBUF (
.I(CLBLM_L_X10Y126_SLICE_X12Y126_DO5),
.O(RIOB33_X105Y161_IOB_X1Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y163_OBUF (
.I(CLBLM_L_X10Y123_SLICE_X13Y123_DO6),
.O(RIOB33_X105Y163_IOB_X1Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y164_OBUF (
.I(CLBLM_L_X10Y123_SLICE_X13Y123_DO5),
.O(RIOB33_X105Y163_IOB_X1Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y165_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_I),
.O(RIOB33_X105Y165_IOB_X1Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y166_OBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.O(RIOB33_X105Y165_IOB_X1Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y167_OBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.O(RIOB33_X105Y167_IOB_X1Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y168_OBUF (
.I(CLBLM_R_X11Y151_SLICE_X14Y151_AO6),
.O(RIOB33_X105Y167_IOB_X1Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y169_OBUF (
.I(CLBLM_R_X103Y169_SLICE_X163Y169_AO6),
.O(RIOB33_X105Y169_IOB_X1Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y170_OBUF (
.I(CLBLM_R_X103Y171_SLICE_X163Y171_AO6),
.O(RIOB33_X105Y169_IOB_X1Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y171_OBUF (
.I(CLBLM_R_X103Y171_SLICE_X163Y171_AO5),
.O(RIOB33_X105Y171_IOB_X1Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y172_OBUF (
.I(CLBLM_R_X103Y171_SLICE_X163Y171_BO6),
.O(RIOB33_X105Y171_IOB_X1Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y173_OBUF (
.I(CLBLM_R_X103Y171_SLICE_X163Y171_BO5),
.O(RIOB33_X105Y173_IOB_X1Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y174_OBUF (
.I(CLBLM_R_X103Y173_SLICE_X163Y173_AO6),
.O(RIOB33_X105Y173_IOB_X1Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y175_OBUF (
.I(CLBLM_L_X10Y136_SLICE_X12Y136_BO6),
.O(RIOB33_X105Y175_IOB_X1Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y176_OBUF (
.I(CLBLM_R_X103Y173_SLICE_X163Y173_AO5),
.O(RIOB33_X105Y175_IOB_X1Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y177_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_AO6),
.O(RIOB33_X105Y177_IOB_X1Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y178_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_AO5),
.O(RIOB33_X105Y177_IOB_X1Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y179_OBUF (
.I(CLBLM_L_X10Y136_SLICE_X12Y136_AO5),
.O(RIOB33_X105Y179_IOB_X1Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y180_OBUF (
.I(CLBLM_R_X11Y124_SLICE_X14Y124_DO6),
.O(RIOB33_X105Y179_IOB_X1Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y181_OBUF (
.I(CLBLM_R_X11Y124_SLICE_X14Y124_DO5),
.O(RIOB33_X105Y181_IOB_X1Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y182_OBUF (
.I(CLBLM_L_X10Y126_SLICE_X12Y126_DO6),
.O(RIOB33_X105Y181_IOB_X1Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y183_OBUF (
.I(CLBLM_L_X10Y126_SLICE_X12Y126_DO5),
.O(RIOB33_X105Y183_IOB_X1Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y184_OBUF (
.I(CLBLM_L_X10Y123_SLICE_X13Y123_DO6),
.O(RIOB33_X105Y183_IOB_X1Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y185_OBUF (
.I(CLBLM_L_X10Y123_SLICE_X13Y123_DO5),
.O(RIOB33_X105Y185_IOB_X1Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y186_OBUF (
.I(CLBLM_R_X11Y125_SLICE_X14Y125_AQ),
.O(RIOB33_X105Y185_IOB_X1Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y187_OBUF (
.I(CLBLM_L_X10Y124_SLICE_X12Y124_AQ),
.O(RIOB33_X105Y187_IOB_X1Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y188_OBUF (
.I(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.O(RIOB33_X105Y187_IOB_X1Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y189_OBUF (
.I(CLBLM_L_X8Y129_SLICE_X10Y129_AQ),
.O(RIOB33_X105Y189_IOB_X1Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y190_OBUF (
.I(CLBLM_L_X12Y126_SLICE_X16Y126_AQ),
.O(RIOB33_X105Y189_IOB_X1Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y191_OBUF (
.I(CLBLM_L_X8Y126_SLICE_X10Y126_AQ),
.O(RIOB33_X105Y191_IOB_X1Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y192_OBUF (
.I(CLBLM_L_X12Y121_SLICE_X16Y121_BQ),
.O(RIOB33_X105Y191_IOB_X1Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y193_OBUF (
.I(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.O(RIOB33_X105Y193_IOB_X1Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y194_OBUF (
.I(CLBLM_R_X11Y131_SLICE_X15Y131_AQ),
.O(RIOB33_X105Y193_IOB_X1Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y195_OBUF (
.I(CLBLM_R_X11Y128_SLICE_X14Y128_AQ),
.O(RIOB33_X105Y195_IOB_X1Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y196_OBUF (
.I(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.O(RIOB33_X105Y195_IOB_X1Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y197_OBUF (
.I(CLBLM_R_X103Y175_SLICE_X163Y175_AO6),
.O(RIOB33_X105Y197_IOB_X1Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y198_OBUF (
.I(CLBLM_R_X103Y175_SLICE_X163Y175_AO6),
.O(RIOB33_X105Y197_IOB_X1Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y100_IOB_X1Y100_IBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_IPAD),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y149_IOB_X1Y149_IBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_IPAD),
.O(RIOB33_SING_X105Y149_IOB_X1Y149_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y150_IOB_X1Y150_OBUF (
.I(LIOB33_X0Y75_IOB_X0Y75_I),
.O(RIOB33_SING_X105Y150_IOB_X1Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y199_IOB_X1Y199_OBUF (
.I(CLBLM_R_X11Y131_SLICE_X15Y131_AQ),
.O(RIOB33_SING_X105Y199_IOB_X1Y199_OPAD)
  );
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B = CLBLL_L_X2Y115_SLICE_X0Y115_BO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C = CLBLL_L_X2Y115_SLICE_X0Y115_CO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D = CLBLL_L_X2Y115_SLICE_X0Y115_DO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_AMUX = CLBLL_L_X2Y115_SLICE_X0Y115_AO5;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A = CLBLL_L_X2Y115_SLICE_X1Y115_AO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B = CLBLL_L_X2Y115_SLICE_X1Y115_BO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C = CLBLL_L_X2Y115_SLICE_X1Y115_CO6;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D = CLBLL_L_X2Y115_SLICE_X1Y115_DO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A = CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B = CLBLL_L_X2Y117_SLICE_X0Y117_BO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C = CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D = CLBLL_L_X2Y117_SLICE_X0Y117_DO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_AMUX = CLBLL_L_X2Y117_SLICE_X0Y117_AO5;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_BMUX = CLBLL_L_X2Y117_SLICE_X0Y117_BO5;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_CMUX = CLBLL_L_X2Y117_SLICE_X0Y117_CO5;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A = CLBLL_L_X2Y117_SLICE_X1Y117_AO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B = CLBLL_L_X2Y117_SLICE_X1Y117_BO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C = CLBLL_L_X2Y117_SLICE_X1Y117_CO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D = CLBLL_L_X2Y117_SLICE_X1Y117_DO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B = CLBLL_L_X2Y118_SLICE_X0Y118_BO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C = CLBLL_L_X2Y118_SLICE_X0Y118_CO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D = CLBLL_L_X2Y118_SLICE_X0Y118_DO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_AMUX = CLBLL_L_X2Y118_SLICE_X0Y118_AO5;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A = CLBLL_L_X2Y118_SLICE_X1Y118_AO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B = CLBLL_L_X2Y118_SLICE_X1Y118_BO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C = CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D = CLBLL_L_X2Y118_SLICE_X1Y118_DO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_AMUX = CLBLL_L_X2Y118_SLICE_X1Y118_A5Q;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_BMUX = CLBLL_L_X2Y118_SLICE_X1Y118_B5Q;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_CMUX = CLBLL_L_X2Y118_SLICE_X1Y118_CO5;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A = CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B = CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C = CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D = CLBLL_L_X2Y119_SLICE_X0Y119_DO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_DMUX = CLBLL_L_X2Y119_SLICE_X0Y119_DO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A = CLBLL_L_X2Y119_SLICE_X1Y119_AO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B = CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C = CLBLL_L_X2Y119_SLICE_X1Y119_CO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D = CLBLL_L_X2Y119_SLICE_X1Y119_DO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A = CLBLL_L_X2Y120_SLICE_X0Y120_AO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B = CLBLL_L_X2Y120_SLICE_X0Y120_BO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C = CLBLL_L_X2Y120_SLICE_X0Y120_CO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D = CLBLL_L_X2Y120_SLICE_X0Y120_DO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A = CLBLL_L_X2Y120_SLICE_X1Y120_AO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B = CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C = CLBLL_L_X2Y120_SLICE_X1Y120_CO6;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D = CLBLL_L_X2Y120_SLICE_X1Y120_DO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A = CLBLL_L_X2Y121_SLICE_X0Y121_AO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B = CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C = CLBLL_L_X2Y121_SLICE_X0Y121_CO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D = CLBLL_L_X2Y121_SLICE_X0Y121_DO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_AMUX = CLBLL_L_X2Y121_SLICE_X0Y121_A5Q;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_BMUX = CLBLL_L_X2Y121_SLICE_X0Y121_BO5;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A = CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B = CLBLL_L_X2Y121_SLICE_X1Y121_BO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C = CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D = CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_AMUX = CLBLL_L_X2Y121_SLICE_X1Y121_AO5;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_BMUX = CLBLL_L_X2Y121_SLICE_X1Y121_B5Q;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_CMUX = CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A = CLBLL_L_X2Y122_SLICE_X0Y122_AO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B = CLBLL_L_X2Y122_SLICE_X0Y122_BO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C = CLBLL_L_X2Y122_SLICE_X0Y122_CO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D = CLBLL_L_X2Y122_SLICE_X0Y122_DO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A = CLBLL_L_X2Y122_SLICE_X1Y122_AO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B = CLBLL_L_X2Y122_SLICE_X1Y122_BO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C = CLBLL_L_X2Y122_SLICE_X1Y122_CO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D = CLBLL_L_X2Y122_SLICE_X1Y122_DO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_AMUX = CLBLL_L_X2Y122_SLICE_X1Y122_A5Q;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A = CLBLL_L_X2Y125_SLICE_X0Y125_AO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B = CLBLL_L_X2Y125_SLICE_X0Y125_BO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C = CLBLL_L_X2Y125_SLICE_X0Y125_CO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D = CLBLL_L_X2Y125_SLICE_X0Y125_DO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A = CLBLL_L_X2Y125_SLICE_X1Y125_AO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B = CLBLL_L_X2Y125_SLICE_X1Y125_BO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C = CLBLL_L_X2Y125_SLICE_X1Y125_CO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D = CLBLL_L_X2Y125_SLICE_X1Y125_DO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_CMUX = CLBLL_L_X2Y125_SLICE_X1Y125_CO5;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_A = CLBLL_L_X2Y126_SLICE_X0Y126_AO6;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_B = CLBLL_L_X2Y126_SLICE_X0Y126_BO6;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_C = CLBLL_L_X2Y126_SLICE_X0Y126_CO6;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_D = CLBLL_L_X2Y126_SLICE_X0Y126_DO6;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_AMUX = CLBLL_L_X2Y126_SLICE_X0Y126_AO5;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_A = CLBLL_L_X2Y126_SLICE_X1Y126_AO6;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_B = CLBLL_L_X2Y126_SLICE_X1Y126_BO6;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_C = CLBLL_L_X2Y126_SLICE_X1Y126_CO6;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_D = CLBLL_L_X2Y126_SLICE_X1Y126_DO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A = CLBLL_L_X2Y127_SLICE_X0Y127_AO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B = CLBLL_L_X2Y127_SLICE_X0Y127_BO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C = CLBLL_L_X2Y127_SLICE_X0Y127_CO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D = CLBLL_L_X2Y127_SLICE_X0Y127_DO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_BMUX = CLBLL_L_X2Y127_SLICE_X0Y127_BO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A = CLBLL_L_X2Y127_SLICE_X1Y127_AO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B = CLBLL_L_X2Y127_SLICE_X1Y127_BO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C = CLBLL_L_X2Y127_SLICE_X1Y127_CO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D = CLBLL_L_X2Y127_SLICE_X1Y127_DO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_A = CLBLL_L_X2Y128_SLICE_X0Y128_AO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_B = CLBLL_L_X2Y128_SLICE_X0Y128_BO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_C = CLBLL_L_X2Y128_SLICE_X0Y128_CO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_D = CLBLL_L_X2Y128_SLICE_X0Y128_DO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_AMUX = CLBLL_L_X2Y128_SLICE_X0Y128_AO5;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_BMUX = CLBLL_L_X2Y128_SLICE_X0Y128_BO5;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_CMUX = CLBLL_L_X2Y128_SLICE_X0Y128_CO6;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_A = CLBLL_L_X2Y128_SLICE_X1Y128_AO6;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_B = CLBLL_L_X2Y128_SLICE_X1Y128_BO6;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_C = CLBLL_L_X2Y128_SLICE_X1Y128_CO6;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_D = CLBLL_L_X2Y128_SLICE_X1Y128_DO6;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_AMUX = CLBLL_L_X2Y128_SLICE_X1Y128_AO5;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_BMUX = CLBLL_L_X2Y128_SLICE_X1Y128_BO5;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A = CLBLL_L_X2Y129_SLICE_X0Y129_AO6;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B = CLBLL_L_X2Y129_SLICE_X0Y129_BO6;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C = CLBLL_L_X2Y129_SLICE_X0Y129_CO6;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D = CLBLL_L_X2Y129_SLICE_X0Y129_DO6;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_AMUX = CLBLL_L_X2Y129_SLICE_X0Y129_AO5;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_CMUX = CLBLL_L_X2Y129_SLICE_X0Y129_CO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A = CLBLL_L_X2Y129_SLICE_X1Y129_AO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B = CLBLL_L_X2Y129_SLICE_X1Y129_BO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C = CLBLL_L_X2Y129_SLICE_X1Y129_CO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D = CLBLL_L_X2Y129_SLICE_X1Y129_DO6;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_A = CLBLL_L_X2Y130_SLICE_X0Y130_AO6;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_B = CLBLL_L_X2Y130_SLICE_X0Y130_BO6;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_C = CLBLL_L_X2Y130_SLICE_X0Y130_CO6;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_D = CLBLL_L_X2Y130_SLICE_X0Y130_DO6;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_AMUX = CLBLL_L_X2Y130_SLICE_X0Y130_AO5;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_BMUX = CLBLL_L_X2Y130_SLICE_X0Y130_BO5;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_CMUX = CLBLL_L_X2Y130_SLICE_X0Y130_CO5;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_DMUX = CLBLL_L_X2Y130_SLICE_X0Y130_DO6;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_A = CLBLL_L_X2Y130_SLICE_X1Y130_AO6;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_B = CLBLL_L_X2Y130_SLICE_X1Y130_BO6;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_C = CLBLL_L_X2Y130_SLICE_X1Y130_CO6;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_D = CLBLL_L_X2Y130_SLICE_X1Y130_DO6;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_AMUX = CLBLL_L_X2Y130_SLICE_X1Y130_AO5;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_BMUX = CLBLL_L_X2Y130_SLICE_X1Y130_BO5;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A = CLBLL_L_X2Y131_SLICE_X0Y131_AO6;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B = CLBLL_L_X2Y131_SLICE_X0Y131_BO6;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C = CLBLL_L_X2Y131_SLICE_X0Y131_CO6;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D = CLBLL_L_X2Y131_SLICE_X0Y131_DO6;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A = CLBLL_L_X2Y131_SLICE_X1Y131_AO6;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B = CLBLL_L_X2Y131_SLICE_X1Y131_BO6;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C = CLBLL_L_X2Y131_SLICE_X1Y131_CO6;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D = CLBLL_L_X2Y131_SLICE_X1Y131_DO6;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_A = CLBLL_L_X2Y132_SLICE_X0Y132_AO6;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_B = CLBLL_L_X2Y132_SLICE_X0Y132_BO6;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_C = CLBLL_L_X2Y132_SLICE_X0Y132_CO6;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_D = CLBLL_L_X2Y132_SLICE_X0Y132_DO6;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_A = CLBLL_L_X2Y132_SLICE_X1Y132_AO6;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_B = CLBLL_L_X2Y132_SLICE_X1Y132_BO6;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_C = CLBLL_L_X2Y132_SLICE_X1Y132_CO6;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_D = CLBLL_L_X2Y132_SLICE_X1Y132_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A = CLBLL_L_X4Y117_SLICE_X4Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B = CLBLL_L_X4Y117_SLICE_X4Y117_BO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C = CLBLL_L_X4Y117_SLICE_X4Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D = CLBLL_L_X4Y117_SLICE_X4Y117_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_AMUX = CLBLL_L_X4Y117_SLICE_X4Y117_AO5;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A = CLBLL_L_X4Y117_SLICE_X5Y117_AO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B = CLBLL_L_X4Y117_SLICE_X5Y117_BO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C = CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D = CLBLL_L_X4Y117_SLICE_X5Y117_DO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_CMUX = CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A = CLBLL_L_X4Y118_SLICE_X4Y118_AO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B = CLBLL_L_X4Y118_SLICE_X4Y118_BO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C = CLBLL_L_X4Y118_SLICE_X4Y118_CO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D = CLBLL_L_X4Y118_SLICE_X4Y118_DO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A = CLBLL_L_X4Y118_SLICE_X5Y118_AO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B = CLBLL_L_X4Y118_SLICE_X5Y118_BO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C = CLBLL_L_X4Y118_SLICE_X5Y118_CO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D = CLBLL_L_X4Y118_SLICE_X5Y118_DO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_CMUX = CLBLL_L_X4Y118_SLICE_X5Y118_C5Q;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A = CLBLL_L_X4Y119_SLICE_X4Y119_AO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B = CLBLL_L_X4Y119_SLICE_X4Y119_BO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C = CLBLL_L_X4Y119_SLICE_X4Y119_CO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D = CLBLL_L_X4Y119_SLICE_X4Y119_DO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A = CLBLL_L_X4Y119_SLICE_X5Y119_AO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B = CLBLL_L_X4Y119_SLICE_X5Y119_BO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C = CLBLL_L_X4Y119_SLICE_X5Y119_CO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D = CLBLL_L_X4Y119_SLICE_X5Y119_DO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_DMUX = CLBLL_L_X4Y119_SLICE_X5Y119_DO5;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A = CLBLL_L_X4Y120_SLICE_X4Y120_AO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B = CLBLL_L_X4Y120_SLICE_X4Y120_BO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C = CLBLL_L_X4Y120_SLICE_X4Y120_CO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D = CLBLL_L_X4Y120_SLICE_X4Y120_DO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_AMUX = CLBLL_L_X4Y120_SLICE_X4Y120_A5Q;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_CMUX = CLBLL_L_X4Y120_SLICE_X4Y120_C5Q;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A = CLBLL_L_X4Y120_SLICE_X5Y120_AO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B = CLBLL_L_X4Y120_SLICE_X5Y120_BO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C = CLBLL_L_X4Y120_SLICE_X5Y120_CO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D = CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_AMUX = CLBLL_L_X4Y120_SLICE_X5Y120_A5Q;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A = CLBLL_L_X4Y121_SLICE_X4Y121_AO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B = CLBLL_L_X4Y121_SLICE_X4Y121_BO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C = CLBLL_L_X4Y121_SLICE_X4Y121_CO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D = CLBLL_L_X4Y121_SLICE_X4Y121_DO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A = CLBLL_L_X4Y121_SLICE_X5Y121_AO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B = CLBLL_L_X4Y121_SLICE_X5Y121_BO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C = CLBLL_L_X4Y121_SLICE_X5Y121_CO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D = CLBLL_L_X4Y121_SLICE_X5Y121_DO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A = CLBLL_L_X4Y122_SLICE_X4Y122_AO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B = CLBLL_L_X4Y122_SLICE_X4Y122_BO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C = CLBLL_L_X4Y122_SLICE_X4Y122_CO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D = CLBLL_L_X4Y122_SLICE_X4Y122_DO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_AMUX = CLBLL_L_X4Y122_SLICE_X4Y122_A5Q;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_CMUX = CLBLL_L_X4Y122_SLICE_X4Y122_CO5;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A = CLBLL_L_X4Y122_SLICE_X5Y122_AO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B = CLBLL_L_X4Y122_SLICE_X5Y122_BO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C = CLBLL_L_X4Y122_SLICE_X5Y122_CO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D = CLBLL_L_X4Y122_SLICE_X5Y122_DO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_CMUX = CLBLL_L_X4Y122_SLICE_X5Y122_C5Q;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A = CLBLL_L_X4Y123_SLICE_X4Y123_AO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B = CLBLL_L_X4Y123_SLICE_X4Y123_BO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C = CLBLL_L_X4Y123_SLICE_X4Y123_CO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D = CLBLL_L_X4Y123_SLICE_X4Y123_DO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A = CLBLL_L_X4Y123_SLICE_X5Y123_AO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B = CLBLL_L_X4Y123_SLICE_X5Y123_BO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C = CLBLL_L_X4Y123_SLICE_X5Y123_CO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D = CLBLL_L_X4Y123_SLICE_X5Y123_DO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_BMUX = CLBLL_L_X4Y123_SLICE_X5Y123_B5Q;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_CMUX = CLBLL_L_X4Y123_SLICE_X5Y123_CO5;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A = CLBLL_L_X4Y124_SLICE_X4Y124_AO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B = CLBLL_L_X4Y124_SLICE_X4Y124_BO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C = CLBLL_L_X4Y124_SLICE_X4Y124_CO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D = CLBLL_L_X4Y124_SLICE_X4Y124_DO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_AMUX = CLBLL_L_X4Y124_SLICE_X4Y124_A5Q;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A = CLBLL_L_X4Y124_SLICE_X5Y124_AO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B = CLBLL_L_X4Y124_SLICE_X5Y124_BO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C = CLBLL_L_X4Y124_SLICE_X5Y124_CO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D = CLBLL_L_X4Y124_SLICE_X5Y124_DO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A = CLBLL_L_X4Y125_SLICE_X4Y125_AO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B = CLBLL_L_X4Y125_SLICE_X4Y125_BO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C = CLBLL_L_X4Y125_SLICE_X4Y125_CO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D = CLBLL_L_X4Y125_SLICE_X4Y125_DO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_CMUX = CLBLL_L_X4Y125_SLICE_X4Y125_C5Q;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A = CLBLL_L_X4Y125_SLICE_X5Y125_AO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B = CLBLL_L_X4Y125_SLICE_X5Y125_BO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C = CLBLL_L_X4Y125_SLICE_X5Y125_CO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D = CLBLL_L_X4Y125_SLICE_X5Y125_DO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A = CLBLL_L_X4Y126_SLICE_X4Y126_AO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B = CLBLL_L_X4Y126_SLICE_X4Y126_BO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C = CLBLL_L_X4Y126_SLICE_X4Y126_CO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D = CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_BMUX = CLBLL_L_X4Y126_SLICE_X4Y126_BO5;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_CMUX = CLBLL_L_X4Y126_SLICE_X4Y126_CO5;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A = CLBLL_L_X4Y126_SLICE_X5Y126_AO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B = CLBLL_L_X4Y126_SLICE_X5Y126_BO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C = CLBLL_L_X4Y126_SLICE_X5Y126_CO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D = CLBLL_L_X4Y126_SLICE_X5Y126_DO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A = CLBLL_L_X4Y127_SLICE_X4Y127_AO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B = CLBLL_L_X4Y127_SLICE_X4Y127_BO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C = CLBLL_L_X4Y127_SLICE_X4Y127_CO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D = CLBLL_L_X4Y127_SLICE_X4Y127_DO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_AMUX = CLBLL_L_X4Y127_SLICE_X4Y127_AO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_CMUX = CLBLL_L_X4Y127_SLICE_X4Y127_CO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A = CLBLL_L_X4Y127_SLICE_X5Y127_AO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B = CLBLL_L_X4Y127_SLICE_X5Y127_BO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C = CLBLL_L_X4Y127_SLICE_X5Y127_CO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D = CLBLL_L_X4Y127_SLICE_X5Y127_DO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_CMUX = CLBLL_L_X4Y127_SLICE_X5Y127_CO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A = CLBLL_L_X4Y128_SLICE_X4Y128_AO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B = CLBLL_L_X4Y128_SLICE_X4Y128_BO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C = CLBLL_L_X4Y128_SLICE_X4Y128_CO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D = CLBLL_L_X4Y128_SLICE_X4Y128_DO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A = CLBLL_L_X4Y128_SLICE_X5Y128_AO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B = CLBLL_L_X4Y128_SLICE_X5Y128_BO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C = CLBLL_L_X4Y128_SLICE_X5Y128_CO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D = CLBLL_L_X4Y128_SLICE_X5Y128_DO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_CMUX = CLBLL_L_X4Y128_SLICE_X5Y128_CO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A = CLBLL_L_X4Y129_SLICE_X4Y129_AO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B = CLBLL_L_X4Y129_SLICE_X4Y129_BO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C = CLBLL_L_X4Y129_SLICE_X4Y129_CO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D = CLBLL_L_X4Y129_SLICE_X4Y129_DO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_BMUX = CLBLL_L_X4Y129_SLICE_X4Y129_BO5;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A = CLBLL_L_X4Y129_SLICE_X5Y129_AO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B = CLBLL_L_X4Y129_SLICE_X5Y129_BO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C = CLBLL_L_X4Y129_SLICE_X5Y129_CO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D = CLBLL_L_X4Y129_SLICE_X5Y129_DO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A = CLBLL_L_X4Y130_SLICE_X4Y130_AO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B = CLBLL_L_X4Y130_SLICE_X4Y130_BO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C = CLBLL_L_X4Y130_SLICE_X4Y130_CO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D = CLBLL_L_X4Y130_SLICE_X4Y130_DO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_AMUX = CLBLL_L_X4Y130_SLICE_X4Y130_AO5;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A = CLBLL_L_X4Y130_SLICE_X5Y130_AO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B = CLBLL_L_X4Y130_SLICE_X5Y130_BO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C = CLBLL_L_X4Y130_SLICE_X5Y130_CO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D = CLBLL_L_X4Y130_SLICE_X5Y130_DO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A = CLBLL_L_X4Y131_SLICE_X4Y131_AO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C = CLBLL_L_X4Y131_SLICE_X4Y131_CO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D = CLBLL_L_X4Y131_SLICE_X4Y131_DO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A = CLBLL_L_X4Y131_SLICE_X5Y131_AO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B = CLBLL_L_X4Y131_SLICE_X5Y131_BO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C = CLBLL_L_X4Y131_SLICE_X5Y131_CO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D = CLBLL_L_X4Y131_SLICE_X5Y131_DO6;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_A = CLBLL_L_X36Y124_SLICE_X54Y124_AO6;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_B = CLBLL_L_X36Y124_SLICE_X54Y124_BO6;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_C = CLBLL_L_X36Y124_SLICE_X54Y124_CO6;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_D = CLBLL_L_X36Y124_SLICE_X54Y124_DO6;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_A = CLBLL_L_X36Y124_SLICE_X55Y124_AO6;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_B = CLBLL_L_X36Y124_SLICE_X55Y124_BO6;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_C = CLBLL_L_X36Y124_SLICE_X55Y124_CO6;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_D = CLBLL_L_X36Y124_SLICE_X55Y124_DO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B = CLBLL_L_X52Y126_SLICE_X78Y126_BO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C = CLBLL_L_X52Y126_SLICE_X78Y126_CO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D = CLBLL_L_X52Y126_SLICE_X78Y126_DO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A = CLBLL_L_X52Y126_SLICE_X79Y126_AO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B = CLBLL_L_X52Y126_SLICE_X79Y126_BO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C = CLBLL_L_X52Y126_SLICE_X79Y126_CO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D = CLBLL_L_X52Y126_SLICE_X79Y126_DO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A = CLBLM_L_X8Y116_SLICE_X10Y116_AO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B = CLBLM_L_X8Y116_SLICE_X10Y116_BO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C = CLBLM_L_X8Y116_SLICE_X10Y116_CO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D = CLBLM_L_X8Y116_SLICE_X10Y116_DO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_AMUX = CLBLM_L_X8Y116_SLICE_X10Y116_AO5;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_CMUX = CLBLM_L_X8Y116_SLICE_X10Y116_CO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A = CLBLM_L_X8Y116_SLICE_X11Y116_AO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C = CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D = CLBLM_L_X8Y116_SLICE_X11Y116_DO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A = CLBLM_L_X8Y117_SLICE_X10Y117_AO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B = CLBLM_L_X8Y117_SLICE_X10Y117_BO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C = CLBLM_L_X8Y117_SLICE_X10Y117_CO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D = CLBLM_L_X8Y117_SLICE_X10Y117_DO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_CMUX = CLBLM_L_X8Y117_SLICE_X10Y117_CO5;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_DMUX = CLBLM_L_X8Y117_SLICE_X10Y117_DO5;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A = CLBLM_L_X8Y117_SLICE_X11Y117_AO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B = CLBLM_L_X8Y117_SLICE_X11Y117_BO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D = CLBLM_L_X8Y117_SLICE_X11Y117_DO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_AMUX = CLBLM_L_X8Y117_SLICE_X11Y117_AO5;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A = CLBLM_L_X8Y118_SLICE_X10Y118_AO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B = CLBLM_L_X8Y118_SLICE_X10Y118_BO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C = CLBLM_L_X8Y118_SLICE_X10Y118_CO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D = CLBLM_L_X8Y118_SLICE_X10Y118_DO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_AMUX = CLBLM_L_X8Y118_SLICE_X10Y118_AO5;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A = CLBLM_L_X8Y118_SLICE_X11Y118_AO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B = CLBLM_L_X8Y118_SLICE_X11Y118_BO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C = CLBLM_L_X8Y118_SLICE_X11Y118_CO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D = CLBLM_L_X8Y118_SLICE_X11Y118_DO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_CMUX = CLBLM_L_X8Y118_SLICE_X11Y118_CO5;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A = CLBLM_L_X8Y119_SLICE_X10Y119_AO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B = CLBLM_L_X8Y119_SLICE_X10Y119_BO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C = CLBLM_L_X8Y119_SLICE_X10Y119_CO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D = CLBLM_L_X8Y119_SLICE_X10Y119_DO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A = CLBLM_L_X8Y119_SLICE_X11Y119_AO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B = CLBLM_L_X8Y119_SLICE_X11Y119_BO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C = CLBLM_L_X8Y119_SLICE_X11Y119_CO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D = CLBLM_L_X8Y119_SLICE_X11Y119_DO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A = CLBLM_L_X8Y120_SLICE_X10Y120_AO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B = CLBLM_L_X8Y120_SLICE_X10Y120_BO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C = CLBLM_L_X8Y120_SLICE_X10Y120_CO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D = CLBLM_L_X8Y120_SLICE_X10Y120_DO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A = CLBLM_L_X8Y120_SLICE_X11Y120_AO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B = CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C = CLBLM_L_X8Y120_SLICE_X11Y120_CO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D = CLBLM_L_X8Y120_SLICE_X11Y120_DO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A = CLBLM_L_X8Y121_SLICE_X10Y121_AO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B = CLBLM_L_X8Y121_SLICE_X10Y121_BO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C = CLBLM_L_X8Y121_SLICE_X10Y121_CO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D = CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_AMUX = CLBLM_L_X8Y121_SLICE_X10Y121_AO5;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_DMUX = CLBLM_L_X8Y121_SLICE_X10Y121_DO5;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A = CLBLM_L_X8Y121_SLICE_X11Y121_AO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B = CLBLM_L_X8Y121_SLICE_X11Y121_BO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C = CLBLM_L_X8Y121_SLICE_X11Y121_CO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D = CLBLM_L_X8Y121_SLICE_X11Y121_DO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_DMUX = CLBLM_L_X8Y121_SLICE_X11Y121_DO5;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A = CLBLM_L_X8Y122_SLICE_X10Y122_AO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B = CLBLM_L_X8Y122_SLICE_X10Y122_BO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C = CLBLM_L_X8Y122_SLICE_X10Y122_CO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D = CLBLM_L_X8Y122_SLICE_X10Y122_DO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_AMUX = CLBLM_L_X8Y122_SLICE_X10Y122_A5Q;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A = CLBLM_L_X8Y122_SLICE_X11Y122_AO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B = CLBLM_L_X8Y122_SLICE_X11Y122_BO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C = CLBLM_L_X8Y122_SLICE_X11Y122_CO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D = CLBLM_L_X8Y122_SLICE_X11Y122_DO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_AMUX = CLBLM_L_X8Y122_SLICE_X11Y122_A5Q;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A = CLBLM_L_X8Y123_SLICE_X10Y123_AO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B = CLBLM_L_X8Y123_SLICE_X10Y123_BO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C = CLBLM_L_X8Y123_SLICE_X10Y123_CO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D = CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_CMUX = CLBLM_L_X8Y123_SLICE_X10Y123_C5Q;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A = CLBLM_L_X8Y123_SLICE_X11Y123_AO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B = CLBLM_L_X8Y123_SLICE_X11Y123_BO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C = CLBLM_L_X8Y123_SLICE_X11Y123_CO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D = CLBLM_L_X8Y123_SLICE_X11Y123_DO6;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_CMUX = CLBLM_L_X8Y123_SLICE_X11Y123_C5Q;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_DMUX = CLBLM_L_X8Y123_SLICE_X11Y123_DO5;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A = CLBLM_L_X8Y124_SLICE_X10Y124_AO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B = CLBLM_L_X8Y124_SLICE_X10Y124_BO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C = CLBLM_L_X8Y124_SLICE_X10Y124_CO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D = CLBLM_L_X8Y124_SLICE_X10Y124_DO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_BMUX = CLBLM_L_X8Y124_SLICE_X10Y124_B5Q;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A = CLBLM_L_X8Y124_SLICE_X11Y124_AO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B = CLBLM_L_X8Y124_SLICE_X11Y124_BO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C = CLBLM_L_X8Y124_SLICE_X11Y124_CO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D = CLBLM_L_X8Y124_SLICE_X11Y124_DO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_CMUX = CLBLM_L_X8Y124_SLICE_X11Y124_CO5;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A = CLBLM_L_X8Y125_SLICE_X10Y125_AO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B = CLBLM_L_X8Y125_SLICE_X10Y125_BO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C = CLBLM_L_X8Y125_SLICE_X10Y125_CO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D = CLBLM_L_X8Y125_SLICE_X10Y125_DO6;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_BMUX = CLBLM_L_X8Y125_SLICE_X10Y125_BO5;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A = CLBLM_L_X8Y125_SLICE_X11Y125_AO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B = CLBLM_L_X8Y125_SLICE_X11Y125_BO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C = CLBLM_L_X8Y125_SLICE_X11Y125_CO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D = CLBLM_L_X8Y125_SLICE_X11Y125_DO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A = CLBLM_L_X8Y126_SLICE_X10Y126_AO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B = CLBLM_L_X8Y126_SLICE_X10Y126_BO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C = CLBLM_L_X8Y126_SLICE_X10Y126_CO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D = CLBLM_L_X8Y126_SLICE_X10Y126_DO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_AMUX = CLBLM_L_X8Y126_SLICE_X10Y126_AO5;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A = CLBLM_L_X8Y126_SLICE_X11Y126_AO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B = CLBLM_L_X8Y126_SLICE_X11Y126_BO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C = CLBLM_L_X8Y126_SLICE_X11Y126_CO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D = CLBLM_L_X8Y126_SLICE_X11Y126_DO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_BMUX = CLBLM_L_X8Y126_SLICE_X11Y126_B5Q;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A = CLBLM_L_X8Y127_SLICE_X10Y127_AO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B = CLBLM_L_X8Y127_SLICE_X10Y127_BO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C = CLBLM_L_X8Y127_SLICE_X10Y127_CO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D = CLBLM_L_X8Y127_SLICE_X10Y127_DO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_DMUX = CLBLM_L_X8Y127_SLICE_X10Y127_DO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A = CLBLM_L_X8Y127_SLICE_X11Y127_AO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B = CLBLM_L_X8Y127_SLICE_X11Y127_BO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C = CLBLM_L_X8Y127_SLICE_X11Y127_CO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D = CLBLM_L_X8Y127_SLICE_X11Y127_DO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A = CLBLM_L_X8Y128_SLICE_X10Y128_AO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B = CLBLM_L_X8Y128_SLICE_X10Y128_BO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C = CLBLM_L_X8Y128_SLICE_X10Y128_CO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D = CLBLM_L_X8Y128_SLICE_X10Y128_DO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A = CLBLM_L_X8Y128_SLICE_X11Y128_AO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B = CLBLM_L_X8Y128_SLICE_X11Y128_BO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C = CLBLM_L_X8Y128_SLICE_X11Y128_CO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D = CLBLM_L_X8Y128_SLICE_X11Y128_DO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A = CLBLM_L_X8Y129_SLICE_X10Y129_AO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B = CLBLM_L_X8Y129_SLICE_X10Y129_BO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C = CLBLM_L_X8Y129_SLICE_X10Y129_CO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D = CLBLM_L_X8Y129_SLICE_X10Y129_DO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_AMUX = CLBLM_L_X8Y129_SLICE_X10Y129_AO5;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_BMUX = CLBLM_L_X8Y129_SLICE_X10Y129_BO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A = CLBLM_L_X8Y129_SLICE_X11Y129_AO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B = CLBLM_L_X8Y129_SLICE_X11Y129_BO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C = CLBLM_L_X8Y129_SLICE_X11Y129_CO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D = CLBLM_L_X8Y129_SLICE_X11Y129_DO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_BMUX = CLBLM_L_X8Y129_SLICE_X11Y129_B5Q;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A = CLBLM_L_X8Y130_SLICE_X10Y130_AO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B = CLBLM_L_X8Y130_SLICE_X10Y130_BO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C = CLBLM_L_X8Y130_SLICE_X10Y130_CO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D = CLBLM_L_X8Y130_SLICE_X10Y130_DO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A = CLBLM_L_X8Y130_SLICE_X11Y130_AO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B = CLBLM_L_X8Y130_SLICE_X11Y130_BO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C = CLBLM_L_X8Y130_SLICE_X11Y130_CO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D = CLBLM_L_X8Y130_SLICE_X11Y130_DO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_AMUX = CLBLM_L_X8Y130_SLICE_X11Y130_AO5;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A = CLBLM_L_X8Y131_SLICE_X10Y131_AO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B = CLBLM_L_X8Y131_SLICE_X10Y131_BO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C = CLBLM_L_X8Y131_SLICE_X10Y131_CO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D = CLBLM_L_X8Y131_SLICE_X10Y131_DO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_AMUX = CLBLM_L_X8Y131_SLICE_X10Y131_AO5;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_BMUX = CLBLM_L_X8Y131_SLICE_X10Y131_BO5;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A = CLBLM_L_X8Y131_SLICE_X11Y131_AO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B = CLBLM_L_X8Y131_SLICE_X11Y131_BO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C = CLBLM_L_X8Y131_SLICE_X11Y131_CO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D = CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A = CLBLM_L_X10Y117_SLICE_X12Y117_AO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B = CLBLM_L_X10Y117_SLICE_X12Y117_BO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C = CLBLM_L_X10Y117_SLICE_X12Y117_CO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D = CLBLM_L_X10Y117_SLICE_X12Y117_DO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A = CLBLM_L_X10Y117_SLICE_X13Y117_AO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B = CLBLM_L_X10Y117_SLICE_X13Y117_BO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C = CLBLM_L_X10Y117_SLICE_X13Y117_CO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D = CLBLM_L_X10Y117_SLICE_X13Y117_DO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A = CLBLM_L_X10Y118_SLICE_X12Y118_AO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B = CLBLM_L_X10Y118_SLICE_X12Y118_BO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C = CLBLM_L_X10Y118_SLICE_X12Y118_CO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D = CLBLM_L_X10Y118_SLICE_X12Y118_DO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A = CLBLM_L_X10Y118_SLICE_X13Y118_AO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B = CLBLM_L_X10Y118_SLICE_X13Y118_BO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C = CLBLM_L_X10Y118_SLICE_X13Y118_CO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D = CLBLM_L_X10Y118_SLICE_X13Y118_DO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A = CLBLM_L_X10Y119_SLICE_X12Y119_AO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B = CLBLM_L_X10Y119_SLICE_X12Y119_BO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C = CLBLM_L_X10Y119_SLICE_X12Y119_CO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D = CLBLM_L_X10Y119_SLICE_X12Y119_DO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A = CLBLM_L_X10Y119_SLICE_X13Y119_AO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B = CLBLM_L_X10Y119_SLICE_X13Y119_BO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C = CLBLM_L_X10Y119_SLICE_X13Y119_CO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D = CLBLM_L_X10Y119_SLICE_X13Y119_DO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A = CLBLM_L_X10Y120_SLICE_X12Y120_AO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B = CLBLM_L_X10Y120_SLICE_X12Y120_BO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C = CLBLM_L_X10Y120_SLICE_X12Y120_CO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D = CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A = CLBLM_L_X10Y120_SLICE_X13Y120_AO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B = CLBLM_L_X10Y120_SLICE_X13Y120_BO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C = CLBLM_L_X10Y120_SLICE_X13Y120_CO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D = CLBLM_L_X10Y120_SLICE_X13Y120_DO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_AMUX = CLBLM_L_X10Y120_SLICE_X13Y120_A5Q;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_BMUX = CLBLM_L_X10Y120_SLICE_X13Y120_BO5;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A = CLBLM_L_X10Y121_SLICE_X12Y121_AO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B = CLBLM_L_X10Y121_SLICE_X12Y121_BO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C = CLBLM_L_X10Y121_SLICE_X12Y121_CO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D = CLBLM_L_X10Y121_SLICE_X12Y121_DO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_CMUX = CLBLM_L_X10Y121_SLICE_X12Y121_C5Q;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A = CLBLM_L_X10Y121_SLICE_X13Y121_AO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B = CLBLM_L_X10Y121_SLICE_X13Y121_BO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C = CLBLM_L_X10Y121_SLICE_X13Y121_CO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D = CLBLM_L_X10Y121_SLICE_X13Y121_DO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_BMUX = CLBLM_L_X10Y121_SLICE_X13Y121_B5Q;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A = CLBLM_L_X10Y122_SLICE_X12Y122_AO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B = CLBLM_L_X10Y122_SLICE_X12Y122_BO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C = CLBLM_L_X10Y122_SLICE_X12Y122_CO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D = CLBLM_L_X10Y122_SLICE_X12Y122_DO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A = CLBLM_L_X10Y122_SLICE_X13Y122_AO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B = CLBLM_L_X10Y122_SLICE_X13Y122_BO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C = CLBLM_L_X10Y122_SLICE_X13Y122_CO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D = CLBLM_L_X10Y122_SLICE_X13Y122_DO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_BMUX = CLBLM_L_X10Y122_SLICE_X13Y122_BO5;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_CMUX = CLBLM_L_X10Y122_SLICE_X13Y122_C5Q;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A = CLBLM_L_X10Y123_SLICE_X12Y123_AO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B = CLBLM_L_X10Y123_SLICE_X12Y123_BO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C = CLBLM_L_X10Y123_SLICE_X12Y123_CO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D = CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_DMUX = CLBLM_L_X10Y123_SLICE_X12Y123_DO5;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A = CLBLM_L_X10Y123_SLICE_X13Y123_AO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B = CLBLM_L_X10Y123_SLICE_X13Y123_BO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C = CLBLM_L_X10Y123_SLICE_X13Y123_CO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D = CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_DMUX = CLBLM_L_X10Y123_SLICE_X13Y123_DO5;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A = CLBLM_L_X10Y124_SLICE_X12Y124_AO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B = CLBLM_L_X10Y124_SLICE_X12Y124_BO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C = CLBLM_L_X10Y124_SLICE_X12Y124_CO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D = CLBLM_L_X10Y124_SLICE_X12Y124_DO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_AMUX = CLBLM_L_X10Y124_SLICE_X12Y124_AO5;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_BMUX = CLBLM_L_X10Y124_SLICE_X12Y124_BO5;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_CMUX = CLBLM_L_X10Y124_SLICE_X12Y124_CO5;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A = CLBLM_L_X10Y124_SLICE_X13Y124_AO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B = CLBLM_L_X10Y124_SLICE_X13Y124_BO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C = CLBLM_L_X10Y124_SLICE_X13Y124_CO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D = CLBLM_L_X10Y124_SLICE_X13Y124_DO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_AMUX = CLBLM_L_X10Y124_SLICE_X13Y124_A5Q;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_BMUX = CLBLM_L_X10Y124_SLICE_X13Y124_B5Q;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_CMUX = CLBLM_L_X10Y124_SLICE_X13Y124_C5Q;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_DMUX = CLBLM_L_X10Y124_SLICE_X13Y124_D5Q;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A = CLBLM_L_X10Y125_SLICE_X12Y125_AO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B = CLBLM_L_X10Y125_SLICE_X12Y125_BO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C = CLBLM_L_X10Y125_SLICE_X12Y125_CO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D = CLBLM_L_X10Y125_SLICE_X12Y125_DO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A = CLBLM_L_X10Y125_SLICE_X13Y125_AO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B = CLBLM_L_X10Y125_SLICE_X13Y125_BO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C = CLBLM_L_X10Y125_SLICE_X13Y125_CO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D = CLBLM_L_X10Y125_SLICE_X13Y125_DO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_DMUX = CLBLM_L_X10Y125_SLICE_X13Y125_DO5;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A = CLBLM_L_X10Y126_SLICE_X12Y126_AO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B = CLBLM_L_X10Y126_SLICE_X12Y126_BO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C = CLBLM_L_X10Y126_SLICE_X12Y126_CO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D = CLBLM_L_X10Y126_SLICE_X12Y126_DO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_AMUX = CLBLM_L_X10Y126_SLICE_X12Y126_A5Q;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_BMUX = CLBLM_L_X10Y126_SLICE_X12Y126_BO5;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_DMUX = CLBLM_L_X10Y126_SLICE_X12Y126_DO5;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A = CLBLM_L_X10Y126_SLICE_X13Y126_AO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B = CLBLM_L_X10Y126_SLICE_X13Y126_BO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C = CLBLM_L_X10Y126_SLICE_X13Y126_CO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D = CLBLM_L_X10Y126_SLICE_X13Y126_DO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A = CLBLM_L_X10Y127_SLICE_X12Y127_AO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B = CLBLM_L_X10Y127_SLICE_X12Y127_BO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C = CLBLM_L_X10Y127_SLICE_X12Y127_CO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D = CLBLM_L_X10Y127_SLICE_X12Y127_DO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A = CLBLM_L_X10Y127_SLICE_X13Y127_AO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B = CLBLM_L_X10Y127_SLICE_X13Y127_BO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C = CLBLM_L_X10Y127_SLICE_X13Y127_CO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D = CLBLM_L_X10Y127_SLICE_X13Y127_DO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A = CLBLM_L_X10Y128_SLICE_X12Y128_AO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B = CLBLM_L_X10Y128_SLICE_X12Y128_BO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C = CLBLM_L_X10Y128_SLICE_X12Y128_CO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D = CLBLM_L_X10Y128_SLICE_X12Y128_DO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A = CLBLM_L_X10Y128_SLICE_X13Y128_AO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B = CLBLM_L_X10Y128_SLICE_X13Y128_BO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C = CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D = CLBLM_L_X10Y128_SLICE_X13Y128_DO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_CMUX = CLBLM_L_X10Y128_SLICE_X13Y128_CO5;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A = CLBLM_L_X10Y129_SLICE_X12Y129_AO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B = CLBLM_L_X10Y129_SLICE_X12Y129_BO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C = CLBLM_L_X10Y129_SLICE_X12Y129_CO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D = CLBLM_L_X10Y129_SLICE_X12Y129_DO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_AMUX = CLBLM_L_X10Y129_SLICE_X12Y129_A5Q;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A = CLBLM_L_X10Y129_SLICE_X13Y129_AO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B = CLBLM_L_X10Y129_SLICE_X13Y129_BO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C = CLBLM_L_X10Y129_SLICE_X13Y129_CO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D = CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_BMUX = CLBLM_L_X10Y129_SLICE_X13Y129_BO5;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A = CLBLM_L_X10Y130_SLICE_X12Y130_AO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B = CLBLM_L_X10Y130_SLICE_X12Y130_BO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C = CLBLM_L_X10Y130_SLICE_X12Y130_CO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D = CLBLM_L_X10Y130_SLICE_X12Y130_DO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A = CLBLM_L_X10Y130_SLICE_X13Y130_AO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B = CLBLM_L_X10Y130_SLICE_X13Y130_BO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C = CLBLM_L_X10Y130_SLICE_X13Y130_CO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D = CLBLM_L_X10Y130_SLICE_X13Y130_DO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A = CLBLM_L_X10Y135_SLICE_X12Y135_AO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B = CLBLM_L_X10Y135_SLICE_X12Y135_BO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C = CLBLM_L_X10Y135_SLICE_X12Y135_CO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A = CLBLM_L_X10Y135_SLICE_X13Y135_AO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B = CLBLM_L_X10Y135_SLICE_X13Y135_BO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C = CLBLM_L_X10Y135_SLICE_X13Y135_CO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D = CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A = CLBLM_L_X10Y136_SLICE_X12Y136_AO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B = CLBLM_L_X10Y136_SLICE_X12Y136_BO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C = CLBLM_L_X10Y136_SLICE_X12Y136_CO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D = CLBLM_L_X10Y136_SLICE_X12Y136_DO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_AMUX = CLBLM_L_X10Y136_SLICE_X12Y136_AO5;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_BMUX = CLBLM_L_X10Y136_SLICE_X12Y136_BO5;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A = CLBLM_L_X10Y136_SLICE_X13Y136_AO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B = CLBLM_L_X10Y136_SLICE_X13Y136_BO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C = CLBLM_L_X10Y136_SLICE_X13Y136_CO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D = CLBLM_L_X10Y136_SLICE_X13Y136_DO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A = CLBLM_L_X12Y121_SLICE_X16Y121_AO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B = CLBLM_L_X12Y121_SLICE_X16Y121_BO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C = CLBLM_L_X12Y121_SLICE_X16Y121_CO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D = CLBLM_L_X12Y121_SLICE_X16Y121_DO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A = CLBLM_L_X12Y121_SLICE_X17Y121_AO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B = CLBLM_L_X12Y121_SLICE_X17Y121_BO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C = CLBLM_L_X12Y121_SLICE_X17Y121_CO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D = CLBLM_L_X12Y121_SLICE_X17Y121_DO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A = CLBLM_L_X12Y126_SLICE_X16Y126_AO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B = CLBLM_L_X12Y126_SLICE_X16Y126_BO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C = CLBLM_L_X12Y126_SLICE_X16Y126_CO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D = CLBLM_L_X12Y126_SLICE_X16Y126_DO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A = CLBLM_L_X12Y126_SLICE_X17Y126_AO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B = CLBLM_L_X12Y126_SLICE_X17Y126_BO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C = CLBLM_L_X12Y126_SLICE_X17Y126_CO6;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D = CLBLM_L_X12Y126_SLICE_X17Y126_DO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A = CLBLM_L_X12Y127_SLICE_X16Y127_AO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B = CLBLM_L_X12Y127_SLICE_X16Y127_BO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C = CLBLM_L_X12Y127_SLICE_X16Y127_CO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D = CLBLM_L_X12Y127_SLICE_X16Y127_DO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A = CLBLM_L_X12Y127_SLICE_X17Y127_AO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B = CLBLM_L_X12Y127_SLICE_X17Y127_BO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C = CLBLM_L_X12Y127_SLICE_X17Y127_CO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D = CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A = CLBLM_R_X3Y118_SLICE_X2Y118_AO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B = CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D = CLBLM_R_X3Y118_SLICE_X2Y118_DO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_BMUX = CLBLM_R_X3Y118_SLICE_X2Y118_BO5;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_CMUX = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A = CLBLM_R_X3Y118_SLICE_X3Y118_AO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B = CLBLM_R_X3Y118_SLICE_X3Y118_BO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D = CLBLM_R_X3Y118_SLICE_X3Y118_DO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_CMUX = CLBLM_R_X3Y118_SLICE_X3Y118_CO5;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A = CLBLM_R_X3Y119_SLICE_X2Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B = CLBLM_R_X3Y119_SLICE_X2Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C = CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D = CLBLM_R_X3Y119_SLICE_X2Y119_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_CMUX = CLBLM_R_X3Y119_SLICE_X2Y119_CO5;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A = CLBLM_R_X3Y119_SLICE_X3Y119_AO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B = CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C = CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_BMUX = CLBLM_R_X3Y119_SLICE_X3Y119_BO5;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A = CLBLM_R_X3Y120_SLICE_X2Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B = CLBLM_R_X3Y120_SLICE_X2Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C = CLBLM_R_X3Y120_SLICE_X2Y120_CO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D = CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A = CLBLM_R_X3Y120_SLICE_X3Y120_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B = CLBLM_R_X3Y120_SLICE_X3Y120_BO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D = CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A = CLBLM_R_X3Y121_SLICE_X2Y121_AO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B = CLBLM_R_X3Y121_SLICE_X2Y121_BO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C = CLBLM_R_X3Y121_SLICE_X2Y121_CO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D = CLBLM_R_X3Y121_SLICE_X2Y121_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_CMUX = CLBLM_R_X3Y121_SLICE_X2Y121_C5Q;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A = CLBLM_R_X3Y121_SLICE_X3Y121_AO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B = CLBLM_R_X3Y121_SLICE_X3Y121_BO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C = CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D = CLBLM_R_X3Y121_SLICE_X3Y121_DO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_CMUX = CLBLM_R_X3Y121_SLICE_X3Y121_CO5;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A = CLBLM_R_X3Y122_SLICE_X2Y122_AO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B = CLBLM_R_X3Y122_SLICE_X2Y122_BO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C = CLBLM_R_X3Y122_SLICE_X2Y122_CO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D = CLBLM_R_X3Y122_SLICE_X2Y122_DO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_AMUX = CLBLM_R_X3Y122_SLICE_X2Y122_A5Q;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_BMUX = CLBLM_R_X3Y122_SLICE_X2Y122_BO5;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A = CLBLM_R_X3Y122_SLICE_X3Y122_AO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B = CLBLM_R_X3Y122_SLICE_X3Y122_BO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C = CLBLM_R_X3Y122_SLICE_X3Y122_CO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D = CLBLM_R_X3Y122_SLICE_X3Y122_DO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_CMUX = CLBLM_R_X3Y122_SLICE_X3Y122_CO5;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A = CLBLM_R_X3Y123_SLICE_X2Y123_AO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B = CLBLM_R_X3Y123_SLICE_X2Y123_BO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C = CLBLM_R_X3Y123_SLICE_X2Y123_CO6;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D = CLBLM_R_X3Y123_SLICE_X2Y123_DO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A = CLBLM_R_X3Y123_SLICE_X3Y123_AO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B = CLBLM_R_X3Y123_SLICE_X3Y123_BO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C = CLBLM_R_X3Y123_SLICE_X3Y123_CO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D = CLBLM_R_X3Y123_SLICE_X3Y123_DO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A = CLBLM_R_X3Y124_SLICE_X2Y124_AO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B = CLBLM_R_X3Y124_SLICE_X2Y124_BO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C = CLBLM_R_X3Y124_SLICE_X2Y124_CO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D = CLBLM_R_X3Y124_SLICE_X2Y124_DO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_AMUX = CLBLM_R_X3Y124_SLICE_X2Y124_A5Q;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_BMUX = CLBLM_R_X3Y124_SLICE_X2Y124_B5Q;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A = CLBLM_R_X3Y124_SLICE_X3Y124_AO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B = CLBLM_R_X3Y124_SLICE_X3Y124_BO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C = CLBLM_R_X3Y124_SLICE_X3Y124_CO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D = CLBLM_R_X3Y124_SLICE_X3Y124_DO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_CMUX = CLBLM_R_X3Y124_SLICE_X3Y124_C5Q;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A = CLBLM_R_X3Y125_SLICE_X2Y125_AO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B = CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C = CLBLM_R_X3Y125_SLICE_X2Y125_CO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D = CLBLM_R_X3Y125_SLICE_X2Y125_DO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A = CLBLM_R_X3Y125_SLICE_X3Y125_AO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B = CLBLM_R_X3Y125_SLICE_X3Y125_BO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C = CLBLM_R_X3Y125_SLICE_X3Y125_CO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D = CLBLM_R_X3Y125_SLICE_X3Y125_DO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_CMUX = CLBLM_R_X3Y125_SLICE_X3Y125_CO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A = CLBLM_R_X3Y126_SLICE_X2Y126_AO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B = CLBLM_R_X3Y126_SLICE_X2Y126_BO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C = CLBLM_R_X3Y126_SLICE_X2Y126_CO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D = CLBLM_R_X3Y126_SLICE_X2Y126_DO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_AMUX = CLBLM_R_X3Y126_SLICE_X2Y126_A5Q;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_DMUX = CLBLM_R_X3Y126_SLICE_X2Y126_DO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A = CLBLM_R_X3Y126_SLICE_X3Y126_AO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B = CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C = CLBLM_R_X3Y126_SLICE_X3Y126_CO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D = CLBLM_R_X3Y126_SLICE_X3Y126_DO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_BMUX = CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B = CLBLM_R_X3Y127_SLICE_X2Y127_BO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C = CLBLM_R_X3Y127_SLICE_X2Y127_CO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D = CLBLM_R_X3Y127_SLICE_X2Y127_DO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_CMUX = CLBLM_R_X3Y127_SLICE_X2Y127_CO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_DMUX = CLBLM_R_X3Y127_SLICE_X2Y127_DO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A = CLBLM_R_X3Y127_SLICE_X3Y127_AO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B = CLBLM_R_X3Y127_SLICE_X3Y127_BO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C = CLBLM_R_X3Y127_SLICE_X3Y127_CO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D = CLBLM_R_X3Y127_SLICE_X3Y127_DO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_AMUX = CLBLM_R_X3Y127_SLICE_X3Y127_AO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_CMUX = CLBLM_R_X3Y127_SLICE_X3Y127_CO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_A = CLBLM_R_X3Y128_SLICE_X2Y128_AO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_B = CLBLM_R_X3Y128_SLICE_X2Y128_BO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_C = CLBLM_R_X3Y128_SLICE_X2Y128_CO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_D = CLBLM_R_X3Y128_SLICE_X2Y128_DO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_A = CLBLM_R_X3Y128_SLICE_X3Y128_AO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_B = CLBLM_R_X3Y128_SLICE_X3Y128_BO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_C = CLBLM_R_X3Y128_SLICE_X3Y128_CO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_D = CLBLM_R_X3Y128_SLICE_X3Y128_DO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_AMUX = CLBLM_R_X3Y128_SLICE_X3Y128_AO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A = CLBLM_R_X3Y129_SLICE_X2Y129_AO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B = CLBLM_R_X3Y129_SLICE_X2Y129_BO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C = CLBLM_R_X3Y129_SLICE_X2Y129_CO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D = CLBLM_R_X3Y129_SLICE_X2Y129_DO6;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A = CLBLM_R_X3Y129_SLICE_X3Y129_AO6;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B = CLBLM_R_X3Y129_SLICE_X3Y129_BO6;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C = CLBLM_R_X3Y129_SLICE_X3Y129_CO6;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_AMUX = CLBLM_R_X3Y129_SLICE_X3Y129_AO5;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_CMUX = CLBLM_R_X3Y129_SLICE_X3Y129_CO6;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_DMUX = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A = CLBLM_R_X3Y130_SLICE_X2Y130_AO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B = CLBLM_R_X3Y130_SLICE_X2Y130_BO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C = CLBLM_R_X3Y130_SLICE_X2Y130_CO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D = CLBLM_R_X3Y130_SLICE_X2Y130_DO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_AMUX = CLBLM_R_X3Y130_SLICE_X2Y130_AO5;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_BMUX = CLBLM_R_X3Y130_SLICE_X2Y130_BO5;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_DMUX = CLBLM_R_X3Y130_SLICE_X2Y130_DO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A = CLBLM_R_X3Y130_SLICE_X3Y130_AO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B = CLBLM_R_X3Y130_SLICE_X3Y130_BO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C = CLBLM_R_X3Y130_SLICE_X3Y130_CO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D = CLBLM_R_X3Y130_SLICE_X3Y130_DO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_AMUX = CLBLM_R_X3Y130_SLICE_X3Y130_AO5;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A = CLBLM_R_X3Y131_SLICE_X2Y131_AO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B = CLBLM_R_X3Y131_SLICE_X2Y131_BO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C = CLBLM_R_X3Y131_SLICE_X2Y131_CO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D = CLBLM_R_X3Y131_SLICE_X2Y131_DO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_CMUX = CLBLM_R_X3Y131_SLICE_X2Y131_CO5;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A = CLBLM_R_X3Y131_SLICE_X3Y131_AO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B = CLBLM_R_X3Y131_SLICE_X3Y131_BO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C = CLBLM_R_X3Y131_SLICE_X3Y131_CO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D = CLBLM_R_X3Y131_SLICE_X3Y131_DO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A = CLBLM_R_X3Y132_SLICE_X2Y132_AO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B = CLBLM_R_X3Y132_SLICE_X2Y132_BO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C = CLBLM_R_X3Y132_SLICE_X2Y132_CO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D = CLBLM_R_X3Y132_SLICE_X2Y132_DO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_AMUX = CLBLM_R_X3Y132_SLICE_X2Y132_A5Q;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_CMUX = CLBLM_R_X3Y132_SLICE_X2Y132_CO5;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A = CLBLM_R_X3Y132_SLICE_X3Y132_AO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B = CLBLM_R_X3Y132_SLICE_X3Y132_BO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C = CLBLM_R_X3Y132_SLICE_X3Y132_CO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D = CLBLM_R_X3Y132_SLICE_X3Y132_DO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A = CLBLM_R_X5Y116_SLICE_X6Y116_AO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B = CLBLM_R_X5Y116_SLICE_X6Y116_BO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C = CLBLM_R_X5Y116_SLICE_X6Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D = CLBLM_R_X5Y116_SLICE_X6Y116_DO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A = CLBLM_R_X5Y116_SLICE_X7Y116_AO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B = CLBLM_R_X5Y116_SLICE_X7Y116_BO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C = CLBLM_R_X5Y116_SLICE_X7Y116_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_DMUX = CLBLM_R_X5Y116_SLICE_X7Y116_DO5;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A = CLBLM_R_X5Y117_SLICE_X6Y117_AO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B = CLBLM_R_X5Y117_SLICE_X6Y117_BO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C = CLBLM_R_X5Y117_SLICE_X6Y117_CO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D = CLBLM_R_X5Y117_SLICE_X6Y117_DO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_AMUX = CLBLM_R_X5Y117_SLICE_X6Y117_A5Q;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_DMUX = CLBLM_R_X5Y117_SLICE_X6Y117_DO5;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A = CLBLM_R_X5Y117_SLICE_X7Y117_AO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B = CLBLM_R_X5Y117_SLICE_X7Y117_BO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C = CLBLM_R_X5Y117_SLICE_X7Y117_CO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D = CLBLM_R_X5Y117_SLICE_X7Y117_DO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_BMUX = CLBLM_R_X5Y117_SLICE_X7Y117_BO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A = CLBLM_R_X5Y118_SLICE_X6Y118_AO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B = CLBLM_R_X5Y118_SLICE_X6Y118_BO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C = CLBLM_R_X5Y118_SLICE_X6Y118_CO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D = CLBLM_R_X5Y118_SLICE_X6Y118_DO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_AMUX = CLBLM_R_X5Y118_SLICE_X6Y118_AO5;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_BMUX = CLBLM_R_X5Y118_SLICE_X6Y118_B5Q;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_CMUX = CLBLM_R_X5Y118_SLICE_X6Y118_CO5;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A = CLBLM_R_X5Y118_SLICE_X7Y118_AO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B = CLBLM_R_X5Y118_SLICE_X7Y118_BO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D = CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_AMUX = CLBLM_R_X5Y118_SLICE_X7Y118_A5Q;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_BMUX = CLBLM_R_X5Y118_SLICE_X7Y118_BO5;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A = CLBLM_R_X5Y119_SLICE_X6Y119_AO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B = CLBLM_R_X5Y119_SLICE_X6Y119_BO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C = CLBLM_R_X5Y119_SLICE_X6Y119_CO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D = CLBLM_R_X5Y119_SLICE_X6Y119_DO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_BMUX = CLBLM_R_X5Y119_SLICE_X6Y119_BO5;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A = CLBLM_R_X5Y119_SLICE_X7Y119_AO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B = CLBLM_R_X5Y119_SLICE_X7Y119_BO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C = CLBLM_R_X5Y119_SLICE_X7Y119_CO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D = CLBLM_R_X5Y119_SLICE_X7Y119_DO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A = CLBLM_R_X5Y120_SLICE_X6Y120_AO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B = CLBLM_R_X5Y120_SLICE_X6Y120_BO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C = CLBLM_R_X5Y120_SLICE_X6Y120_CO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D = CLBLM_R_X5Y120_SLICE_X6Y120_DO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A = CLBLM_R_X5Y120_SLICE_X7Y120_AO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B = CLBLM_R_X5Y120_SLICE_X7Y120_BO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C = CLBLM_R_X5Y120_SLICE_X7Y120_CO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D = CLBLM_R_X5Y120_SLICE_X7Y120_DO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_AMUX = CLBLM_R_X5Y120_SLICE_X7Y120_A5Q;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A = CLBLM_R_X5Y121_SLICE_X6Y121_AO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B = CLBLM_R_X5Y121_SLICE_X6Y121_BO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C = CLBLM_R_X5Y121_SLICE_X6Y121_CO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D = CLBLM_R_X5Y121_SLICE_X6Y121_DO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_CMUX = CLBLM_R_X5Y121_SLICE_X6Y121_CO5;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A = CLBLM_R_X5Y121_SLICE_X7Y121_AO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B = CLBLM_R_X5Y121_SLICE_X7Y121_BO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C = CLBLM_R_X5Y121_SLICE_X7Y121_CO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D = CLBLM_R_X5Y121_SLICE_X7Y121_DO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_BMUX = CLBLM_R_X5Y121_SLICE_X7Y121_BO5;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A = CLBLM_R_X5Y122_SLICE_X6Y122_AO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B = CLBLM_R_X5Y122_SLICE_X6Y122_BO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C = CLBLM_R_X5Y122_SLICE_X6Y122_CO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D = CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_DMUX = CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A = CLBLM_R_X5Y122_SLICE_X7Y122_AO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B = CLBLM_R_X5Y122_SLICE_X7Y122_BO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C = CLBLM_R_X5Y122_SLICE_X7Y122_CO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D = CLBLM_R_X5Y122_SLICE_X7Y122_DO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A = CLBLM_R_X5Y123_SLICE_X6Y123_AO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B = CLBLM_R_X5Y123_SLICE_X6Y123_BO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C = CLBLM_R_X5Y123_SLICE_X6Y123_CO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D = CLBLM_R_X5Y123_SLICE_X6Y123_DO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_BMUX = CLBLM_R_X5Y123_SLICE_X6Y123_B5Q;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A = CLBLM_R_X5Y123_SLICE_X7Y123_AO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B = CLBLM_R_X5Y123_SLICE_X7Y123_BO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C = CLBLM_R_X5Y123_SLICE_X7Y123_CO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D = CLBLM_R_X5Y123_SLICE_X7Y123_DO6;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_CMUX = CLBLM_R_X5Y123_SLICE_X7Y123_C5Q;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A = CLBLM_R_X5Y124_SLICE_X6Y124_AO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B = CLBLM_R_X5Y124_SLICE_X6Y124_BO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C = CLBLM_R_X5Y124_SLICE_X6Y124_CO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D = CLBLM_R_X5Y124_SLICE_X6Y124_DO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_AMUX = CLBLM_R_X5Y124_SLICE_X6Y124_A5Q;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_DMUX = CLBLM_R_X5Y124_SLICE_X6Y124_DO5;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A = CLBLM_R_X5Y124_SLICE_X7Y124_AO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B = CLBLM_R_X5Y124_SLICE_X7Y124_BO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C = CLBLM_R_X5Y124_SLICE_X7Y124_CO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D = CLBLM_R_X5Y124_SLICE_X7Y124_DO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_CMUX = CLBLM_R_X5Y124_SLICE_X7Y124_C5Q;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A = CLBLM_R_X5Y125_SLICE_X6Y125_AO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B = CLBLM_R_X5Y125_SLICE_X6Y125_BO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C = CLBLM_R_X5Y125_SLICE_X6Y125_CO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D = CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_AMUX = CLBLM_R_X5Y125_SLICE_X6Y125_A5Q;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_CMUX = CLBLM_R_X5Y125_SLICE_X6Y125_CO5;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A = CLBLM_R_X5Y125_SLICE_X7Y125_AO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B = CLBLM_R_X5Y125_SLICE_X7Y125_BO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C = CLBLM_R_X5Y125_SLICE_X7Y125_CO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D = CLBLM_R_X5Y125_SLICE_X7Y125_DO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A = CLBLM_R_X5Y126_SLICE_X6Y126_AO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B = CLBLM_R_X5Y126_SLICE_X6Y126_BO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C = CLBLM_R_X5Y126_SLICE_X6Y126_CO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D = CLBLM_R_X5Y126_SLICE_X6Y126_DO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A = CLBLM_R_X5Y126_SLICE_X7Y126_AO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B = CLBLM_R_X5Y126_SLICE_X7Y126_BO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C = CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D = CLBLM_R_X5Y126_SLICE_X7Y126_DO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_AMUX = CLBLM_R_X5Y126_SLICE_X7Y126_A5Q;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_CMUX = CLBLM_R_X5Y126_SLICE_X7Y126_CO5;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A = CLBLM_R_X5Y127_SLICE_X6Y127_AO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B = CLBLM_R_X5Y127_SLICE_X6Y127_BO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C = CLBLM_R_X5Y127_SLICE_X6Y127_CO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D = CLBLM_R_X5Y127_SLICE_X6Y127_DO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A = CLBLM_R_X5Y127_SLICE_X7Y127_AO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B = CLBLM_R_X5Y127_SLICE_X7Y127_BO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C = CLBLM_R_X5Y127_SLICE_X7Y127_CO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D = CLBLM_R_X5Y127_SLICE_X7Y127_DO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_BMUX = CLBLM_R_X5Y127_SLICE_X7Y127_B5Q;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A = CLBLM_R_X5Y128_SLICE_X6Y128_AO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B = CLBLM_R_X5Y128_SLICE_X6Y128_BO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C = CLBLM_R_X5Y128_SLICE_X6Y128_CO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D = CLBLM_R_X5Y128_SLICE_X6Y128_DO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_AMUX = CLBLM_R_X5Y128_SLICE_X6Y128_A5Q;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_CMUX = CLBLM_R_X5Y128_SLICE_X6Y128_CO5;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A = CLBLM_R_X5Y128_SLICE_X7Y128_AO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B = CLBLM_R_X5Y128_SLICE_X7Y128_BO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C = CLBLM_R_X5Y128_SLICE_X7Y128_CO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D = CLBLM_R_X5Y128_SLICE_X7Y128_DO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_AMUX = CLBLM_R_X5Y128_SLICE_X7Y128_A5Q;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_BMUX = CLBLM_R_X5Y128_SLICE_X7Y128_B5Q;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A = CLBLM_R_X5Y129_SLICE_X6Y129_AO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B = CLBLM_R_X5Y129_SLICE_X6Y129_BO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C = CLBLM_R_X5Y129_SLICE_X6Y129_CO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D = CLBLM_R_X5Y129_SLICE_X6Y129_DO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A = CLBLM_R_X5Y129_SLICE_X7Y129_AO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B = CLBLM_R_X5Y129_SLICE_X7Y129_BO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C = CLBLM_R_X5Y129_SLICE_X7Y129_CO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D = CLBLM_R_X5Y129_SLICE_X7Y129_DO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A = CLBLM_R_X5Y130_SLICE_X6Y130_AO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B = CLBLM_R_X5Y130_SLICE_X6Y130_BO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C = CLBLM_R_X5Y130_SLICE_X6Y130_CO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D = CLBLM_R_X5Y130_SLICE_X6Y130_DO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A = CLBLM_R_X5Y130_SLICE_X7Y130_AO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B = CLBLM_R_X5Y130_SLICE_X7Y130_BO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C = CLBLM_R_X5Y130_SLICE_X7Y130_CO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D = CLBLM_R_X5Y130_SLICE_X7Y130_DO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_CMUX = CLBLM_R_X5Y130_SLICE_X7Y130_CO5;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A = CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B = CLBLM_R_X7Y115_SLICE_X8Y115_BO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C = CLBLM_R_X7Y115_SLICE_X8Y115_CO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D = CLBLM_R_X7Y115_SLICE_X8Y115_DO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_AMUX = CLBLM_R_X7Y115_SLICE_X8Y115_AO5;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A = CLBLM_R_X7Y115_SLICE_X9Y115_AO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B = CLBLM_R_X7Y115_SLICE_X9Y115_BO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C = CLBLM_R_X7Y115_SLICE_X9Y115_CO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D = CLBLM_R_X7Y115_SLICE_X9Y115_DO6;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_AMUX = CLBLM_R_X7Y115_SLICE_X9Y115_AO5;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A = CLBLM_R_X7Y116_SLICE_X8Y116_AO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C = CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_BMUX = CLBLM_R_X7Y116_SLICE_X8Y116_BO5;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A = CLBLM_R_X7Y116_SLICE_X9Y116_AO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B = CLBLM_R_X7Y116_SLICE_X9Y116_BO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C = CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D = CLBLM_R_X7Y116_SLICE_X9Y116_DO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A = CLBLM_R_X7Y117_SLICE_X8Y117_AO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B = CLBLM_R_X7Y117_SLICE_X8Y117_BO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C = CLBLM_R_X7Y117_SLICE_X8Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D = CLBLM_R_X7Y117_SLICE_X8Y117_DO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A = CLBLM_R_X7Y117_SLICE_X9Y117_AO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B = CLBLM_R_X7Y117_SLICE_X9Y117_BO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C = CLBLM_R_X7Y117_SLICE_X9Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D = CLBLM_R_X7Y117_SLICE_X9Y117_DO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_AMUX = CLBLM_R_X7Y117_SLICE_X9Y117_AO5;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_BMUX = CLBLM_R_X7Y117_SLICE_X9Y117_BO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A = CLBLM_R_X7Y118_SLICE_X8Y118_AO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B = CLBLM_R_X7Y118_SLICE_X8Y118_BO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C = CLBLM_R_X7Y118_SLICE_X8Y118_CO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D = CLBLM_R_X7Y118_SLICE_X8Y118_DO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_CMUX = CLBLM_R_X7Y118_SLICE_X8Y118_C5Q;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A = CLBLM_R_X7Y118_SLICE_X9Y118_AO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B = CLBLM_R_X7Y118_SLICE_X9Y118_BO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C = CLBLM_R_X7Y118_SLICE_X9Y118_CO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D = CLBLM_R_X7Y118_SLICE_X9Y118_DO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_BMUX = CLBLM_R_X7Y118_SLICE_X9Y118_BO5;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A = CLBLM_R_X7Y119_SLICE_X8Y119_AO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B = CLBLM_R_X7Y119_SLICE_X8Y119_BO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C = CLBLM_R_X7Y119_SLICE_X8Y119_CO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D = CLBLM_R_X7Y119_SLICE_X8Y119_DO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A = CLBLM_R_X7Y119_SLICE_X9Y119_AO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B = CLBLM_R_X7Y119_SLICE_X9Y119_BO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C = CLBLM_R_X7Y119_SLICE_X9Y119_CO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D = CLBLM_R_X7Y119_SLICE_X9Y119_DO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A = CLBLM_R_X7Y120_SLICE_X8Y120_AO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B = CLBLM_R_X7Y120_SLICE_X8Y120_BO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C = CLBLM_R_X7Y120_SLICE_X8Y120_CO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D = CLBLM_R_X7Y120_SLICE_X8Y120_DO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A = CLBLM_R_X7Y120_SLICE_X9Y120_AO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B = CLBLM_R_X7Y120_SLICE_X9Y120_BO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C = CLBLM_R_X7Y120_SLICE_X9Y120_CO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D = CLBLM_R_X7Y120_SLICE_X9Y120_DO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A = CLBLM_R_X7Y121_SLICE_X8Y121_AO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B = CLBLM_R_X7Y121_SLICE_X8Y121_BO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C = CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_AMUX = CLBLM_R_X7Y121_SLICE_X8Y121_A5Q;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_DMUX = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A = CLBLM_R_X7Y121_SLICE_X9Y121_AO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B = CLBLM_R_X7Y121_SLICE_X9Y121_BO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C = CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D = CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_BMUX = CLBLM_R_X7Y121_SLICE_X9Y121_B5Q;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A = CLBLM_R_X7Y122_SLICE_X8Y122_AO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B = CLBLM_R_X7Y122_SLICE_X8Y122_BO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C = CLBLM_R_X7Y122_SLICE_X8Y122_CO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D = CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_DMUX = CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A = CLBLM_R_X7Y122_SLICE_X9Y122_AO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B = CLBLM_R_X7Y122_SLICE_X9Y122_BO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C = CLBLM_R_X7Y122_SLICE_X9Y122_CO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D = CLBLM_R_X7Y122_SLICE_X9Y122_DO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A = CLBLM_R_X7Y123_SLICE_X8Y123_AO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B = CLBLM_R_X7Y123_SLICE_X8Y123_BO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C = CLBLM_R_X7Y123_SLICE_X8Y123_CO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D = CLBLM_R_X7Y123_SLICE_X8Y123_DO6;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_BMUX = CLBLM_R_X7Y123_SLICE_X8Y123_B5Q;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_CMUX = CLBLM_R_X7Y123_SLICE_X8Y123_CO5;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A = CLBLM_R_X7Y123_SLICE_X9Y123_AO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B = CLBLM_R_X7Y123_SLICE_X9Y123_BO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C = CLBLM_R_X7Y123_SLICE_X9Y123_CO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D = CLBLM_R_X7Y123_SLICE_X9Y123_DO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_AMUX = CLBLM_R_X7Y123_SLICE_X9Y123_A5Q;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_DMUX = CLBLM_R_X7Y123_SLICE_X9Y123_DO5;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A = CLBLM_R_X7Y124_SLICE_X8Y124_AO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B = CLBLM_R_X7Y124_SLICE_X8Y124_BO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C = CLBLM_R_X7Y124_SLICE_X8Y124_CO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D = CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_BMUX = CLBLM_R_X7Y124_SLICE_X8Y124_B5Q;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_CMUX = CLBLM_R_X7Y124_SLICE_X8Y124_CO5;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A = CLBLM_R_X7Y124_SLICE_X9Y124_AO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B = CLBLM_R_X7Y124_SLICE_X9Y124_BO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C = CLBLM_R_X7Y124_SLICE_X9Y124_CO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D = CLBLM_R_X7Y124_SLICE_X9Y124_DO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_BMUX = CLBLM_R_X7Y124_SLICE_X9Y124_BO5;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A = CLBLM_R_X7Y125_SLICE_X8Y125_AO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B = CLBLM_R_X7Y125_SLICE_X8Y125_BO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C = CLBLM_R_X7Y125_SLICE_X8Y125_CO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D = CLBLM_R_X7Y125_SLICE_X8Y125_DO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A = CLBLM_R_X7Y125_SLICE_X9Y125_AO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B = CLBLM_R_X7Y125_SLICE_X9Y125_BO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C = CLBLM_R_X7Y125_SLICE_X9Y125_CO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D = CLBLM_R_X7Y125_SLICE_X9Y125_DO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_AMUX = CLBLM_R_X7Y125_SLICE_X9Y125_A5Q;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_BMUX = CLBLM_R_X7Y125_SLICE_X9Y125_B5Q;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A = CLBLM_R_X7Y126_SLICE_X8Y126_AO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B = CLBLM_R_X7Y126_SLICE_X8Y126_BO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C = CLBLM_R_X7Y126_SLICE_X8Y126_CO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D = CLBLM_R_X7Y126_SLICE_X8Y126_DO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A = CLBLM_R_X7Y126_SLICE_X9Y126_AO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B = CLBLM_R_X7Y126_SLICE_X9Y126_BO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C = CLBLM_R_X7Y126_SLICE_X9Y126_CO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D = CLBLM_R_X7Y126_SLICE_X9Y126_DO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_BMUX = CLBLM_R_X7Y126_SLICE_X9Y126_B5Q;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_CMUX = CLBLM_R_X7Y126_SLICE_X9Y126_C5Q;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_DMUX = CLBLM_R_X7Y126_SLICE_X9Y126_D5Q;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A = CLBLM_R_X7Y127_SLICE_X8Y127_AO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B = CLBLM_R_X7Y127_SLICE_X8Y127_BO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C = CLBLM_R_X7Y127_SLICE_X8Y127_CO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D = CLBLM_R_X7Y127_SLICE_X8Y127_DO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A = CLBLM_R_X7Y127_SLICE_X9Y127_AO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B = CLBLM_R_X7Y127_SLICE_X9Y127_BO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C = CLBLM_R_X7Y127_SLICE_X9Y127_CO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D = CLBLM_R_X7Y127_SLICE_X9Y127_DO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_DMUX = CLBLM_R_X7Y127_SLICE_X9Y127_DO5;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A = CLBLM_R_X7Y128_SLICE_X8Y128_AO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B = CLBLM_R_X7Y128_SLICE_X8Y128_BO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C = CLBLM_R_X7Y128_SLICE_X8Y128_CO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D = CLBLM_R_X7Y128_SLICE_X8Y128_DO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A = CLBLM_R_X7Y128_SLICE_X9Y128_AO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B = CLBLM_R_X7Y128_SLICE_X9Y128_BO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C = CLBLM_R_X7Y128_SLICE_X9Y128_CO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D = CLBLM_R_X7Y128_SLICE_X9Y128_DO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_BMUX = CLBLM_R_X7Y128_SLICE_X9Y128_BO5;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A = CLBLM_R_X7Y129_SLICE_X8Y129_AO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B = CLBLM_R_X7Y129_SLICE_X8Y129_BO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C = CLBLM_R_X7Y129_SLICE_X8Y129_CO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D = CLBLM_R_X7Y129_SLICE_X8Y129_DO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_AMUX = CLBLM_R_X7Y129_SLICE_X8Y129_A5Q;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A = CLBLM_R_X7Y129_SLICE_X9Y129_AO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B = CLBLM_R_X7Y129_SLICE_X9Y129_BO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C = CLBLM_R_X7Y129_SLICE_X9Y129_CO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D = CLBLM_R_X7Y129_SLICE_X9Y129_DO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A = CLBLM_R_X7Y130_SLICE_X8Y130_AO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B = CLBLM_R_X7Y130_SLICE_X8Y130_BO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D = CLBLM_R_X7Y130_SLICE_X8Y130_DO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_CMUX = CLBLM_R_X7Y130_SLICE_X8Y130_CO5;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A = CLBLM_R_X7Y130_SLICE_X9Y130_AO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B = CLBLM_R_X7Y130_SLICE_X9Y130_BO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C = CLBLM_R_X7Y130_SLICE_X9Y130_CO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D = CLBLM_R_X7Y130_SLICE_X9Y130_DO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_BMUX = CLBLM_R_X7Y130_SLICE_X9Y130_BO5;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_CMUX = CLBLM_R_X7Y130_SLICE_X9Y130_CO5;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_DMUX = CLBLM_R_X7Y130_SLICE_X9Y130_DO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A = CLBLM_R_X7Y131_SLICE_X8Y131_AO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B = CLBLM_R_X7Y131_SLICE_X8Y131_BO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C = CLBLM_R_X7Y131_SLICE_X8Y131_CO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D = CLBLM_R_X7Y131_SLICE_X8Y131_DO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_BMUX = CLBLM_R_X7Y131_SLICE_X8Y131_BO5;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_CMUX = CLBLM_R_X7Y131_SLICE_X8Y131_CO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A = CLBLM_R_X7Y131_SLICE_X9Y131_AO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B = CLBLM_R_X7Y131_SLICE_X9Y131_BO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C = CLBLM_R_X7Y131_SLICE_X9Y131_CO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D = CLBLM_R_X7Y131_SLICE_X9Y131_DO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_BMUX = CLBLM_R_X7Y131_SLICE_X9Y131_BO5;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A = CLBLM_R_X11Y119_SLICE_X14Y119_AO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B = CLBLM_R_X11Y119_SLICE_X14Y119_BO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C = CLBLM_R_X11Y119_SLICE_X14Y119_CO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D = CLBLM_R_X11Y119_SLICE_X14Y119_DO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A = CLBLM_R_X11Y119_SLICE_X15Y119_AO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B = CLBLM_R_X11Y119_SLICE_X15Y119_BO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C = CLBLM_R_X11Y119_SLICE_X15Y119_CO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D = CLBLM_R_X11Y119_SLICE_X15Y119_DO6;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_AMUX = CLBLM_R_X11Y119_SLICE_X15Y119_AO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A = CLBLM_R_X11Y120_SLICE_X14Y120_AO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B = CLBLM_R_X11Y120_SLICE_X14Y120_BO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C = CLBLM_R_X11Y120_SLICE_X14Y120_CO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A = CLBLM_R_X11Y120_SLICE_X15Y120_AO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B = CLBLM_R_X11Y120_SLICE_X15Y120_BO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C = CLBLM_R_X11Y120_SLICE_X15Y120_CO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D = CLBLM_R_X11Y120_SLICE_X15Y120_DO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_BMUX = CLBLM_R_X11Y120_SLICE_X15Y120_BO5;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_CMUX = CLBLM_R_X11Y120_SLICE_X15Y120_CO5;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A = CLBLM_R_X11Y121_SLICE_X14Y121_AO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B = CLBLM_R_X11Y121_SLICE_X14Y121_BO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C = CLBLM_R_X11Y121_SLICE_X14Y121_CO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A = CLBLM_R_X11Y121_SLICE_X15Y121_AO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B = CLBLM_R_X11Y121_SLICE_X15Y121_BO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C = CLBLM_R_X11Y121_SLICE_X15Y121_CO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D = CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A = CLBLM_R_X11Y122_SLICE_X14Y122_AO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B = CLBLM_R_X11Y122_SLICE_X14Y122_BO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C = CLBLM_R_X11Y122_SLICE_X14Y122_CO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D = CLBLM_R_X11Y122_SLICE_X14Y122_DO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A = CLBLM_R_X11Y122_SLICE_X15Y122_AO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B = CLBLM_R_X11Y122_SLICE_X15Y122_BO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C = CLBLM_R_X11Y122_SLICE_X15Y122_CO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D = CLBLM_R_X11Y122_SLICE_X15Y122_DO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A = CLBLM_R_X11Y123_SLICE_X14Y123_AO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B = CLBLM_R_X11Y123_SLICE_X14Y123_BO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C = CLBLM_R_X11Y123_SLICE_X14Y123_CO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D = CLBLM_R_X11Y123_SLICE_X14Y123_DO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A = CLBLM_R_X11Y123_SLICE_X15Y123_AO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B = CLBLM_R_X11Y123_SLICE_X15Y123_BO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C = CLBLM_R_X11Y123_SLICE_X15Y123_CO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D = CLBLM_R_X11Y123_SLICE_X15Y123_DO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A = CLBLM_R_X11Y124_SLICE_X14Y124_AO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B = CLBLM_R_X11Y124_SLICE_X14Y124_BO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C = CLBLM_R_X11Y124_SLICE_X14Y124_CO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D = CLBLM_R_X11Y124_SLICE_X14Y124_DO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_AMUX = CLBLM_R_X11Y124_SLICE_X14Y124_A5Q;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_DMUX = CLBLM_R_X11Y124_SLICE_X14Y124_DO5;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A = CLBLM_R_X11Y124_SLICE_X15Y124_AO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B = CLBLM_R_X11Y124_SLICE_X15Y124_BO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C = CLBLM_R_X11Y124_SLICE_X15Y124_CO6;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D = CLBLM_R_X11Y124_SLICE_X15Y124_DO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A = CLBLM_R_X11Y125_SLICE_X14Y125_AO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B = CLBLM_R_X11Y125_SLICE_X14Y125_BO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C = CLBLM_R_X11Y125_SLICE_X14Y125_CO6;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D = CLBLM_R_X11Y125_SLICE_X14Y125_DO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A = CLBLM_R_X11Y125_SLICE_X15Y125_AO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B = CLBLM_R_X11Y125_SLICE_X15Y125_BO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C = CLBLM_R_X11Y125_SLICE_X15Y125_CO6;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D = CLBLM_R_X11Y125_SLICE_X15Y125_DO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A = CLBLM_R_X11Y126_SLICE_X14Y126_AO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B = CLBLM_R_X11Y126_SLICE_X14Y126_BO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C = CLBLM_R_X11Y126_SLICE_X14Y126_CO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D = CLBLM_R_X11Y126_SLICE_X14Y126_DO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_AMUX = CLBLM_R_X11Y126_SLICE_X14Y126_AO5;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A = CLBLM_R_X11Y126_SLICE_X15Y126_AO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B = CLBLM_R_X11Y126_SLICE_X15Y126_BO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C = CLBLM_R_X11Y126_SLICE_X15Y126_CO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D = CLBLM_R_X11Y126_SLICE_X15Y126_DO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_DMUX = CLBLM_R_X11Y126_SLICE_X15Y126_DO5;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A = CLBLM_R_X11Y127_SLICE_X14Y127_AO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B = CLBLM_R_X11Y127_SLICE_X14Y127_BO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C = CLBLM_R_X11Y127_SLICE_X14Y127_CO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D = CLBLM_R_X11Y127_SLICE_X14Y127_DO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_BMUX = CLBLM_R_X11Y127_SLICE_X14Y127_BO5;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A = CLBLM_R_X11Y127_SLICE_X15Y127_AO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B = CLBLM_R_X11Y127_SLICE_X15Y127_BO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C = CLBLM_R_X11Y127_SLICE_X15Y127_CO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D = CLBLM_R_X11Y127_SLICE_X15Y127_DO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_BMUX = CLBLM_R_X11Y127_SLICE_X15Y127_BO5;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_CMUX = CLBLM_R_X11Y127_SLICE_X15Y127_CO5;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_DMUX = CLBLM_R_X11Y127_SLICE_X15Y127_DO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A = CLBLM_R_X11Y128_SLICE_X14Y128_AO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B = CLBLM_R_X11Y128_SLICE_X14Y128_BO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C = CLBLM_R_X11Y128_SLICE_X14Y128_CO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D = CLBLM_R_X11Y128_SLICE_X14Y128_DO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_AMUX = CLBLM_R_X11Y128_SLICE_X14Y128_AO5;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A = CLBLM_R_X11Y128_SLICE_X15Y128_AO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B = CLBLM_R_X11Y128_SLICE_X15Y128_BO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C = CLBLM_R_X11Y128_SLICE_X15Y128_CO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D = CLBLM_R_X11Y128_SLICE_X15Y128_DO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A = CLBLM_R_X11Y129_SLICE_X14Y129_AO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B = CLBLM_R_X11Y129_SLICE_X14Y129_BO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C = CLBLM_R_X11Y129_SLICE_X14Y129_CO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D = CLBLM_R_X11Y129_SLICE_X14Y129_DO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_DMUX = CLBLM_R_X11Y129_SLICE_X14Y129_DO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A = CLBLM_R_X11Y129_SLICE_X15Y129_AO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B = CLBLM_R_X11Y129_SLICE_X15Y129_BO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C = CLBLM_R_X11Y129_SLICE_X15Y129_CO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D = CLBLM_R_X11Y129_SLICE_X15Y129_DO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_AMUX = CLBLM_R_X11Y129_SLICE_X15Y129_AO5;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A = CLBLM_R_X11Y130_SLICE_X14Y130_AO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B = CLBLM_R_X11Y130_SLICE_X14Y130_BO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C = CLBLM_R_X11Y130_SLICE_X14Y130_CO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D = CLBLM_R_X11Y130_SLICE_X14Y130_DO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_BMUX = CLBLM_R_X11Y130_SLICE_X14Y130_BO5;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A = CLBLM_R_X11Y130_SLICE_X15Y130_AO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B = CLBLM_R_X11Y130_SLICE_X15Y130_BO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C = CLBLM_R_X11Y130_SLICE_X15Y130_CO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D = CLBLM_R_X11Y130_SLICE_X15Y130_DO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A = CLBLM_R_X11Y131_SLICE_X14Y131_AO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B = CLBLM_R_X11Y131_SLICE_X14Y131_BO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D = CLBLM_R_X11Y131_SLICE_X14Y131_DO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A = CLBLM_R_X11Y131_SLICE_X15Y131_AO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B = CLBLM_R_X11Y131_SLICE_X15Y131_BO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C = CLBLM_R_X11Y131_SLICE_X15Y131_CO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D = CLBLM_R_X11Y131_SLICE_X15Y131_DO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A = CLBLM_R_X11Y151_SLICE_X14Y151_AO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B = CLBLM_R_X11Y151_SLICE_X14Y151_BO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C = CLBLM_R_X11Y151_SLICE_X14Y151_CO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D = CLBLM_R_X11Y151_SLICE_X14Y151_DO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A = CLBLM_R_X11Y151_SLICE_X15Y151_AO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B = CLBLM_R_X11Y151_SLICE_X15Y151_BO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C = CLBLM_R_X11Y151_SLICE_X15Y151_CO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D = CLBLM_R_X11Y151_SLICE_X15Y151_DO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A = CLBLM_R_X13Y127_SLICE_X18Y127_AO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B = CLBLM_R_X13Y127_SLICE_X18Y127_BO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C = CLBLM_R_X13Y127_SLICE_X18Y127_CO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D = CLBLM_R_X13Y127_SLICE_X18Y127_DO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A = CLBLM_R_X13Y127_SLICE_X19Y127_AO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B = CLBLM_R_X13Y127_SLICE_X19Y127_BO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C = CLBLM_R_X13Y127_SLICE_X19Y127_CO6;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D = CLBLM_R_X13Y127_SLICE_X19Y127_DO6;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_A = CLBLM_R_X103Y140_SLICE_X162Y140_AO6;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_B = CLBLM_R_X103Y140_SLICE_X162Y140_BO6;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_C = CLBLM_R_X103Y140_SLICE_X162Y140_CO6;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_D = CLBLM_R_X103Y140_SLICE_X162Y140_DO6;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_A = CLBLM_R_X103Y140_SLICE_X163Y140_AO6;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_B = CLBLM_R_X103Y140_SLICE_X163Y140_BO6;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_C = CLBLM_R_X103Y140_SLICE_X163Y140_CO6;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_D = CLBLM_R_X103Y140_SLICE_X163Y140_DO6;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_AMUX = CLBLM_R_X103Y140_SLICE_X163Y140_AO5;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A = CLBLM_R_X103Y169_SLICE_X162Y169_AO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B = CLBLM_R_X103Y169_SLICE_X162Y169_BO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C = CLBLM_R_X103Y169_SLICE_X162Y169_CO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D = CLBLM_R_X103Y169_SLICE_X162Y169_DO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B = CLBLM_R_X103Y169_SLICE_X163Y169_BO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C = CLBLM_R_X103Y169_SLICE_X163Y169_CO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D = CLBLM_R_X103Y169_SLICE_X163Y169_DO6;
  assign CLBLM_R_X103Y171_SLICE_X162Y171_A = CLBLM_R_X103Y171_SLICE_X162Y171_AO6;
  assign CLBLM_R_X103Y171_SLICE_X162Y171_B = CLBLM_R_X103Y171_SLICE_X162Y171_BO6;
  assign CLBLM_R_X103Y171_SLICE_X162Y171_C = CLBLM_R_X103Y171_SLICE_X162Y171_CO6;
  assign CLBLM_R_X103Y171_SLICE_X162Y171_D = CLBLM_R_X103Y171_SLICE_X162Y171_DO6;
  assign CLBLM_R_X103Y171_SLICE_X163Y171_A = CLBLM_R_X103Y171_SLICE_X163Y171_AO6;
  assign CLBLM_R_X103Y171_SLICE_X163Y171_B = CLBLM_R_X103Y171_SLICE_X163Y171_BO6;
  assign CLBLM_R_X103Y171_SLICE_X163Y171_C = CLBLM_R_X103Y171_SLICE_X163Y171_CO6;
  assign CLBLM_R_X103Y171_SLICE_X163Y171_D = CLBLM_R_X103Y171_SLICE_X163Y171_DO6;
  assign CLBLM_R_X103Y171_SLICE_X163Y171_AMUX = CLBLM_R_X103Y171_SLICE_X163Y171_AO5;
  assign CLBLM_R_X103Y171_SLICE_X163Y171_BMUX = CLBLM_R_X103Y171_SLICE_X163Y171_BO5;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_A = CLBLM_R_X103Y173_SLICE_X162Y173_AO6;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_B = CLBLM_R_X103Y173_SLICE_X162Y173_BO6;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_C = CLBLM_R_X103Y173_SLICE_X162Y173_CO6;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_D = CLBLM_R_X103Y173_SLICE_X162Y173_DO6;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_A = CLBLM_R_X103Y173_SLICE_X163Y173_AO6;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_B = CLBLM_R_X103Y173_SLICE_X163Y173_BO6;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_C = CLBLM_R_X103Y173_SLICE_X163Y173_CO6;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_D = CLBLM_R_X103Y173_SLICE_X163Y173_DO6;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_AMUX = CLBLM_R_X103Y173_SLICE_X163Y173_AO5;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_A = CLBLM_R_X103Y175_SLICE_X162Y175_AO6;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_B = CLBLM_R_X103Y175_SLICE_X162Y175_BO6;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_C = CLBLM_R_X103Y175_SLICE_X162Y175_CO6;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_D = CLBLM_R_X103Y175_SLICE_X162Y175_DO6;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_A = CLBLM_R_X103Y175_SLICE_X163Y175_AO6;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_B = CLBLM_R_X103Y175_SLICE_X163Y175_BO6;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_C = CLBLM_R_X103Y175_SLICE_X163Y175_CO6;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_D = CLBLM_R_X103Y175_SLICE_X163Y175_DO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A = CLBLM_R_X103Y177_SLICE_X162Y177_AO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B = CLBLM_R_X103Y177_SLICE_X162Y177_BO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C = CLBLM_R_X103Y177_SLICE_X162Y177_CO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D = CLBLM_R_X103Y177_SLICE_X162Y177_DO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B = CLBLM_R_X103Y177_SLICE_X163Y177_BO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C = CLBLM_R_X103Y177_SLICE_X163Y177_CO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D = CLBLM_R_X103Y177_SLICE_X163Y177_DO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_AMUX = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_O = LIOB33_X0Y51_IOB_X0Y51_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_O = LIOB33_X0Y53_IOB_X0Y53_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_O = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_O = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_O = LIOB33_X0Y65_IOB_X0Y65_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_O = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_O = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_O = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_O = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_O = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y73_O = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_O = LIOB33_X0Y75_IOB_X0Y76_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_O = LIOB33_X0Y75_IOB_X0Y75_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_O = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_O = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_O = LIOB33_X0Y79_IOB_X0Y79_I;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_OQ = CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_OQ = CLBLL_L_X2Y117_SLICE_X0Y117_BO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_OQ = CLBLL_L_X2Y118_SLICE_X0Y118_AO5;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_OQ = CLBLL_L_X2Y117_SLICE_X0Y117_AO5;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_OQ = CLBLL_L_X2Y125_SLICE_X1Y125_CO6;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_OQ = CLBLL_L_X2Y117_SLICE_X0Y117_CO5;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_OQ = CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_OQ = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_OQ = CLBLL_L_X2Y118_SLICE_X1Y118_CO5;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_OQ = CLBLM_L_X10Y121_SLICE_X13Y121_B5Q;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_OQ = 1'b0;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_OQ = CLBLM_R_X5Y128_SLICE_X7Y128_BQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_OQ = CLBLM_L_X10Y121_SLICE_X13Y121_BQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_OQ = CLBLL_L_X4Y122_SLICE_X5Y122_CQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_OQ = CLBLL_L_X2Y122_SLICE_X1Y122_AQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = CLBLM_R_X5Y126_SLICE_X7Y126_AQ;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = CLBLM_R_X5Y128_SLICE_X7Y128_B5Q;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = CLBLL_L_X4Y122_SLICE_X5Y122_C5Q;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = CLBLL_L_X4Y118_SLICE_X5Y118_C5Q;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_OQ = CLBLM_R_X3Y125_SLICE_X2Y125_AQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_OQ = CLBLM_L_X8Y123_SLICE_X10Y123_C5Q;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_OQ = CLBLL_L_X2Y118_SLICE_X1Y118_B5Q;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_OQ = CLBLL_L_X4Y126_SLICE_X4Y126_AQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_OQ = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_OQ = CLBLM_R_X3Y123_SLICE_X3Y123_CQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_OQ = CLBLM_R_X3Y123_SLICE_X2Y123_CQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_OQ = CLBLM_R_X3Y132_SLICE_X2Y132_A5Q;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = CLBLM_R_X3Y132_SLICE_X2Y132_BQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_OQ = CLBLM_R_X3Y129_SLICE_X2Y129_AQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = CLBLL_L_X2Y125_SLICE_X1Y125_AQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_OQ = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_OQ = CLBLL_L_X2Y126_SLICE_X1Y126_AQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_OQ = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_OQ = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_OQ = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_OQ = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_OQ = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_OQ = LIOB33_X0Y65_IOB_X0Y65_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_OQ = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_OQ = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_OQ = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_OQ = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_OQ = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_OQ = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_OQ = RIOB33_X105Y109_IOB_X1Y109_I;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_OQ = RIOB33_X105Y107_IOB_X1Y108_I;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_OQ = RIOB33_X105Y113_IOB_X1Y113_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_OQ = RIOB33_X105Y111_IOB_X1Y112_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_OQ = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_OQ = RIOB33_X105Y113_IOB_X1Y114_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_OQ = CLBLM_R_X103Y140_SLICE_X163Y140_AO6;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_OQ = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_OQ = CLBLM_R_X11Y151_SLICE_X14Y151_AO6;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_OQ = CLBLM_R_X103Y140_SLICE_X163Y140_AO5;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_OQ = RIOB33_X105Y127_IOB_X1Y128_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_OQ = RIOB33_X105Y127_IOB_X1Y127_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_OQ = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_OQ = RIOB33_X105Y129_IOB_X1Y129_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_OQ = RIOB33_X105Y131_IOB_X1Y132_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_OQ = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_OQ = RIOB33_X105Y135_IOB_X1Y136_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_OQ = RIOB33_X105Y135_IOB_X1Y135_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_OQ = RIOB33_X105Y143_IOB_X1Y143_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_OQ = RIOB33_X105Y137_IOB_X1Y137_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_OQ = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_OQ = RIOB33_X105Y145_IOB_X1Y146_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_OQ = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_OQ = RIOB33_X105Y147_IOB_X1Y148_I;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_OQ = LIOB33_X0Y69_IOB_X0Y69_I;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_OQ = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_OQ = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_OQ = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_TQ = 1'b1;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ = 1'b1;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_O = LIOB33_X0Y69_IOB_X0Y69_I;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ = CLBLL_L_X2Y117_SLICE_X0Y117_BO5;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ = CLBLL_L_X2Y115_SLICE_X0Y115_AO5;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = CLBLM_L_X10Y120_SLICE_X13Y120_AQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ = CLBLM_R_X5Y118_SLICE_X6Y118_AO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ = RIOB33_X105Y115_IOB_X1Y115_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ = RIOB33_X105Y121_IOB_X1Y122_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_O = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ = CLBLL_L_X4Y118_SLICE_X5Y118_CQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = CLBLM_R_X3Y131_SLICE_X2Y131_BQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = CLBLM_R_X3Y131_SLICE_X2Y131_AQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ = RIOB33_X105Y111_IOB_X1Y111_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ = RIOB33_X105Y109_IOB_X1Y110_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ = RIOB33_X105Y143_IOB_X1Y144_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_O = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_O = RIOB33_X105Y123_IOB_X1Y124_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_O = RIOB33_X105Y135_IOB_X1Y136_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_O = RIOB33_X105Y135_IOB_X1Y135_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_O = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_O = RIOB33_X105Y139_IOB_X1Y139_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_O = RIOB33_X105Y141_IOB_X1Y142_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_O = RIOB33_X105Y141_IOB_X1Y141_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_O = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_O = RIOB33_X105Y145_IOB_X1Y145_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_O = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_O = RIOB33_X105Y147_IOB_X1Y147_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_OQ = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_TQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_OQ = LIOB33_X0Y75_IOB_X0Y76_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_OQ = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_OQ = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_OQ = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_OQ = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_OQ = CLBLM_R_X11Y124_SLICE_X14Y124_DO5;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_OQ = CLBLM_R_X11Y124_SLICE_X14Y124_DO6;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_OQ = CLBLM_L_X10Y126_SLICE_X12Y126_DO5;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_OQ = CLBLM_L_X10Y126_SLICE_X12Y126_DO6;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_OQ = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_OQ = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_OQ = CLBLM_R_X11Y151_SLICE_X14Y151_AO6;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_OQ = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_OQ = CLBLM_R_X103Y171_SLICE_X163Y171_BO6;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_OQ = CLBLM_R_X103Y171_SLICE_X163Y171_AO5;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_OQ = CLBLM_R_X103Y173_SLICE_X163Y173_AO6;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_OQ = CLBLM_R_X103Y171_SLICE_X163Y171_BO5;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_OQ = CLBLM_R_X103Y173_SLICE_X163Y173_AO5;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_OQ = CLBLM_L_X10Y136_SLICE_X12Y136_BO6;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_OQ = CLBLM_R_X11Y124_SLICE_X14Y124_DO6;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_OQ = CLBLM_L_X10Y136_SLICE_X12Y136_AO5;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_OQ = CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_OQ = CLBLM_L_X10Y126_SLICE_X12Y126_DO5;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_OQ = CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_OQ = CLBLM_L_X10Y123_SLICE_X13Y123_DO5;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_OQ = CLBLM_L_X12Y126_SLICE_X16Y126_AQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_OQ = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_OQ = CLBLM_L_X12Y121_SLICE_X16Y121_BQ;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_OQ = CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_OQ = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_OQ = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_OQ = CLBLM_R_X103Y175_SLICE_X163Y175_AO6;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_OQ = CLBLM_R_X103Y175_SLICE_X163Y175_AO6;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_TQ = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ = LIOB33_X0Y75_IOB_X0Y75_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ = CLBLM_R_X11Y131_SLICE_X15Y131_AQ;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O = RIOB33_X105Y119_IOB_X1Y119_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O = RIOB33_X105Y131_IOB_X1Y131_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O = RIOB33_X105Y143_IOB_X1Y144_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O = RIOB33_X105Y143_IOB_X1Y143_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ = CLBLL_L_X36Y124_SLICE_X54Y124_AO6;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ = CLBLM_R_X103Y171_SLICE_X163Y171_AO6;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ = CLBLM_L_X10Y126_SLICE_X12Y126_DO6;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ = CLBLM_R_X11Y124_SLICE_X14Y124_DO5;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ = CLBLM_R_X11Y131_SLICE_X15Y131_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O = RIOB33_X105Y137_IOB_X1Y137_I;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ = CLBLM_L_X10Y123_SLICE_X13Y123_DO5;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ = CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ = 1'b1;
  assign LIOB33_X0Y147_IOB_X0Y148_O = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOB33_X0Y147_IOB_X0Y147_O = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_D1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_T1 = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_D1 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A1 = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A2 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A4 = CLBLM_R_X7Y130_SLICE_X9Y130_BO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A6 = CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B1 = CLBLM_R_X5Y128_SLICE_X6Y128_CO5;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B2 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B3 = CLBLM_L_X8Y129_SLICE_X11Y129_B5Q;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B4 = CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B5 = CLBLM_R_X5Y130_SLICE_X7Y130_CO5;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B6 = CLBLM_L_X8Y131_SLICE_X10Y131_DO6;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_T1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A2 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A3 = CLBLM_R_X3Y119_SLICE_X3Y119_AQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A4 = CLBLM_R_X3Y124_SLICE_X2Y124_AQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C2 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C3 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C4 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B1 = CLBLM_R_X3Y118_SLICE_X3Y118_AQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B2 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B3 = CLBLL_L_X4Y118_SLICE_X5Y118_BQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B4 = CLBLM_R_X3Y118_SLICE_X3Y118_BQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B5 = CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_B6 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C1 = CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C2 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C3 = CLBLM_R_X3Y118_SLICE_X3Y118_AQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C4 = CLBLM_R_X7Y117_SLICE_X9Y117_DO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C5 = CLBLL_L_X4Y118_SLICE_X5Y118_BQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_C6 = CLBLM_R_X3Y118_SLICE_X3Y118_BQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D3 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D4 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A1 = CLBLM_R_X7Y131_SLICE_X9Y131_BO5;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A2 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A4 = CLBLM_R_X7Y129_SLICE_X8Y129_BQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A5 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D1 = CLBLL_L_X2Y127_SLICE_X0Y127_CO6;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D3 = CLBLM_R_X3Y123_SLICE_X3Y123_CQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D4 = CLBLL_L_X4Y120_SLICE_X4Y120_CQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D5 = CLBLM_L_X10Y120_SLICE_X12Y120_AQ;
  assign CLBLM_R_X3Y119_SLICE_X3Y119_D6 = CLBLM_R_X3Y128_SLICE_X3Y128_BO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A6 = CLBLM_R_X5Y119_SLICE_X6Y119_CQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B1 = CLBLM_R_X7Y131_SLICE_X9Y131_BO5;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B2 = CLBLM_L_X10Y129_SLICE_X13Y129_AQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B3 = CLBLM_R_X5Y129_SLICE_X6Y129_AQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B4 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A1 = CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A3 = CLBLM_R_X3Y119_SLICE_X2Y119_AQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A4 = CLBLL_L_X2Y119_SLICE_X1Y119_AQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A5 = CLBLL_L_X4Y119_SLICE_X4Y119_DQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_A6 = CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C2 = CLBLM_R_X5Y129_SLICE_X6Y129_CQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C3 = CLBLM_R_X5Y123_SLICE_X7Y123_AQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B1 = CLBLM_R_X3Y119_SLICE_X2Y119_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B2 = CLBLM_R_X3Y119_SLICE_X2Y119_BQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B3 = CLBLM_R_X3Y119_SLICE_X2Y119_AQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B4 = CLBLM_L_X10Y119_SLICE_X12Y119_CQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_B6 = CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D1 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D2 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C1 = CLBLM_L_X8Y123_SLICE_X11Y123_CQ;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C3 = CLBLL_L_X2Y118_SLICE_X1Y118_B5Q;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C4 = CLBLL_L_X2Y118_SLICE_X1Y118_A5Q;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C5 = CLBLM_R_X5Y120_SLICE_X7Y120_A5Q;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_C6 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D3 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D4 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D5 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D6 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D1 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D2 = CLBLM_R_X7Y117_SLICE_X9Y117_DO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D3 = CLBLM_R_X3Y119_SLICE_X3Y119_BO5;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D4 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D5 = 1'b1;
  assign CLBLM_R_X3Y119_SLICE_X2Y119_D6 = CLBLL_L_X2Y119_SLICE_X1Y119_AQ;
  assign RIOB33_X105Y157_IOB_X1Y158_O = CLBLL_L_X36Y124_SLICE_X54Y124_AO6;
  assign RIOB33_X105Y157_IOB_X1Y157_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B2 = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1 = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOB33_X0Y151_IOB_X0Y152_O = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOB33_X0Y151_IOB_X0Y151_O = LIOB33_X0Y65_IOB_X0Y65_I;
  assign RIOB33_SING_X105Y199_IOB_X1Y199_O = CLBLM_R_X11Y131_SLICE_X15Y131_AQ;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C4 = 1'b1;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_D = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_D = RIOB33_X105Y139_IOB_X1Y139_I;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_D = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_D = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A2 = CLBLM_R_X7Y129_SLICE_X9Y129_CQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A3 = CLBLM_R_X5Y130_SLICE_X7Y130_AQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A4 = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A5 = CLBLM_R_X5Y130_SLICE_X7Y130_BQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A6 = CLBLM_R_X5Y130_SLICE_X7Y130_CO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B1 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B2 = CLBLM_R_X7Y129_SLICE_X9Y129_CQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B4 = CLBLM_R_X7Y128_SLICE_X8Y128_BQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B5 = CLBLM_R_X5Y130_SLICE_X7Y130_BQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B6 = CLBLM_R_X5Y130_SLICE_X7Y130_CO6;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_D1 = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A2 = CLBLL_L_X4Y117_SLICE_X4Y117_AO5;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A3 = CLBLM_R_X3Y120_SLICE_X3Y120_AQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A4 = CLBLL_L_X4Y120_SLICE_X4Y120_BQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A5 = CLBLM_R_X3Y126_SLICE_X3Y126_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C1 = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C2 = CLBLM_R_X5Y130_SLICE_X7Y130_AQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C3 = CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B1 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B3 = CLBLM_R_X3Y120_SLICE_X3Y120_AQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B4 = CLBLM_R_X5Y121_SLICE_X7Y121_AQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_B6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D1 = CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C2 = CLBLL_L_X4Y125_SLICE_X4Y125_BQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C3 = CLBLM_R_X3Y119_SLICE_X3Y119_DO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C4 = CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C5 = CLBLM_R_X3Y120_SLICE_X3Y120_DO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_C6 = CLBLM_R_X3Y127_SLICE_X2Y127_DO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D3 = CLBLM_R_X5Y130_SLICE_X7Y130_BQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D4 = CLBLM_L_X8Y129_SLICE_X11Y129_B5Q;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A1 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A2 = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A3 = CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A5 = CLBLM_R_X5Y120_SLICE_X6Y120_BQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D1 = CLBLM_R_X3Y126_SLICE_X3Y126_AO6;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D2 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D3 = CLBLM_R_X3Y121_SLICE_X2Y121_CQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D4 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D5 = CLBLM_R_X3Y125_SLICE_X2Y125_AQ;
  assign CLBLM_R_X3Y120_SLICE_X3Y120_D6 = CLBLM_R_X3Y130_SLICE_X3Y130_BO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A6 = CLBLM_R_X5Y130_SLICE_X6Y130_CO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B1 = CLBLM_L_X8Y131_SLICE_X10Y131_DO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B2 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A1 = CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A3 = CLBLM_R_X3Y120_SLICE_X2Y120_AQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A4 = CLBLM_R_X3Y121_SLICE_X3Y121_BQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A5 = CLBLM_R_X3Y118_SLICE_X3Y118_AQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_A6 = CLBLL_L_X4Y125_SLICE_X4Y125_BQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C1 = CLBLM_R_X5Y130_SLICE_X7Y130_AQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C2 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C3 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B1 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B2 = CLBLM_R_X3Y120_SLICE_X2Y120_BQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B3 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B5 = CLBLL_L_X4Y120_SLICE_X4Y120_C5Q;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D1 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D2 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C1 = CLBLL_L_X4Y120_SLICE_X4Y120_BQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C2 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C3 = CLBLL_L_X2Y121_SLICE_X1Y121_B5Q;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C5 = CLBLM_R_X3Y120_SLICE_X2Y120_DO6;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D5 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D6 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D2 = CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D1 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D2 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D3 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D5 = 1'b1;
  assign CLBLM_R_X3Y120_SLICE_X2Y120_D6 = CLBLM_R_X5Y124_SLICE_X6Y124_CQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D5 = CLBLM_R_X11Y129_SLICE_X14Y129_BQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D6 = CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  assign LIOB33_X0Y153_IOB_X0Y154_O = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOB33_X0Y153_IOB_X0Y153_O = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C3 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C4 = CLBLM_L_X8Y129_SLICE_X11Y129_B5Q;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C5 = CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C6 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B4 = CLBLM_L_X10Y128_SLICE_X13Y128_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B5 = CLBLM_R_X11Y130_SLICE_X14Y130_BO5;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B6 = CLBLM_R_X11Y128_SLICE_X14Y128_CO6;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_A3 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_A4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_A5 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D1 = CLBLM_R_X7Y130_SLICE_X9Y130_CO5;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C1 = CLBLM_L_X12Y127_SLICE_X16Y127_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D2 = CLBLM_R_X7Y128_SLICE_X9Y128_CO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C2 = CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D3 = CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C3 = CLBLM_R_X11Y129_SLICE_X14Y129_BQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A1 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A2 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A3 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D4 = CLBLM_R_X7Y130_SLICE_X9Y130_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C4 = CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A4 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A5 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A6 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D5 = CLBLM_R_X7Y131_SLICE_X9Y131_BO5;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C5 = CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B1 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B2 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D6 = CLBLM_R_X5Y129_SLICE_X6Y129_BQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_C6 = CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B3 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B4 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B5 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B6 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C1 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C2 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C3 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C4 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C5 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C6 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D1 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D2 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D3 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D4 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D5 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D6 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A1 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A2 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A3 = CLBLM_R_X11Y124_SLICE_X14Y124_A5Q;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A4 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A5 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A6 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B1 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A1 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A2 = CLBLM_R_X5Y123_SLICE_X7Y123_BQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A3 = CLBLM_R_X3Y121_SLICE_X3Y121_AQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A5 = CLBLM_R_X3Y121_SLICE_X3Y121_CO5;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_A6 = CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B2 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B3 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B4 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B1 = CLBLM_R_X3Y121_SLICE_X3Y121_DO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B2 = CLBLM_R_X3Y121_SLICE_X3Y121_BQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B4 = CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B5 = CLBLM_R_X3Y121_SLICE_X3Y121_CO5;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_B6 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D1 = CLBLM_L_X12Y127_SLICE_X16Y127_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D2 = CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C1 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C2 = CLBLM_R_X5Y122_SLICE_X7Y122_AQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C3 = CLBLM_R_X3Y121_SLICE_X3Y121_BQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C4 = CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C5 = CLBLM_R_X3Y121_SLICE_X3Y121_AQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_C6 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A6 = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D1 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D2 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D3 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D5 = CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D4 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D1 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D2 = CLBLM_R_X5Y122_SLICE_X7Y122_AQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D3 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D4 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D5 = CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  assign CLBLM_R_X3Y121_SLICE_X3Y121_D6 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A1 = CLBLL_L_X2Y121_SLICE_X1Y121_AO5;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A2 = CLBLM_R_X3Y120_SLICE_X2Y120_BQ;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A3 = CLBLM_R_X3Y121_SLICE_X2Y121_AQ;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A5 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_A6 = CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B1 = CLBLL_L_X2Y121_SLICE_X1Y121_AO5;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B3 = CLBLM_R_X3Y121_SLICE_X2Y121_AQ;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B4 = CLBLL_L_X2Y121_SLICE_X1Y121_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B5 = CLBLM_L_X10Y125_SLICE_X13Y125_BQ;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_B6 = CLBLM_R_X3Y121_SLICE_X2Y121_BQ;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_D1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C1 = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C2 = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C4 = CLBLM_L_X10Y120_SLICE_X12Y120_CQ;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C5 = CLBLM_R_X3Y121_SLICE_X2Y121_DO6;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_C6 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_T1 = 1'b1;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D1 = CLBLM_R_X3Y121_SLICE_X2Y121_C5Q;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D2 = CLBLL_L_X2Y121_SLICE_X0Y121_BQ;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D3 = CLBLM_R_X3Y121_SLICE_X2Y121_BQ;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D4 = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D5 = CLBLM_R_X3Y121_SLICE_X2Y121_AQ;
  assign CLBLM_R_X3Y121_SLICE_X2Y121_D6 = CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_D1 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_T1 = 1'b1;
  assign LIOB33_X0Y155_IOB_X0Y156_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOB33_X0Y155_IOB_X0Y155_O = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C3 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C4 = CLBLM_R_X5Y130_SLICE_X7Y130_CO5;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C5 = CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1 = CLBLM_R_X11Y131_SLICE_X15Y131_AQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D2 = CLBLM_R_X3Y128_SLICE_X2Y128_AO6;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D5 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1 = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1 = 1'b1;
  assign RIOB33_X105Y181_IOB_X1Y182_O = CLBLM_L_X10Y126_SLICE_X12Y126_DO6;
  assign RIOB33_X105Y181_IOB_X1Y181_O = CLBLM_R_X11Y124_SLICE_X14Y124_DO5;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_D = RIOB33_X105Y141_IOB_X1Y142_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_D = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A1 = CLBLM_R_X5Y123_SLICE_X6Y123_B5Q;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A2 = CLBLL_L_X4Y125_SLICE_X4Y125_BQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A4 = CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A5 = CLBLM_R_X3Y121_SLICE_X3Y121_AQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_A6 = CLBLM_R_X3Y122_SLICE_X3Y122_AQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B1 = CLBLM_R_X5Y120_SLICE_X6Y120_DQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B2 = CLBLM_R_X3Y122_SLICE_X3Y122_BQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B3 = CLBLM_R_X3Y123_SLICE_X3Y123_AQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B5 = CLBLM_R_X7Y123_SLICE_X9Y123_A5Q;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_B6 = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C1 = CLBLM_R_X3Y121_SLICE_X3Y121_AQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C2 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C3 = CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C4 = CLBLM_R_X3Y121_SLICE_X3Y121_BQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C5 = CLBLM_R_X5Y122_SLICE_X7Y122_AQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_C6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A1 = CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_D2 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_D3 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_D4 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D2 = CLBLL_L_X2Y129_SLICE_X0Y129_AO6;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D1 = CLBLM_R_X3Y121_SLICE_X3Y121_AQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D2 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D3 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D4 = CLBLM_R_X3Y122_SLICE_X2Y122_CQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D5 = CLBLM_R_X5Y123_SLICE_X7Y123_BQ;
  assign CLBLM_R_X3Y122_SLICE_X3Y122_D6 = CLBLM_R_X3Y121_SLICE_X3Y121_BQ;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_D5 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_D6 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A1 = CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A2 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A3 = CLBLM_R_X3Y122_SLICE_X2Y122_AQ;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A4 = CLBLL_L_X4Y122_SLICE_X5Y122_CQ;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_A6 = CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A2 = CLBLM_R_X5Y117_SLICE_X6Y117_CQ;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_AX = CLBLM_R_X3Y122_SLICE_X2Y122_BO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D3 = CLBLM_L_X10Y121_SLICE_X12Y121_C5Q;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B1 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B4 = CLBLL_L_X2Y126_SLICE_X1Y126_AQ;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B5 = CLBLM_R_X7Y122_SLICE_X8Y122_DO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_B6 = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_T1 = 1'b1;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C1 = CLBLM_L_X10Y121_SLICE_X12Y121_C5Q;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C2 = CLBLM_R_X3Y122_SLICE_X2Y122_CQ;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C3 = CLBLM_R_X5Y123_SLICE_X7Y123_BQ;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C4 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C5 = CLBLM_R_X3Y122_SLICE_X2Y122_BO5;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A3 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign LIOB33_X0Y157_IOB_X0Y157_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign LIOB33_X0Y157_IOB_X0Y158_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D4 = CLBLL_L_X4Y121_SLICE_X4Y121_AQ;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D1 = CLBLM_R_X7Y123_SLICE_X9Y123_A5Q;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D2 = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D3 = CLBLM_R_X3Y122_SLICE_X2Y122_DQ;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D4 = CLBLM_R_X5Y122_SLICE_X7Y122_AQ;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D5 = CLBLM_R_X3Y121_SLICE_X3Y121_BQ;
  assign CLBLM_R_X3Y122_SLICE_X2Y122_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D5 = CLBLL_L_X4Y126_SLICE_X4Y126_BO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D6 = CLBLM_R_X3Y125_SLICE_X3Y125_AQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_A6 = CLBLM_L_X10Y120_SLICE_X12Y120_CQ;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_D1 = CLBLM_R_X11Y124_SLICE_X14Y124_DO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A1 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A3 = CLBLM_R_X3Y123_SLICE_X3Y123_AQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A4 = CLBLM_R_X3Y125_SLICE_X3Y125_AQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A5 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_A6 = CLBLM_R_X3Y121_SLICE_X3Y121_CO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B1 = CLBLM_R_X3Y123_SLICE_X3Y123_DO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B2 = CLBLM_R_X3Y122_SLICE_X3Y122_DO6;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B3 = CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B4 = CLBLM_R_X5Y126_SLICE_X7Y126_BQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B5 = CLBLM_R_X3Y122_SLICE_X3Y122_CO5;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C1 = CLBLM_R_X5Y124_SLICE_X7Y124_C5Q;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C3 = CLBLM_R_X3Y121_SLICE_X2Y121_C5Q;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C4 = CLBLL_L_X2Y121_SLICE_X0Y121_BQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C5 = CLBLM_R_X3Y121_SLICE_X2Y121_AQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_C6 = CLBLM_R_X3Y121_SLICE_X2Y121_BQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D1 = CLBLL_L_X4Y120_SLICE_X5Y120_BQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D2 = CLBLM_R_X3Y123_SLICE_X3Y123_AQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D3 = CLBLM_R_X5Y123_SLICE_X6Y123_B5Q;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D4 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D5 = CLBLL_L_X4Y120_SLICE_X5Y120_AQ;
  assign CLBLM_R_X3Y123_SLICE_X3Y123_D6 = 1'b1;
  assign LIOB33_X0Y159_IOB_X0Y160_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOB33_X0Y159_IOB_X0Y159_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A1 = CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A2 = CLBLL_L_X4Y125_SLICE_X4Y125_BQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A3 = CLBLM_R_X3Y123_SLICE_X2Y123_AQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A4 = CLBLM_R_X3Y122_SLICE_X2Y122_AQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A5 = CLBLM_R_X3Y122_SLICE_X2Y122_CQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B1 = CLBLM_R_X3Y122_SLICE_X2Y122_DQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B2 = CLBLM_R_X3Y123_SLICE_X2Y123_BQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B3 = CLBLM_R_X5Y126_SLICE_X7Y126_CO5;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B4 = 1'b1;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B5 = CLBLL_L_X4Y120_SLICE_X4Y120_BQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C2 = CLBLM_R_X3Y123_SLICE_X2Y123_CQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C3 = CLBLL_L_X2Y118_SLICE_X1Y118_AQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C4 = CLBLM_R_X3Y132_SLICE_X2Y132_A5Q;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_C6 = CLBLM_R_X5Y117_SLICE_X6Y117_A5Q;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D1 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D2 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D3 = CLBLM_R_X3Y123_SLICE_X2Y123_DQ;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D4 = CLBLM_R_X3Y132_SLICE_X2Y132_A5Q;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X3Y123_SLICE_X2Y123_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D5 = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_D1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_T1 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_D1 = CLBLL_L_X2Y117_SLICE_X0Y117_BO6;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_D1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_T1 = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_T1 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_D1 = CLBLL_L_X2Y118_SLICE_X0Y118_AO5;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_T1 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A3 = CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A1 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A2 = CLBLL_L_X4Y124_SLICE_X4Y124_AQ;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A3 = CLBLM_R_X3Y124_SLICE_X3Y124_AQ;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A5 = CLBLM_L_X8Y124_SLICE_X11Y124_BQ;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_A6 = CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A4 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B1 = CLBLM_R_X5Y126_SLICE_X7Y126_CO5;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B2 = CLBLM_R_X3Y124_SLICE_X3Y124_BQ;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B3 = CLBLM_R_X3Y124_SLICE_X3Y124_AQ;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B4 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_B6 = CLBLL_L_X4Y121_SLICE_X4Y121_DQ;
  assign LIOB33_X0Y161_IOB_X0Y161_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign LIOB33_X0Y161_IOB_X0Y162_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C3 = CLBLL_L_X4Y120_SLICE_X5Y120_A5Q;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C4 = CLBLM_R_X3Y124_SLICE_X2Y124_CQ;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C5 = CLBLL_L_X4Y124_SLICE_X4Y124_A5Q;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_C6 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D1 = CLBLM_R_X3Y125_SLICE_X3Y125_CO6;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D3 = CLBLM_R_X3Y124_SLICE_X2Y124_B5Q;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D4 = CLBLL_L_X4Y123_SLICE_X5Y123_B5Q;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D5 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X3Y124_D6 = CLBLM_R_X5Y125_SLICE_X6Y125_A5Q;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A1 = CLBLM_R_X3Y124_SLICE_X2Y124_CQ;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A2 = CLBLM_R_X3Y127_SLICE_X2Y127_DO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A4 = CLBLM_R_X3Y128_SLICE_X3Y128_BO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A5 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_A6 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B1 = CLBLL_L_X2Y118_SLICE_X1Y118_AQ;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B2 = CLBLM_R_X5Y123_SLICE_X6Y123_AQ;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B4 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B5 = CLBLM_R_X3Y126_SLICE_X3Y126_AO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_B6 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C2 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C3 = CLBLL_L_X4Y121_SLICE_X4Y121_BQ;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C5 = CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_C6 = CLBLL_L_X4Y125_SLICE_X4Y125_BQ;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D2 = CLBLL_L_X4Y120_SLICE_X5Y120_A5Q;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D3 = CLBLM_R_X3Y124_SLICE_X2Y124_DQ;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D4 = 1'b1;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D5 = CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  assign CLBLM_R_X3Y124_SLICE_X2Y124_D6 = CLBLM_R_X3Y132_SLICE_X2Y132_BQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B5 = CLBLM_R_X5Y126_SLICE_X7Y126_CO5;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_D = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_D = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_D = LIOB33_X0Y63_IOB_X0Y64_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B5 = CLBLL_L_X4Y118_SLICE_X4Y118_AQ;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B6 = CLBLM_L_X8Y121_SLICE_X10Y121_BQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B6 = CLBLM_R_X5Y122_SLICE_X6Y122_CQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B1 = CLBLM_R_X7Y118_SLICE_X8Y118_DQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D5 = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D5 = CLBLL_L_X4Y123_SLICE_X4Y123_BQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D6 = CLBLL_L_X4Y124_SLICE_X4Y124_AQ;
  assign LIOB33_X0Y163_IOB_X0Y164_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign LIOB33_X0Y163_IOB_X0Y163_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A1 = CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A2 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A3 = CLBLM_R_X3Y125_SLICE_X3Y125_AQ;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A4 = CLBLL_L_X4Y125_SLICE_X4Y125_AQ;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_A6 = CLBLL_L_X2Y121_SLICE_X0Y121_BQ;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B1 = CLBLM_R_X5Y122_SLICE_X6Y122_CQ;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B2 = CLBLM_R_X3Y125_SLICE_X3Y125_BQ;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B4 = CLBLL_L_X2Y125_SLICE_X1Y125_AQ;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_B6 = CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C3 = CLBLM_L_X12Y126_SLICE_X16Y126_BQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C4 = CLBLM_L_X10Y129_SLICE_X13Y129_BO5;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C1 = CLBLM_R_X5Y127_SLICE_X7Y127_B5Q;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C2 = CLBLM_R_X7Y126_SLICE_X9Y126_D5Q;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C3 = CLBLM_R_X3Y126_SLICE_X2Y126_A5Q;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C4 = CLBLL_L_X2Y122_SLICE_X1Y122_A5Q;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C5 = CLBLM_R_X5Y123_SLICE_X7Y123_C5Q;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_C6 = CLBLL_L_X2Y121_SLICE_X1Y121_BQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C5 = CLBLM_L_X10Y128_SLICE_X13Y128_AQ;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C6 = CLBLM_R_X11Y129_SLICE_X14Y129_BQ;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D1 = CLBLM_R_X3Y124_SLICE_X3Y124_AQ;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D2 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D3 = CLBLL_L_X4Y126_SLICE_X4Y126_BO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D4 = CLBLL_L_X2Y129_SLICE_X0Y129_AO6;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X3Y125_D6 = CLBLM_R_X3Y120_SLICE_X2Y120_AQ;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A1 = CLBLL_L_X2Y126_SLICE_X1Y126_AQ;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A2 = CLBLM_R_X3Y130_SLICE_X2Y130_AO5;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A3 = CLBLL_L_X2Y118_SLICE_X1Y118_AQ;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A4 = CLBLM_R_X3Y122_SLICE_X2Y122_CQ;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_A6 = CLBLL_L_X2Y125_SLICE_X1Y125_AQ;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B1 = CLBLM_R_X3Y125_SLICE_X2Y125_DO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B2 = CLBLM_R_X3Y126_SLICE_X2Y126_BO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B3 = CLBLM_R_X5Y127_SLICE_X7Y127_B5Q;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B4 = CLBLM_R_X7Y126_SLICE_X9Y126_D5Q;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_B6 = CLBLL_L_X2Y125_SLICE_X1Y125_DO6;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C1 = CLBLL_L_X2Y121_SLICE_X1Y121_BQ;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C2 = CLBLM_R_X5Y123_SLICE_X7Y123_C5Q;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C4 = CLBLM_R_X3Y124_SLICE_X2Y124_B5Q;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C5 = CLBLM_R_X5Y127_SLICE_X7Y127_B5Q;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_C6 = CLBLM_R_X7Y126_SLICE_X9Y126_D5Q;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D1 = CLBLM_R_X5Y123_SLICE_X7Y123_C5Q;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D2 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D3 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D4 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D5 = 1'b1;
  assign CLBLM_R_X3Y125_SLICE_X2Y125_D6 = CLBLM_R_X3Y124_SLICE_X2Y124_B5Q;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D5 = CLBLM_L_X12Y127_SLICE_X16Y127_AQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D6 = CLBLM_R_X11Y129_SLICE_X14Y129_BQ;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D6 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C3 = CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C4 = CLBLM_R_X5Y130_SLICE_X7Y130_CO5;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C5 = CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C6 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B5 = CLBLM_L_X10Y125_SLICE_X13Y125_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C2 = CLBLM_L_X10Y123_SLICE_X13Y123_CQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B6 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C3 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D2 = CLBLM_L_X8Y129_SLICE_X11Y129_B5Q;
  assign LIOB33_X0Y165_IOB_X0Y166_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign LIOB33_X0Y165_IOB_X0Y165_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C4 = CLBLM_L_X12Y127_SLICE_X16Y127_AQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D5 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C5 = CLBLM_L_X10Y129_SLICE_X13Y129_CO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D6 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C6 = CLBLM_L_X10Y129_SLICE_X13Y129_BO5;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_D1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_T1 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_D1 = CLBLL_L_X2Y117_SLICE_X0Y117_AO5;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1 = CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A1 = CLBLM_R_X3Y126_SLICE_X3Y126_DO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A2 = CLBLM_R_X3Y126_SLICE_X2Y126_DO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A3 = CLBLL_L_X2Y129_SLICE_X1Y129_CO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A4 = CLBLL_L_X4Y127_SLICE_X5Y127_AO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A5 = CLBLL_L_X4Y125_SLICE_X4Y125_DO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_A6 = CLBLL_L_X2Y126_SLICE_X1Y126_DO6;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_D1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_D1 = CLBLM_R_X11Y151_SLICE_X14Y151_AO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B1 = CLBLM_R_X7Y126_SLICE_X8Y126_AQ;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B2 = CLBLM_R_X3Y127_SLICE_X3Y127_CO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B3 = CLBLM_R_X3Y122_SLICE_X3Y122_AQ;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B4 = CLBLL_L_X4Y126_SLICE_X4Y126_BO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B5 = CLBLL_L_X2Y129_SLICE_X0Y129_AO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_B6 = CLBLM_R_X3Y126_SLICE_X3Y126_CO6;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_T1 = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_T1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C1 = CLBLL_L_X2Y130_SLICE_X0Y130_BO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C2 = CLBLL_L_X2Y130_SLICE_X0Y130_CO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C3 = CLBLM_R_X5Y126_SLICE_X6Y126_DQ;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C4 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C5 = CLBLL_L_X2Y125_SLICE_X1Y125_CO5;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_C6 = CLBLL_L_X2Y128_SLICE_X1Y128_AO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D2 = CLBLM_R_X11Y126_SLICE_X14Y126_DQ;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_D1 = CLBLL_L_X2Y125_SLICE_X1Y125_CO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D3 = CLBLM_L_X12Y127_SLICE_X16Y127_AQ;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_T1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D1 = CLBLM_R_X3Y130_SLICE_X3Y130_AO6;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D2 = CLBLM_L_X10Y128_SLICE_X12Y128_DQ;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D3 = CLBLL_L_X4Y126_SLICE_X4Y126_BO5;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D4 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D5 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X3Y126_D6 = CLBLM_R_X3Y120_SLICE_X3Y120_AQ;
  assign RIOB33_X105Y197_IOB_X1Y198_O = CLBLM_R_X103Y175_SLICE_X163Y175_AO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A3 = CLBLM_R_X3Y126_SLICE_X2Y126_AQ;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A4 = CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A5 = CLBLM_R_X3Y126_SLICE_X2Y126_A5Q;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_A6 = CLBLM_R_X3Y124_SLICE_X2Y124_A5Q;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_AX = CLBLM_R_X3Y130_SLICE_X2Y130_AO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B1 = CLBLM_R_X3Y129_SLICE_X2Y129_CO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B2 = CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B3 = CLBLM_R_X3Y126_SLICE_X3Y126_AO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B4 = CLBLM_R_X3Y128_SLICE_X3Y128_BO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B5 = CLBLL_L_X4Y128_SLICE_X4Y128_AO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_B6 = CLBLL_L_X2Y127_SLICE_X1Y127_CO6;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C1 = CLBLM_R_X3Y124_SLICE_X2Y124_AQ;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C2 = CLBLM_R_X3Y126_SLICE_X2Y126_AQ;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C3 = CLBLL_L_X2Y130_SLICE_X0Y130_CO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C4 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_C6 = CLBLL_L_X2Y128_SLICE_X1Y128_AO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B4 = CLBLM_L_X8Y129_SLICE_X11Y129_B5Q;
  assign RIOB33_X105Y197_IOB_X1Y197_O = CLBLM_R_X103Y175_SLICE_X163Y175_AO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B5 = CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B6 = 1'b1;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D1 = CLBLL_L_X2Y126_SLICE_X0Y126_AO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D2 = CLBLL_L_X4Y119_SLICE_X4Y119_DQ;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D3 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D4 = CLBLL_L_X2Y130_SLICE_X1Y130_BO6;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D5 = CLBLL_L_X2Y126_SLICE_X0Y126_AO5;
  assign CLBLM_R_X3Y126_SLICE_X2Y126_D6 = CLBLL_L_X4Y124_SLICE_X5Y124_DQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A1 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A2 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A3 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A4 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A5 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_A6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C5 = CLBLM_L_X8Y124_SLICE_X11Y124_DO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B1 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B2 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C6 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B3 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B4 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B5 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_B6 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C1 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C2 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C3 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C4 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C5 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_C6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C2 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C3 = CLBLM_L_X8Y131_SLICE_X10Y131_DO6;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D1 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D2 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D3 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D4 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D5 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X17Y121_D6 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C4 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C5 = CLBLM_R_X7Y131_SLICE_X8Y131_BO5;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A2 = CLBLM_L_X12Y121_SLICE_X16Y121_BQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A3 = CLBLM_L_X12Y121_SLICE_X16Y121_AQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A4 = CLBLM_R_X11Y121_SLICE_X15Y121_CO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A5 = CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C6 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B2 = CLBLM_L_X12Y121_SLICE_X16Y121_BQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B3 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B4 = CLBLM_L_X10Y120_SLICE_X13Y120_A5Q;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B5 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_B6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D2 = CLBLM_R_X3Y123_SLICE_X2Y123_DQ;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C1 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C2 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C3 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C4 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C5 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_C6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D3 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D4 = CLBLM_R_X3Y128_SLICE_X2Y128_AO6;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D5 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D1 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D2 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D3 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D4 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D5 = 1'b1;
  assign CLBLM_L_X12Y121_SLICE_X16Y121_D6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_D6 = CLBLM_R_X5Y125_SLICE_X6Y125_CO6;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_A1 = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_A3 = RIOB33_X105Y137_IOB_X1Y138_I;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_A4 = RIOB33_X105Y139_IOB_X1Y140_I;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_A5 = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_A6 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D5 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_B1 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_B2 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_B3 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_B4 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_B5 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_B6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A2 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_C1 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_C2 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_C3 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_C4 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A3 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_C5 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_C6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A4 = CLBLM_R_X11Y126_SLICE_X15Y126_CQ;
  assign LIOB33_X0Y167_IOB_X0Y168_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOB33_X0Y167_IOB_X0Y167_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A5 = CLBLM_R_X7Y122_SLICE_X9Y122_AQ;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_D1 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_D2 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_D3 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_D4 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_D5 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X163Y140_D6 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_A1 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_A2 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_A3 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_A4 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_A5 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_A6 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_B1 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_B2 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_B3 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_B4 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_B5 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_B6 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_C1 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_C2 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_C3 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_C4 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_C5 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_C6 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_D1 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_D2 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_D3 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_D4 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_D5 = 1'b1;
  assign CLBLM_R_X103Y140_SLICE_X162Y140_D6 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_T1 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A3 = CLBLM_L_X10Y123_SLICE_X12Y123_AQ;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A4 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_A6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B1 = CLBLL_L_X4Y127_SLICE_X5Y127_DO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B2 = CLBLL_L_X4Y121_SLICE_X4Y121_BQ;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B4 = CLBLL_L_X2Y128_SLICE_X0Y128_AO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B5 = CLBLM_R_X3Y129_SLICE_X3Y129_AO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_B6 = CLBLM_R_X3Y127_SLICE_X3Y127_AO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C1 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C2 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C4 = CLBLL_L_X2Y130_SLICE_X0Y130_BO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C5 = CLBLL_L_X2Y130_SLICE_X0Y130_CO5;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_C6 = CLBLL_L_X2Y128_SLICE_X1Y128_AO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D1 = CLBLL_L_X2Y130_SLICE_X0Y130_CO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D2 = CLBLL_L_X2Y128_SLICE_X1Y128_AO5;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D3 = CLBLM_R_X3Y119_SLICE_X2Y119_AQ;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D4 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D5 = CLBLL_L_X2Y130_SLICE_X0Y130_AO6;
  assign CLBLM_R_X3Y127_SLICE_X3Y127_D6 = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A1 = CLBLL_L_X2Y130_SLICE_X0Y130_AO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A2 = CLBLL_L_X4Y125_SLICE_X5Y125_BQ;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A3 = CLBLL_L_X4Y130_SLICE_X4Y130_AO5;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A4 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A5 = CLBLL_L_X4Y120_SLICE_X4Y120_AQ;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_A6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B2 = CLBLL_L_X4Y125_SLICE_X5Y125_BQ;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B3 = CLBLM_R_X3Y129_SLICE_X3Y129_AO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B4 = CLBLL_L_X4Y129_SLICE_X4Y129_BO5;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B5 = CLBLL_L_X4Y120_SLICE_X4Y120_AQ;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_B6 = CLBLL_L_X2Y128_SLICE_X0Y128_AO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C1 = CLBLM_R_X3Y122_SLICE_X3Y122_BQ;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C2 = CLBLM_R_X3Y126_SLICE_X2Y126_CO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C3 = CLBLL_L_X4Y129_SLICE_X4Y129_BO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C4 = CLBLM_R_X3Y130_SLICE_X2Y130_BO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C5 = CLBLM_R_X3Y125_SLICE_X3Y125_BQ;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_C6 = CLBLL_L_X2Y127_SLICE_X1Y127_DO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D1 = CLBLM_R_X3Y127_SLICE_X2Y127_CO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D2 = CLBLL_L_X2Y129_SLICE_X1Y129_BO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D3 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D4 = CLBLL_L_X4Y125_SLICE_X5Y125_CO6;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D5 = 1'b1;
  assign CLBLM_R_X3Y127_SLICE_X2Y127_D6 = CLBLM_R_X3Y127_SLICE_X2Y127_BO6;
  assign LIOB33_X0Y169_IOB_X0Y170_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOB33_X0Y169_IOB_X0Y169_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_D1 = CLBLM_L_X10Y123_SLICE_X13Y123_DO5;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A4 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A5 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A6 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B1 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B2 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B3 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B4 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B5 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B6 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_A1 = CLBLL_L_X2Y130_SLICE_X0Y130_CO5;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_A2 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_A3 = CLBLL_L_X2Y130_SLICE_X0Y130_AO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_A4 = CLBLM_R_X3Y124_SLICE_X3Y124_BQ;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_A5 = CLBLL_L_X2Y130_SLICE_X0Y130_BO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_A6 = CLBLL_L_X2Y121_SLICE_X0Y121_BQ;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_B1 = CLBLM_R_X3Y125_SLICE_X3Y125_DO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_B2 = CLBLL_L_X4Y126_SLICE_X5Y126_CO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_B3 = CLBLM_R_X3Y127_SLICE_X3Y127_BO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_B4 = CLBLL_L_X2Y128_SLICE_X1Y128_DO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_B5 = CLBLL_L_X2Y129_SLICE_X1Y129_DO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_B6 = CLBLM_R_X3Y128_SLICE_X3Y128_CO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_C1 = CLBLL_L_X2Y126_SLICE_X0Y126_AO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_C2 = CLBLL_L_X2Y126_SLICE_X0Y126_CO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C2 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_C3 = CLBLL_L_X4Y129_SLICE_X4Y129_AQ;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_C4 = CLBLM_R_X3Y130_SLICE_X3Y130_CO6;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_C5 = CLBLL_L_X4Y120_SLICE_X4Y120_DQ;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_C6 = CLBLL_L_X4Y129_SLICE_X4Y129_BO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C3 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C4 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_D1 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_D2 = CLBLM_R_X3Y129_SLICE_X3Y129_AO5;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C5 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_D3 = CLBLM_R_X5Y128_SLICE_X6Y128_DQ;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_D4 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_D5 = CLBLL_L_X2Y126_SLICE_X0Y126_AO5;
  assign CLBLM_R_X3Y128_SLICE_X3Y128_D6 = CLBLL_L_X2Y130_SLICE_X0Y130_DO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C6 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_A1 = CLBLM_L_X8Y130_SLICE_X11Y130_DO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_A2 = CLBLL_L_X4Y126_SLICE_X5Y126_AO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_A3 = CLBLM_R_X3Y128_SLICE_X2Y128_BO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_A4 = CLBLL_L_X4Y128_SLICE_X5Y128_CO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_A5 = CLBLL_L_X2Y129_SLICE_X1Y129_CO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_A6 = CLBLM_R_X3Y128_SLICE_X2Y128_CO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_B1 = CLBLL_L_X2Y129_SLICE_X0Y129_CO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_B2 = CLBLL_L_X4Y124_SLICE_X4Y124_A5Q;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_B3 = CLBLL_L_X4Y129_SLICE_X5Y129_AQ;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_B4 = CLBLL_L_X2Y126_SLICE_X0Y126_AO5;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_B5 = CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_B6 = CLBLL_L_X2Y128_SLICE_X0Y128_DO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_C1 = CLBLL_L_X2Y126_SLICE_X0Y126_AO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_C2 = CLBLM_R_X5Y127_SLICE_X7Y127_CQ;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_C3 = CLBLL_L_X2Y129_SLICE_X0Y129_DO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_C4 = CLBLM_R_X3Y129_SLICE_X3Y129_AO5;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_C5 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_C6 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_D1 = CLBLL_L_X2Y128_SLICE_X0Y128_BO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_D3 = CLBLM_R_X3Y129_SLICE_X3Y129_DO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_D4 = CLBLL_L_X2Y130_SLICE_X1Y130_BO6;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_D5 = 1'b1;
  assign CLBLM_R_X3Y128_SLICE_X2Y128_D6 = CLBLM_R_X3Y119_SLICE_X2Y119_BQ;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_D1 = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_T1 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D5 = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_D1 = CLBLL_L_X2Y117_SLICE_X0Y117_CO5;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D6 = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_D1 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_D1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_T1 = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_D1 = CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1 = CLBLL_L_X4Y118_SLICE_X5Y118_CQ;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_D1 = LIOB33_X0Y75_IOB_X0Y76_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOB33_X0Y171_IOB_X0Y172_O = CLBLM_R_X103Y140_SLICE_X163Y140_AO6;
  assign LIOB33_X0Y171_IOB_X0Y171_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B5 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C1 = CLBLM_R_X5Y123_SLICE_X6Y123_AQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C2 = CLBLL_L_X4Y124_SLICE_X4Y124_AQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A1 = CLBLL_L_X2Y130_SLICE_X0Y130_CO5;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_A6 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B1 = CLBLL_L_X4Y124_SLICE_X4Y124_A5Q;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B2 = CLBLM_R_X7Y128_SLICE_X9Y128_BO5;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B3 = CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B4 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B5 = CLBLL_L_X2Y130_SLICE_X1Y130_AO5;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_B6 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C2 = CLBLL_L_X2Y130_SLICE_X0Y130_CO6;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C3 = CLBLL_L_X4Y129_SLICE_X5Y129_AQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_C6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C3 = CLBLL_L_X4Y123_SLICE_X4Y123_BQ;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D1 = CLBLL_L_X2Y128_SLICE_X1Y128_AO5;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D4 = CLBLM_R_X7Y129_SLICE_X8Y129_A5Q;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D5 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X3Y129_SLICE_X3Y129_D6 = CLBLL_L_X2Y130_SLICE_X0Y130_CO5;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C4 = CLBLL_L_X4Y122_SLICE_X4Y122_A5Q;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A1 = CLBLM_R_X3Y123_SLICE_X2Y123_CQ;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A2 = CLBLM_R_X3Y132_SLICE_X2Y132_CO5;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A3 = CLBLM_R_X3Y129_SLICE_X2Y129_AQ;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A4 = CLBLM_R_X3Y132_SLICE_X2Y132_A5Q;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A5 = CLBLL_L_X4Y129_SLICE_X4Y129_AQ;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B1 = CLBLM_L_X8Y130_SLICE_X11Y130_DO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B2 = CLBLM_R_X3Y129_SLICE_X3Y129_BO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B3 = CLBLM_R_X3Y129_SLICE_X3Y129_CO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B4 = CLBLL_L_X2Y128_SLICE_X1Y128_CO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B5 = CLBLL_L_X2Y128_SLICE_X0Y128_DO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_B6 = CLBLL_L_X2Y129_SLICE_X0Y129_DO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C1 = CLBLL_L_X4Y128_SLICE_X5Y128_CO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C2 = CLBLL_L_X2Y129_SLICE_X1Y129_CO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C3 = CLBLL_L_X4Y126_SLICE_X5Y126_AO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C4 = CLBLL_L_X4Y130_SLICE_X4Y130_CO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C5 = CLBLM_R_X3Y129_SLICE_X2Y129_DO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_C6 = CLBLM_R_X3Y129_SLICE_X2Y129_BO6;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C5 = CLBLL_L_X4Y123_SLICE_X5Y123_DO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D1 = CLBLL_L_X2Y128_SLICE_X0Y128_CO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D2 = 1'b1;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D3 = CLBLM_R_X3Y130_SLICE_X2Y130_BO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D4 = CLBLM_R_X3Y130_SLICE_X3Y130_AO5;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D5 = CLBLL_L_X2Y130_SLICE_X1Y130_CO6;
  assign CLBLM_R_X3Y129_SLICE_X2Y129_D6 = CLBLL_L_X2Y129_SLICE_X0Y129_CO6;
  assign LIOB33_X0Y173_IOB_X0Y174_O = CLBLM_R_X11Y151_SLICE_X14Y151_AO6;
  assign LIOB33_X0Y173_IOB_X0Y173_O = CLBLM_R_X103Y140_SLICE_X163Y140_AO5;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_T1 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A2 = CLBLL_L_X2Y130_SLICE_X0Y130_CO5;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A6 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B1 = CLBLM_R_X3Y130_SLICE_X3Y130_DO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B2 = CLBLM_R_X3Y130_SLICE_X2Y130_DO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B3 = CLBLL_L_X4Y129_SLICE_X4Y129_DO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B4 = CLBLM_R_X3Y130_SLICE_X2Y130_CO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B5 = CLBLM_R_X7Y129_SLICE_X8Y129_DQ;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B6 = CLBLL_L_X4Y126_SLICE_X4Y126_BO6;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_D = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C3 = CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C6 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C4 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C5 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D1 = CLBLM_R_X3Y130_SLICE_X3Y130_AO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D2 = CLBLL_L_X2Y130_SLICE_X1Y130_BO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D3 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D4 = CLBLL_L_X4Y130_SLICE_X4Y130_DO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D5 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D6 = CLBLM_R_X3Y123_SLICE_X2Y123_AQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C6 = 1'b1;
  assign LIOB33_X0Y109_IOB_X0Y110_O = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_D = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOB33_X0Y109_IOB_X0Y109_O = CLBLL_L_X2Y118_SLICE_X1Y118_CO5;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A1 = CLBLL_L_X4Y124_SLICE_X4Y124_CQ;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A2 = CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A4 = CLBLM_R_X3Y131_SLICE_X2Y131_BQ;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A5 = CLBLM_R_X3Y131_SLICE_X2Y131_CO5;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A6 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B4 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B6 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C3 = CLBLL_L_X2Y130_SLICE_X0Y130_CO5;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C6 = CLBLL_L_X2Y129_SLICE_X0Y129_CO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D2 = CLBLL_L_X2Y128_SLICE_X0Y128_BO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D3 = CLBLL_L_X2Y130_SLICE_X1Y130_CO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D5 = CLBLM_R_X3Y130_SLICE_X2Y130_BO5;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D6 = CLBLM_R_X3Y130_SLICE_X2Y130_BO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D5 = 1'b1;
  assign LIOB33_X0Y175_IOB_X0Y176_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign LIOB33_X0Y175_IOB_X0Y175_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D6 = 1'b1;
  assign RIOB33_X105Y191_IOB_X1Y192_O = CLBLM_L_X12Y121_SLICE_X16Y121_BQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_D1 = CLBLM_R_X3Y123_SLICE_X2Y123_CQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B5 = CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_D1 = CLBLM_R_X103Y140_SLICE_X163Y140_AO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_T1 = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_D = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_BX = CLBLM_L_X10Y124_SLICE_X12Y124_BO6;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_T1 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_D1 = CLBLL_L_X2Y115_SLICE_X0Y115_AO6;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_D1 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B6 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_T1 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_D1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C4 = CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_T1 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C5 = CLBLM_L_X10Y124_SLICE_X12Y124_CO5;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_D1 = CLBLL_L_X2Y118_SLICE_X1Y118_CO5;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = CLBLM_R_X3Y131_SLICE_X2Y131_BQ;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_T1 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_D1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1 = CLBLL_L_X2Y117_SLICE_X0Y117_BO5;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_D1 = CLBLM_R_X3Y132_SLICE_X2Y132_A5Q;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_T1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C4 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = CLBLM_R_X3Y131_SLICE_X2Y131_AQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C5 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A2 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A3 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A4 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A6 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B2 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B3 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B4 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C2 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C3 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C4 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C6 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_T1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D2 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D3 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D4 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D6 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A3 = CLBLM_R_X3Y131_SLICE_X2Y131_AQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A4 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A5 = CLBLL_L_X2Y118_SLICE_X1Y118_AQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A6 = CLBLM_R_X3Y131_SLICE_X2Y131_CO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B2 = CLBLM_R_X3Y131_SLICE_X2Y131_BQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B3 = CLBLL_L_X2Y118_SLICE_X1Y118_AQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B5 = CLBLM_R_X3Y131_SLICE_X2Y131_CO5;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B6 = CLBLM_R_X7Y125_SLICE_X9Y125_A5Q;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C1 = CLBLM_R_X3Y129_SLICE_X2Y129_AQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C2 = CLBLM_R_X3Y131_SLICE_X2Y131_AQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C3 = CLBLM_R_X3Y132_SLICE_X2Y132_BQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C4 = CLBLM_R_X3Y132_SLICE_X2Y132_A5Q;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C5 = CLBLM_R_X3Y123_SLICE_X2Y123_CQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C6 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y177_IOB_X0Y178_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOB33_X0Y177_IOB_X0Y177_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D2 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D3 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D4 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D6 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A1 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A2 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A3 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A4 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A5 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_A6 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B1 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C4 = CLBLM_L_X8Y126_SLICE_X11Y126_BQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B2 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B3 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B4 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B5 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C5 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_B6 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C1 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C6 = CLBLM_L_X8Y124_SLICE_X11Y124_BQ;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C2 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C3 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C4 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C5 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_C6 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D1 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D2 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D3 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D4 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D5 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X17Y126_D6 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A1 = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A3 = CLBLM_L_X12Y126_SLICE_X16Y126_AQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A4 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A5 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_A6 = 1'b1;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_D = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B1 = CLBLM_L_X12Y126_SLICE_X16Y126_BQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B2 = CLBLM_R_X7Y127_SLICE_X8Y127_BQ;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B4 = CLBLM_L_X12Y127_SLICE_X16Y127_BO6;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B5 = CLBLM_R_X11Y130_SLICE_X14Y130_BO5;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_B6 = CLBLM_R_X11Y127_SLICE_X15Y127_BO5;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C1 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C2 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C3 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C4 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C5 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_C6 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D1 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D2 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D3 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D4 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D5 = 1'b1;
  assign CLBLM_L_X12Y126_SLICE_X16Y126_D6 = 1'b1;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_D = RIOB33_X105Y111_IOB_X1Y112_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1 = 1'b1;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_D = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D1 = CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D2 = 1'b1;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_D = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_D1 = LIOB33_X0Y69_IOB_X0Y69_I;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A1 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A2 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A3 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A4 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A5 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A6 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B1 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B2 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B3 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B4 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B5 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B6 = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_T1 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C1 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C2 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C3 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C4 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C5 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C6 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D1 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D2 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D3 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D4 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D5 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D6 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A1 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A3 = CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A5 = CLBLL_L_X2Y118_SLICE_X1Y118_AQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A6 = CLBLL_L_X2Y132_SLICE_X1Y132_AO6;
  assign LIOB33_X0Y179_IOB_X0Y179_O = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOB33_X0Y179_IOB_X0Y180_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_AX = CLBLM_R_X3Y132_SLICE_X2Y132_CO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B1 = CLBLM_R_X3Y132_SLICE_X2Y132_DO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B2 = CLBLM_R_X3Y132_SLICE_X2Y132_BQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B3 = CLBLL_L_X2Y118_SLICE_X1Y118_AQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B6 = CLBLM_R_X5Y129_SLICE_X6Y129_BQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C2 = CLBLL_L_X2Y118_SLICE_X1Y118_AQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C3 = CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C4 = CLBLM_R_X3Y132_SLICE_X2Y132_A5Q;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C6 = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_D1 = LIOB33_X0Y63_IOB_X0Y64_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D1 = CLBLM_R_X3Y123_SLICE_X2Y123_CQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D2 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D3 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D4 = CLBLM_R_X3Y132_SLICE_X2Y132_A5Q;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D5 = CLBLM_R_X3Y129_SLICE_X2Y129_AQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D6 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A1 = CLBLM_L_X12Y127_SLICE_X17Y127_DO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A2 = CLBLM_R_X11Y128_SLICE_X14Y128_AO5;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A3 = CLBLM_R_X11Y126_SLICE_X15Y126_CQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A4 = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A5 = CLBLM_L_X10Y129_SLICE_X13Y129_CO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_A6 = CLBLM_L_X12Y127_SLICE_X17Y127_CO6;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B1 = CLBLM_R_X11Y126_SLICE_X15Y126_AQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B2 = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B3 = CLBLM_L_X12Y126_SLICE_X16Y126_BQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B4 = CLBLM_L_X10Y128_SLICE_X13Y128_AQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B5 = CLBLM_R_X11Y128_SLICE_X14Y128_DO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_B6 = CLBLM_R_X11Y126_SLICE_X14Y126_CQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C1 = CLBLM_L_X12Y126_SLICE_X16Y126_BQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C2 = CLBLM_R_X11Y126_SLICE_X14Y126_CQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C3 = CLBLM_R_X11Y126_SLICE_X15Y126_AQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A4 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A5 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A6 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C4 = CLBLM_R_X11Y128_SLICE_X14Y128_DO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C5 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_C6 = CLBLM_L_X10Y128_SLICE_X13Y128_AQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B1 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B2 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B3 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B4 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B5 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_B6 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D1 = CLBLM_R_X11Y128_SLICE_X15Y128_DO6;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D2 = CLBLM_R_X11Y126_SLICE_X14Y126_CQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D3 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D4 = CLBLM_L_X12Y126_SLICE_X16Y126_BQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D5 = CLBLM_R_X11Y126_SLICE_X15Y126_AQ;
  assign CLBLM_L_X12Y127_SLICE_X17Y127_D6 = CLBLM_L_X10Y128_SLICE_X13Y128_AQ;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C2 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C3 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C5 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A1 = CLBLM_L_X12Y127_SLICE_X16Y127_DO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A2 = CLBLM_R_X5Y116_SLICE_X7Y116_BQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A4 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A5 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_A6 = CLBLM_R_X11Y127_SLICE_X15Y127_BO5;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D1 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D2 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D3 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D4 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D5 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_D6 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B1 = CLBLM_R_X11Y128_SLICE_X14Y128_AO5;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B2 = CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B3 = CLBLM_R_X11Y128_SLICE_X15Y128_DO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B4 = CLBLM_L_X10Y128_SLICE_X13Y128_AQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B5 = CLBLM_L_X10Y129_SLICE_X13Y129_CO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_B6 = CLBLM_R_X11Y128_SLICE_X14Y128_DO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C1 = CLBLM_L_X12Y126_SLICE_X16Y126_BQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C2 = CLBLM_R_X11Y126_SLICE_X15Y126_AQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C3 = CLBLM_R_X13Y127_SLICE_X18Y127_AQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A6 = CLBLM_L_X8Y117_SLICE_X10Y117_CO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C4 = CLBLM_R_X11Y126_SLICE_X14Y126_CQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C5 = CLBLM_R_X11Y128_SLICE_X15Y128_DO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_C6 = CLBLM_L_X10Y128_SLICE_X13Y128_AQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A2 = CLBLM_L_X12Y126_SLICE_X16Y126_BQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B2 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B3 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B4 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B5 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B6 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D1 = CLBLM_L_X10Y129_SLICE_X13Y129_CO6;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D2 = CLBLM_L_X12Y127_SLICE_X16Y127_AQ;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D3 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D4 = CLBLM_R_X11Y128_SLICE_X14Y128_AO5;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D5 = CLBLM_R_X11Y130_SLICE_X14Y130_BO5;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C2 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C3 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C4 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C5 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C6 = 1'b1;
  assign CLBLM_L_X12Y127_SLICE_X16Y127_D6 = CLBLM_L_X10Y128_SLICE_X12Y128_BQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_C1 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D1 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D2 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D3 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D4 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D5 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_D6 = 1'b1;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1 = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A1 = CLBLM_L_X8Y117_SLICE_X11Y117_BO6;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C4 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A5 = CLBLM_L_X8Y116_SLICE_X10Y116_DO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A6 = CLBLM_L_X8Y116_SLICE_X11Y116_CO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D5 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B1 = CLBLM_R_X7Y118_SLICE_X9Y118_BO5;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B2 = CLBLM_R_X5Y118_SLICE_X7Y118_BO5;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B5 = CLBLM_R_X7Y119_SLICE_X8Y119_CQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C3 = CLBLM_R_X7Y118_SLICE_X9Y118_BO5;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_D1 = CLBLM_R_X11Y151_SLICE_X14Y151_AO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C4 = CLBLM_R_X7Y115_SLICE_X9Y115_AO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C5 = CLBLM_R_X3Y124_SLICE_X3Y124_DO6;
  assign LIOB33_X0Y181_IOB_X0Y182_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOB33_X0Y181_IOB_X0Y181_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_T1 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_D1 = CLBLM_L_X10Y121_SLICE_X13Y121_B5Q;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_D1 = CLBLM_R_X103Y140_SLICE_X163Y140_AO5;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_T1 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_D1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_T1 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_D1 = 1'b0;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_T1 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_D1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A2 = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A3 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A4 = CLBLM_L_X10Y118_SLICE_X13Y118_BO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A5 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_A6 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B1 = CLBLM_L_X10Y120_SLICE_X13Y120_A5Q;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B2 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B3 = CLBLM_L_X10Y118_SLICE_X13Y118_AQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B4 = CLBLM_L_X8Y117_SLICE_X11Y117_AO6;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B5 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_B6 = CLBLM_R_X5Y119_SLICE_X6Y119_CQ;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C1 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C2 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C3 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C4 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C5 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_C6 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D1 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D2 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D3 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D4 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D5 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X13Y118_D6 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A1 = CLBLM_L_X10Y128_SLICE_X12Y128_DQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A3 = CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A4 = CLBLM_L_X10Y118_SLICE_X12Y118_BO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A5 = CLBLM_L_X8Y116_SLICE_X11Y116_AO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_A6 = CLBLM_R_X7Y118_SLICE_X9Y118_BO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A6 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C6 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B1 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B2 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B3 = CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B4 = CLBLM_R_X7Y118_SLICE_X9Y118_BO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B5 = CLBLM_L_X8Y118_SLICE_X11Y118_CO5;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_B6 = CLBLM_L_X10Y121_SLICE_X12Y121_CQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C1 = CLBLM_L_X8Y118_SLICE_X11Y118_CO5;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C2 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C3 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C4 = CLBLM_L_X10Y121_SLICE_X12Y121_CQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C5 = CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_C6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B1 = CLBLM_R_X3Y123_SLICE_X2Y123_DQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B2 = CLBLM_L_X8Y116_SLICE_X10Y116_BQ;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D1 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D2 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D3 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D4 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D5 = 1'b1;
  assign CLBLM_L_X10Y118_SLICE_X12Y118_D6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B3 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_D = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_D = LIOB33_X0Y51_IOB_X0Y51_I;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1 = CLBLM_R_X11Y131_SLICE_X15Y131_AQ;
  assign RIOB33_X105Y151_IOB_X1Y152_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOB33_X105Y151_IOB_X1Y151_O = LIOB33_X0Y75_IOB_X0Y76_I;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOB33_X0Y183_IOB_X0Y184_O = RIOB33_X105Y135_IOB_X1Y136_I;
  assign LIOB33_X0Y183_IOB_X0Y183_O = RIOB33_X105Y135_IOB_X1Y135_I;
  assign RIOB33_SING_X105Y150_IOB_X1Y150_O = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C4 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C5 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C6 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A6 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_AX = CLBLL_L_X4Y122_SLICE_X4Y122_CO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B3 = CLBLL_L_X4Y122_SLICE_X5Y122_C5Q;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B4 = CLBLM_R_X5Y122_SLICE_X7Y122_BQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D1 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B6 = CLBLM_R_X5Y122_SLICE_X7Y122_CO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D2 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D3 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D4 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A1 = CLBLM_L_X10Y120_SLICE_X13Y120_BQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D5 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A3 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A5 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A6 = CLBLM_L_X8Y119_SLICE_X11Y119_CQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_A2 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B1 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B2 = CLBLM_L_X10Y119_SLICE_X13Y119_BQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B3 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B4 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_B6 = CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C3 = CLBLM_R_X5Y123_SLICE_X6Y123_AQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C1 = CLBLM_L_X8Y117_SLICE_X11Y117_AO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C2 = CLBLM_L_X10Y124_SLICE_X13Y124_D5Q;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C4 = CLBLM_L_X10Y123_SLICE_X13Y123_BQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C5 = CLBLM_L_X10Y119_SLICE_X12Y119_DQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C3 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_C6 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C4 = CLBLL_L_X4Y122_SLICE_X4Y122_A5Q;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C5 = CLBLM_R_X5Y124_SLICE_X6Y124_DO5;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C6 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D1 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D2 = CLBLM_L_X10Y120_SLICE_X13Y120_CQ;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D3 = CLBLM_L_X10Y120_SLICE_X13Y120_DO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D4 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D5 = CLBLM_L_X8Y119_SLICE_X10Y119_DO6;
  assign CLBLM_L_X10Y119_SLICE_X13Y119_D6 = CLBLM_L_X10Y121_SLICE_X13Y121_AQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A1 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A2 = CLBLM_L_X10Y118_SLICE_X12Y118_CO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A3 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A4 = CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A5 = CLBLM_L_X8Y116_SLICE_X11Y116_AO6;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_A6 = CLBLM_L_X10Y121_SLICE_X12Y121_CQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A2 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A3 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B3 = CLBLM_R_X3Y118_SLICE_X3Y118_BQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A4 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B4 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B5 = CLBLM_L_X10Y122_SLICE_X12Y122_AQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_B6 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A5 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C2 = CLBLM_L_X10Y119_SLICE_X12Y119_CQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C3 = CLBLM_R_X11Y122_SLICE_X14Y122_DQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C4 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C5 = CLBLM_R_X5Y119_SLICE_X6Y119_CQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_C6 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A6 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D1 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D2 = CLBLM_L_X10Y119_SLICE_X12Y119_CQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D3 = CLBLM_L_X10Y119_SLICE_X12Y119_DQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D4 = 1'b1;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D5 = CLBLM_L_X8Y127_SLICE_X10Y127_CQ;
  assign CLBLM_L_X10Y119_SLICE_X12Y119_D6 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_AX = CLBLM_L_X10Y136_SLICE_X12Y136_BO5;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D2 = CLBLM_L_X10Y121_SLICE_X12Y121_DQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D3 = CLBLM_R_X3Y123_SLICE_X2Y123_AQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D4 = 1'b1;
  assign LIOB33_X0Y111_IOB_X0Y111_O = 1'b0;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B1 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B2 = 1'b1;
  assign RIOB33_X105Y153_IOB_X1Y154_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOB33_X105Y153_IOB_X1Y153_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B3 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B4 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B5 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B6 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_BX = CLBLM_L_X10Y136_SLICE_X12Y136_AO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C1 = 1'b1;
  assign LIOB33_X0Y185_IOB_X0Y186_O = RIOB33_X105Y143_IOB_X1Y143_I;
  assign LIOB33_X0Y185_IOB_X0Y185_O = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C2 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C3 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C4 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C5 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D = RIOB33_X105Y119_IOB_X1Y119_I;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = CLBLL_L_X4Y122_SLICE_X5Y122_C5Q;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D1 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C4 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D2 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C5 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D3 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C6 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D5 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D2 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = CLBLL_L_X4Y118_SLICE_X5Y118_C5Q;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A1 = CLBLM_R_X7Y125_SLICE_X9Y125_B5Q;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A2 = CLBLM_L_X10Y121_SLICE_X13Y121_AQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A4 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_A6 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B3 = CLBLL_L_X4Y123_SLICE_X5Y123_AQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D5 = 1'b1;
  assign RIOB33_X105Y187_IOB_X1Y187_O = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B1 = CLBLM_L_X10Y121_SLICE_X12Y121_BQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B2 = CLBLM_L_X10Y120_SLICE_X13Y120_BQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B3 = CLBLM_L_X10Y119_SLICE_X13Y119_BQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B4 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_B6 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B4 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D6 = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_D1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C1 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C2 = CLBLM_L_X10Y121_SLICE_X13Y121_AQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C3 = CLBLM_R_X7Y125_SLICE_X9Y125_B5Q;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C4 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C5 = CLBLM_L_X10Y120_SLICE_X13Y120_CQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B6 = CLBLL_L_X4Y123_SLICE_X5Y123_CO5;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_D1 = CLBLM_R_X5Y128_SLICE_X7Y128_BQ;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_T1 = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_D1 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D1 = CLBLM_L_X10Y122_SLICE_X13Y122_AQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D2 = CLBLM_R_X5Y119_SLICE_X6Y119_CQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D3 = CLBLM_R_X7Y118_SLICE_X8Y118_DQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D4 = CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D5 = CLBLM_L_X10Y120_SLICE_X13Y120_BO5;
  assign CLBLM_L_X10Y120_SLICE_X13Y120_D6 = CLBLM_L_X10Y124_SLICE_X13Y124_AQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_T1 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_D1 = CLBLM_R_X11Y124_SLICE_X14Y124_DO5;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_T1 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A1 = CLBLM_L_X10Y120_SLICE_X12Y120_DO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A3 = CLBLM_R_X7Y118_SLICE_X9Y118_BO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A5 = CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_A6 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C2 = CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_D1 = CLBLM_L_X10Y121_SLICE_X13Y121_BQ;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1 = RIOB33_X105Y145_IOB_X1Y145_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B2 = CLBLM_L_X10Y120_SLICE_X12Y120_BQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B4 = CLBLM_R_X7Y120_SLICE_X9Y120_AO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B5 = CLBLM_L_X10Y119_SLICE_X13Y119_BQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_B6 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_T1 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C2 = CLBLM_L_X10Y120_SLICE_X12Y120_CQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C3 = CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C4 = CLBLM_L_X10Y121_SLICE_X12Y121_BQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_C6 = CLBLM_L_X8Y128_SLICE_X10Y128_BQ;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A6 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_T1 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y193_IOB_X0Y194_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign RIOB33_X105Y155_IOB_X1Y155_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign RIOB33_X105Y155_IOB_X1Y156_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D1 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D2 = CLBLM_L_X10Y120_SLICE_X12Y120_AQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D3 = 1'b1;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D4 = CLBLM_L_X8Y120_SLICE_X10Y120_CO6;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D5 = CLBLM_R_X11Y123_SLICE_X14Y123_AQ;
  assign CLBLM_L_X10Y120_SLICE_X12Y120_D6 = CLBLM_L_X8Y120_SLICE_X11Y120_BO6;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1 = 1'b1;
  assign LIOB33_X0Y193_IOB_X0Y193_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B3 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B4 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B5 = 1'b1;
  assign LIOB33_X0Y187_IOB_X0Y188_O = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOB33_X0Y187_IOB_X0Y187_O = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C2 = CLBLM_L_X10Y125_SLICE_X13Y125_CQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A1 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C2 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A4 = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A5 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A6 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C6 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D1 = CLBLM_L_X8Y126_SLICE_X11Y126_CQ;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B2 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D5 = CLBLM_L_X10Y124_SLICE_X13Y124_C5Q;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B4 = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_D = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B6 = 1'b1;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_D = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D2 = 1'b1;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_D = LIOB33_X0Y53_IOB_X0Y53_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_D = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D3 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D4 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D5 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B4 = CLBLM_L_X8Y118_SLICE_X11Y118_BQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B5 = CLBLM_L_X8Y128_SLICE_X11Y128_AQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B6 = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_D = LIOB33_X0Y69_IOB_X0Y69_I;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_D1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A1 = CLBLM_L_X8Y125_SLICE_X10Y125_CQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C4 = CLBLM_L_X8Y127_SLICE_X11Y127_BQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A2 = CLBLM_L_X10Y124_SLICE_X13Y124_AQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A3 = CLBLM_L_X10Y121_SLICE_X13Y121_AQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A5 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C5 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_A6 = CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B2 = CLBLM_L_X8Y122_SLICE_X11Y122_A5Q;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B3 = CLBLM_R_X7Y117_SLICE_X8Y117_DQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B6 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_B5 = CLBLM_R_X11Y123_SLICE_X14Y123_BQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C2 = CLBLM_L_X10Y121_SLICE_X13Y121_CQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C3 = CLBLM_R_X5Y120_SLICE_X7Y120_DO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C4 = CLBLL_L_X4Y119_SLICE_X4Y119_CQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_C6 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A1 = CLBLL_L_X4Y122_SLICE_X4Y122_BQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A3 = CLBLL_L_X4Y117_SLICE_X5Y117_CO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A4 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_A6 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D1 = CLBLM_R_X11Y123_SLICE_X14Y123_AQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D2 = CLBLM_L_X8Y120_SLICE_X10Y120_DO6;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B2 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B3 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B4 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B5 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_B6 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D4 = CLBLM_R_X11Y122_SLICE_X15Y122_BQ;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D5 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C2 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C3 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C4 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C5 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_C6 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A1 = CLBLM_L_X8Y121_SLICE_X11Y121_DO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A2 = CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A6 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B1 = CLBLL_L_X4Y121_SLICE_X4Y121_DQ;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D2 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D3 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D4 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D5 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X4Y117_D6 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C5 = CLBLM_R_X11Y127_SLICE_X14Y127_AQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C6 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C1 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C3 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_C4 = CLBLM_L_X10Y126_SLICE_X12Y126_A5Q;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D1 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D2 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D4 = CLBLL_L_X4Y123_SLICE_X5Y123_BQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D5 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOB33_X0Y189_IOB_X0Y190_O = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOB33_X0Y189_IOB_X0Y189_O = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A2 = CLBLM_R_X5Y117_SLICE_X6Y117_AQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A3 = CLBLL_L_X4Y117_SLICE_X5Y117_AQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A5 = CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_A6 = CLBLL_L_X4Y118_SLICE_X5Y118_CQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B1 = CLBLL_L_X4Y119_SLICE_X5Y119_DO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B2 = CLBLL_L_X4Y117_SLICE_X5Y117_BQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B3 = CLBLM_R_X3Y124_SLICE_X2Y124_DQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B5 = CLBLM_R_X5Y116_SLICE_X7Y116_DO5;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_B6 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_D1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign RIOB33_X105Y175_IOB_X1Y176_O = CLBLM_R_X103Y173_SLICE_X163Y173_AO5;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C1 = CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C2 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C4 = CLBLM_R_X3Y123_SLICE_X2Y123_DQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C5 = CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_C6 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D1 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D2 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D3 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D4 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D5 = 1'b1;
  assign CLBLL_L_X4Y117_SLICE_X5Y117_D6 = 1'b1;
  assign RIOB33_X105Y175_IOB_X1Y175_O = CLBLM_L_X10Y136_SLICE_X12Y136_BO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D3 = CLBLM_L_X10Y125_SLICE_X12Y125_DQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D4 = CLBLM_L_X10Y124_SLICE_X13Y124_AQ;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_T1 = 1'b1;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_D = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A6 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_D1 = CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B3 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1 = CLBLM_R_X11Y124_SLICE_X14Y124_DO5;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B6 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_T1 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A1 = CLBLM_L_X10Y128_SLICE_X12Y128_CQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A2 = CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A3 = CLBLM_L_X10Y122_SLICE_X13Y122_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A4 = CLBLM_L_X10Y120_SLICE_X13Y120_BQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_A6 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D2 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B1 = CLBLM_R_X7Y121_SLICE_X9Y121_B5Q;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B2 = CLBLM_L_X10Y119_SLICE_X12Y119_DQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D3 = CLBLL_L_X4Y125_SLICE_X4Y125_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B4 = CLBLM_L_X10Y121_SLICE_X13Y121_CQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_B6 = 1'b1;
  assign RIOB33_X105Y159_IOB_X1Y160_O = CLBLM_R_X11Y124_SLICE_X14Y124_DO5;
  assign RIOB33_X105Y159_IOB_X1Y159_O = CLBLM_R_X11Y124_SLICE_X14Y124_DO6;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C2 = CLBLL_L_X4Y122_SLICE_X4Y122_DQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C4 = CLBLM_L_X10Y123_SLICE_X13Y123_BQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C5 = CLBLM_L_X10Y122_SLICE_X12Y122_BQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_C6 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A2 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A3 = CLBLL_L_X4Y118_SLICE_X4Y118_AQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A5 = CLBLM_L_X10Y118_SLICE_X13Y118_AQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_A6 = CLBLL_L_X2Y118_SLICE_X1Y118_A5Q;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D2 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D3 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D4 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D5 = CLBLM_R_X7Y121_SLICE_X9Y121_B5Q;
  assign CLBLM_L_X10Y122_SLICE_X13Y122_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B1 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B2 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B3 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B4 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B5 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_B6 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A1 = CLBLM_L_X10Y123_SLICE_X12Y123_CQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A2 = CLBLM_L_X8Y123_SLICE_X11Y123_C5Q;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A3 = CLBLM_L_X10Y122_SLICE_X12Y122_AQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_A6 = CLBLM_L_X10Y122_SLICE_X12Y122_CO6;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C1 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C2 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C3 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C4 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B1 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B4 = CLBLM_L_X10Y124_SLICE_X13Y124_D5Q;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B5 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_B6 = CLBLM_L_X10Y123_SLICE_X12Y123_CQ;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D1 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D2 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D3 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D4 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D5 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_D6 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C1 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C5 = CLBLM_L_X10Y126_SLICE_X13Y126_DQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C6 = CLBLM_L_X8Y122_SLICE_X10Y122_BO6;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C2 = CLBLM_L_X10Y122_SLICE_X12Y122_AQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C3 = CLBLM_L_X10Y122_SLICE_X12Y122_BQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_C4 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D1 = CLBLL_L_X4Y122_SLICE_X5Y122_DQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D2 = CLBLM_L_X10Y123_SLICE_X12Y123_CQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D3 = CLBLM_R_X11Y123_SLICE_X14Y123_DQ;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D4 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D5 = 1'b1;
  assign CLBLM_L_X10Y122_SLICE_X12Y122_D6 = CLBLM_R_X5Y124_SLICE_X6Y124_CQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A1 = CLBLL_L_X4Y120_SLICE_X5Y120_CQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A3 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A4 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A5 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B1 = CLBLM_R_X3Y119_SLICE_X3Y119_BO5;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B2 = CLBLL_L_X4Y118_SLICE_X5Y118_BQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B3 = CLBLM_R_X5Y130_SLICE_X7Y130_AQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B4 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B5 = CLBLM_R_X5Y118_SLICE_X6Y118_CO5;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A1 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A2 = CLBLL_L_X4Y117_SLICE_X5Y117_BQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C2 = CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C3 = CLBLM_R_X5Y118_SLICE_X6Y118_DQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C4 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_C6 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A3 = CLBLM_R_X5Y116_SLICE_X7Y116_CQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_D1 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A5 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D1 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D2 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D3 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D4 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D5 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X5Y118_D6 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A6 = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_T1 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_D1 = CLBLL_L_X4Y122_SLICE_X5Y122_CQ;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_D1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_T1 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_D1 = CLBLM_L_X10Y126_SLICE_X12Y126_DO5;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B1 = CLBLM_R_X3Y124_SLICE_X3Y124_DO6;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_T1 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B2 = CLBLM_L_X8Y117_SLICE_X10Y117_DO5;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_D1 = CLBLL_L_X2Y122_SLICE_X1Y122_AQ;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B3 = CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_T1 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B4 = CLBLM_L_X10Y124_SLICE_X13Y124_D5Q;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B5 = CLBLM_R_X3Y126_SLICE_X2Y126_BO6;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_T1 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_D1 = CLBLM_L_X10Y126_SLICE_X12Y126_DO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_B6 = CLBLM_L_X8Y117_SLICE_X11Y117_AO5;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_T1 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C3 = CLBLM_R_X7Y118_SLICE_X8Y118_C5Q;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1 = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOB33_X105Y161_IOB_X1Y162_O = CLBLM_L_X10Y126_SLICE_X12Y126_DO5;
  assign RIOB33_X105Y161_IOB_X1Y161_O = CLBLM_L_X10Y126_SLICE_X12Y126_DO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A1 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A3 = CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A4 = CLBLM_L_X10Y121_SLICE_X13Y121_CQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_A6 = CLBLM_L_X10Y126_SLICE_X13Y126_CQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C3 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B1 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B2 = CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B3 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B4 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_B6 = CLBLM_L_X10Y119_SLICE_X13Y119_CO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A2 = CLBLM_R_X5Y126_SLICE_X7Y126_CO5;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C4 = CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_C6 = CLBLM_R_X11Y126_SLICE_X14Y126_BQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A3 = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A4 = CLBLM_R_X3Y120_SLICE_X3Y120_BQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A5 = CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_A6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B1 = CLBLM_L_X8Y123_SLICE_X11Y123_CQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B2 = CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B3 = CLBLM_R_X3Y119_SLICE_X3Y119_BO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D1 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D2 = CLBLM_L_X10Y123_SLICE_X13Y123_CQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D3 = CLBLL_L_X4Y121_SLICE_X5Y121_CQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D4 = CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D5 = CLBLL_L_X4Y117_SLICE_X4Y117_AQ;
  assign CLBLM_L_X10Y123_SLICE_X13Y123_D6 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B5 = CLBLM_L_X10Y120_SLICE_X12Y120_BQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C1 = CLBLL_L_X4Y122_SLICE_X4Y122_AQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C2 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A1 = CLBLM_L_X8Y127_SLICE_X10Y127_CQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A2 = CLBLM_R_X11Y121_SLICE_X14Y121_CQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A3 = CLBLM_L_X10Y123_SLICE_X12Y123_AQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A5 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_A6 = CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_C6 = CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B1 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B2 = CLBLM_L_X10Y123_SLICE_X12Y123_BQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D1 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D2 = CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D3 = CLBLL_L_X4Y119_SLICE_X4Y119_DQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D4 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y119_SLICE_X4Y119_D6 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B4 = CLBLM_R_X7Y123_SLICE_X9Y123_DO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_B6 = CLBLM_L_X10Y123_SLICE_X13Y123_CQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C4 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C5 = 1'b1;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C6 = CLBLM_L_X10Y119_SLICE_X12Y119_BQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C1 = CLBLM_R_X7Y119_SLICE_X9Y119_BQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B5 = CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_AX = CLBLM_L_X10Y126_SLICE_X12Y126_BO6;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D1 = CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D4 = CLBLM_L_X10Y122_SLICE_X13Y122_CQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D5 = CLBLM_R_X3Y125_SLICE_X2Y125_AQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A1 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A2 = CLBLL_L_X4Y117_SLICE_X5Y117_BQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A3 = CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A5 = CLBLM_R_X5Y126_SLICE_X7Y126_CO5;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_A6 = CLBLL_L_X4Y119_SLICE_X4Y119_CQ;
  assign CLBLM_L_X10Y123_SLICE_X12Y123_D6 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B2 = CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B1 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B2 = CLBLL_L_X4Y119_SLICE_X5Y119_BQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B3 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B4 = CLBLM_R_X3Y121_SLICE_X2Y121_C5Q;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_B6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B3 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B5 = 1'b1;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C1 = CLBLL_L_X4Y128_SLICE_X4Y128_AO6;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C2 = CLBLL_L_X4Y119_SLICE_X5Y119_CQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C4 = CLBLL_L_X4Y117_SLICE_X4Y117_AO5;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C5 = CLBLM_R_X7Y119_SLICE_X8Y119_DQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_B6 = CLBLL_L_X4Y117_SLICE_X5Y117_AQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D2 = CLBLM_R_X5Y120_SLICE_X6Y120_BQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D4 = CLBLM_R_X7Y126_SLICE_X9Y126_BQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D5 = CLBLM_R_X3Y119_SLICE_X3Y119_AQ;
  assign CLBLL_L_X4Y119_SLICE_X5Y119_D6 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A1 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A2 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A3 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A4 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A5 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_A6 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B1 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B2 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B3 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B4 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B5 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_B6 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C1 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C2 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C3 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C4 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C5 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_C6 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D1 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D2 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D3 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D4 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D5 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X19Y127_D6 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A1 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A2 = CLBLM_R_X11Y127_SLICE_X15Y127_BO5;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A4 = CLBLM_L_X12Y127_SLICE_X17Y127_AO6;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A5 = CLBLM_R_X11Y130_SLICE_X14Y130_BO5;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_A6 = CLBLM_R_X11Y120_SLICE_X14Y120_CQ;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B1 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B2 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B3 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B4 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B5 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_B6 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C1 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C2 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C3 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C4 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C5 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_C6 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D1 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D2 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D3 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D4 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D5 = 1'b1;
  assign CLBLM_R_X13Y127_SLICE_X18Y127_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1 = CLBLM_L_X10Y126_SLICE_X12Y126_DO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C4 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C5 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C6 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B3 = CLBLL_L_X4Y122_SLICE_X4Y122_CO5;
  assign RIOB33_X105Y163_IOB_X1Y164_O = CLBLM_L_X10Y123_SLICE_X13Y123_DO5;
  assign RIOB33_X105Y163_IOB_X1Y163_O = CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B4 = CLBLL_L_X4Y124_SLICE_X4Y124_AQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B5 = CLBLM_R_X5Y124_SLICE_X6Y124_DO5;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B6 = CLBLL_L_X4Y123_SLICE_X4Y123_BQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D1 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C1 = CLBLM_R_X5Y123_SLICE_X6Y123_AQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D2 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A1 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D3 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A2 = CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A3 = CLBLM_L_X10Y124_SLICE_X13Y124_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A5 = CLBLM_L_X10Y122_SLICE_X13Y122_AQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D4 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_A6 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_AX = CLBLM_L_X10Y123_SLICE_X12Y123_DO6;
  assign LIOB33_X0Y195_IOB_X0Y195_O = LIOB33_X0Y63_IOB_X0Y64_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B1 = CLBLM_R_X7Y129_SLICE_X9Y129_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B2 = CLBLM_L_X10Y124_SLICE_X13Y124_BQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B4 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D5 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A1 = CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A2 = CLBLM_R_X5Y120_SLICE_X6Y120_BQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A3 = CLBLL_L_X4Y120_SLICE_X4Y120_AQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C1 = CLBLM_R_X11Y119_SLICE_X14Y119_BQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C2 = CLBLM_L_X10Y124_SLICE_X13Y124_CQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C3 = CLBLM_L_X10Y125_SLICE_X13Y125_CQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A5 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_A6 = CLBLL_L_X4Y121_SLICE_X5Y121_CQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_AX = CLBLM_R_X7Y123_SLICE_X8Y123_CO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B1 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_CX = CLBLM_L_X10Y124_SLICE_X12Y124_AO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_B4 = CLBLM_R_X5Y121_SLICE_X7Y121_BO6;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D1 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D2 = CLBLM_L_X8Y125_SLICE_X10Y125_CQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D4 = CLBLM_L_X10Y122_SLICE_X13Y122_BO5;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D5 = CLBLM_L_X10Y124_SLICE_X13Y124_B5Q;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C1 = CLBLM_R_X3Y123_SLICE_X3Y123_CQ;
  assign CLBLM_L_X10Y124_SLICE_X13Y124_DX = CLBLM_L_X10Y124_SLICE_X12Y124_CO6;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C2 = CLBLL_L_X4Y120_SLICE_X4Y120_AQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C4 = CLBLL_L_X4Y120_SLICE_X4Y120_A5Q;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_C5 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A1 = CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A2 = CLBLM_L_X8Y126_SLICE_X11Y126_CQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A3 = CLBLM_L_X10Y124_SLICE_X13Y124_C5Q;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A4 = CLBLM_L_X8Y121_SLICE_X11Y121_CQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_A6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D2 = CLBLL_L_X4Y120_SLICE_X4Y120_CQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_AX = CLBLM_L_X10Y121_SLICE_X13Y121_BQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D3 = CLBLL_L_X4Y120_SLICE_X4Y120_DQ;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D4 = CLBLM_R_X3Y121_SLICE_X3Y121_BQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B3 = CLBLL_L_X4Y123_SLICE_X5Y123_BQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B4 = CLBLM_R_X11Y122_SLICE_X15Y122_BQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B6 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X4Y120_D6 = CLBLM_R_X7Y123_SLICE_X9Y123_A5Q;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_B1 = CLBLM_R_X11Y124_SLICE_X14Y124_CQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C1 = CLBLM_L_X8Y126_SLICE_X11Y126_CQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C2 = CLBLM_L_X10Y125_SLICE_X12Y125_BQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C3 = CLBLM_L_X10Y124_SLICE_X13Y124_B5Q;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C5 = CLBLM_L_X10Y124_SLICE_X13Y124_C5Q;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_C6 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A1 = CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A2 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D3 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D4 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D5 = 1'b1;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_D6 = CLBLM_L_X8Y124_SLICE_X10Y124_AQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A3 = CLBLL_L_X4Y120_SLICE_X5Y120_AQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A5 = CLBLM_L_X10Y122_SLICE_X13Y122_AQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_A6 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_AX = CLBLL_L_X4Y119_SLICE_X5Y119_DO5;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B1 = CLBLL_L_X4Y120_SLICE_X5Y120_DO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B2 = CLBLL_L_X4Y120_SLICE_X5Y120_BQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B3 = CLBLL_L_X4Y120_SLICE_X5Y120_AQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B4 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_B6 = CLBLM_R_X5Y124_SLICE_X6Y124_CQ;
  assign CLBLM_L_X10Y124_SLICE_X12Y124_SR = CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C2 = CLBLL_L_X4Y120_SLICE_X5Y120_CQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C3 = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C4 = CLBLM_L_X12Y121_SLICE_X16Y121_AQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C5 = CLBLM_R_X3Y122_SLICE_X2Y122_CQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_C6 = CLBLM_R_X7Y123_SLICE_X9Y123_A5Q;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B1 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B2 = CLBLM_L_X10Y129_SLICE_X12Y129_A5Q;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D1 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D3 = CLBLM_R_X5Y123_SLICE_X7Y123_BQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D4 = 1'b1;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D5 = CLBLM_R_X3Y122_SLICE_X2Y122_CQ;
  assign CLBLL_L_X4Y120_SLICE_X5Y120_D6 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B3 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B4 = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B6 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C1 = 1'b1;
  assign RIOB33_X105Y189_IOB_X1Y190_O = CLBLM_L_X12Y126_SLICE_X16Y126_AQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C2 = 1'b1;
  assign RIOB33_X105Y189_IOB_X1Y189_O = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C3 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C4 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C5 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C6 = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_D1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOB33_X105Y165_IOB_X1Y165_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOB33_X105Y165_IOB_X1Y166_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D1 = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_T1 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D2 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = CLBLM_R_X5Y126_SLICE_X7Y126_AQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D3 = 1'b1;
  assign LIOI3_X0Y73_ILOGIC_X0Y73_D = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_D1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A5 = CLBLL_L_X4Y123_SLICE_X5Y123_CO5;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D5 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_D1 = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A6 = CLBLL_L_X4Y124_SLICE_X5Y124_CQ;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_T1 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = CLBLM_R_X5Y128_SLICE_X7Y128_B5Q;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_T1 = 1'b1;
  assign LIOB33_X0Y197_IOB_X0Y198_O = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOB33_X0Y197_IOB_X0Y197_O = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_D1 = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B3 = CLBLL_L_X4Y122_SLICE_X5Y122_BQ;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_T1 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A2 = CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A3 = CLBLM_L_X10Y125_SLICE_X13Y125_AQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A4 = CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_A6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B1 = CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A1 = CLBLM_R_X5Y122_SLICE_X7Y122_AQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A2 = CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B4 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B6 = CLBLM_L_X8Y125_SLICE_X10Y125_CQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A3 = CLBLL_L_X4Y121_SLICE_X4Y121_AQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A4 = CLBLL_L_X4Y121_SLICE_X4Y121_CQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_A6 = CLBLL_L_X4Y125_SLICE_X4Y125_BQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B2 = CLBLM_L_X10Y125_SLICE_X13Y125_BQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_B3 = CLBLM_L_X10Y125_SLICE_X13Y125_CQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C3 = CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C4 = CLBLL_L_X4Y120_SLICE_X4Y120_DQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C5 = CLBLM_L_X10Y125_SLICE_X13Y125_DO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_C6 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B1 = CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B2 = CLBLL_L_X4Y121_SLICE_X4Y121_BQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B3 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B5 = CLBLL_L_X4Y118_SLICE_X5Y118_BQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_B6 = CLBLM_R_X3Y124_SLICE_X3Y124_CQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C2 = CLBLL_L_X4Y121_SLICE_X4Y121_CQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C3 = CLBLM_R_X5Y122_SLICE_X7Y122_CO6;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C4 = CLBLM_R_X3Y121_SLICE_X2Y121_BQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D6 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_C6 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D2 = CLBLM_L_X10Y125_SLICE_X13Y125_CQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D3 = CLBLM_L_X10Y125_SLICE_X12Y125_BQ;
  assign CLBLM_L_X10Y125_SLICE_X13Y125_D4 = CLBLM_L_X10Y124_SLICE_X13Y124_CQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D2 = CLBLL_L_X4Y121_SLICE_X4Y121_AQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D4 = CLBLM_R_X3Y120_SLICE_X3Y120_BQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A6 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D5 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X4Y121_D6 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A1 = CLBLM_L_X8Y121_SLICE_X11Y121_DO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A3 = CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_A4 = CLBLM_R_X7Y125_SLICE_X9Y125_CQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B1 = CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B2 = CLBLM_L_X10Y125_SLICE_X12Y125_BQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B3 = CLBLM_L_X10Y124_SLICE_X12Y124_AO5;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B5 = CLBLM_L_X10Y125_SLICE_X13Y125_DO5;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_B6 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C2 = CLBLM_R_X11Y129_SLICE_X14Y129_BQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C3 = CLBLM_L_X8Y127_SLICE_X10Y127_CQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C4 = CLBLM_L_X10Y123_SLICE_X12Y123_DO5;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C5 = 1'b1;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_X105Y171_IOB_X1Y172_O = CLBLM_R_X103Y171_SLICE_X163Y171_BO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A1 = CLBLL_L_X4Y120_SLICE_X4Y120_CQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A3 = CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A5 = CLBLM_R_X3Y121_SLICE_X2Y121_CQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_A6 = CLBLM_R_X3Y123_SLICE_X3Y123_CQ;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D5 = CLBLM_L_X8Y125_SLICE_X11Y125_DO6;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B2 = CLBLL_L_X4Y121_SLICE_X5Y121_BQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B4 = CLBLM_R_X11Y121_SLICE_X15Y121_AQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B5 = CLBLM_R_X3Y128_SLICE_X2Y128_AO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_B6 = CLBLL_L_X4Y117_SLICE_X4Y117_AO5;
  assign CLBLM_L_X10Y125_SLICE_X12Y125_D6 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C2 = CLBLL_L_X4Y121_SLICE_X5Y121_CQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C3 = CLBLL_L_X4Y118_SLICE_X5Y118_C5Q;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C4 = CLBLM_R_X5Y121_SLICE_X7Y121_DO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_C6 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign LIOB33_SING_X0Y100_IOB_X0Y100_O = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D1 = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D2 = CLBLM_R_X5Y122_SLICE_X6Y122_CQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D3 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D4 = CLBLL_L_X4Y119_SLICE_X4Y119_CQ;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D5 = 1'b1;
  assign CLBLL_L_X4Y121_SLICE_X5Y121_D6 = CLBLL_L_X4Y120_SLICE_X4Y120_BQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D3 = CLBLL_L_X4Y124_SLICE_X4Y124_CQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A1 = CLBLM_L_X10Y124_SLICE_X13Y124_BQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A2 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A3 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A4 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A5 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_A6 = CLBLM_L_X10Y120_SLICE_X12Y120_CQ;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B1 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B2 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B3 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B4 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B5 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_B6 = 1'b1;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_D = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_D = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C1 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C2 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C3 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C4 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C5 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_C6 = 1'b1;
  assign LIOB33_X0Y79_IOB_X0Y80_O = CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_D = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_D = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D1 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D2 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D3 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D4 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D5 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X15Y119_D6 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A1 = CLBLM_R_X11Y123_SLICE_X14Y123_CQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A3 = CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A4 = CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A5 = CLBLM_L_X10Y122_SLICE_X12Y122_AQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B1 = CLBLM_R_X7Y117_SLICE_X8Y117_DQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B2 = CLBLM_R_X11Y119_SLICE_X14Y119_BQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B3 = CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B4 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_B6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOB33_X105Y167_IOB_X1Y167_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign RIOB33_X105Y167_IOB_X1Y168_O = CLBLM_R_X11Y151_SLICE_X14Y151_AO6;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C1 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C2 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C3 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C4 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C5 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_C6 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D1 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D2 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D3 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D4 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D5 = 1'b1;
  assign CLBLM_R_X11Y119_SLICE_X14Y119_D6 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B2 = CLBLM_L_X8Y128_SLICE_X11Y128_BQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B3 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B6 = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C1 = CLBLM_R_X7Y131_SLICE_X8Y131_CO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A1 = CLBLM_R_X3Y119_SLICE_X2Y119_AQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C2 = CLBLM_L_X8Y129_SLICE_X11Y129_CO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A3 = CLBLM_L_X10Y126_SLICE_X13Y126_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A4 = CLBLM_R_X11Y126_SLICE_X15Y126_DO5;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A6 = CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_A5 = CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A1 = CLBLM_R_X5Y126_SLICE_X7Y126_CO5;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A2 = CLBLM_L_X10Y121_SLICE_X12Y121_DQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B1 = CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B2 = CLBLM_L_X10Y126_SLICE_X13Y126_BQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B3 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B5 = CLBLM_R_X11Y126_SLICE_X15Y126_DO5;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_B6 = CLBLM_R_X11Y126_SLICE_X14Y126_DQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A3 = CLBLL_L_X4Y122_SLICE_X4Y122_AQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_A5 = CLBLM_R_X5Y121_SLICE_X7Y121_AQ;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_B5 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C1 = CLBLM_L_X10Y123_SLICE_X13Y123_BQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C2 = CLBLM_L_X10Y126_SLICE_X13Y126_CQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_C1 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C5 = CLBLM_L_X10Y126_SLICE_X13Y126_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_C6 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A2 = CLBLM_R_X7Y116_SLICE_X9Y116_CO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A3 = CLBLM_L_X8Y116_SLICE_X10Y116_CO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_A4 = CLBLM_L_X8Y116_SLICE_X11Y116_BO6;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D2 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D3 = CLBLM_L_X12Y127_SLICE_X16Y127_AQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D4 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D5 = CLBLL_L_X4Y122_SLICE_X5Y122_DQ;
  assign CLBLM_L_X10Y126_SLICE_X13Y126_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B3 = CLBLM_R_X3Y124_SLICE_X3Y124_DO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B4 = CLBLM_R_X7Y118_SLICE_X8Y118_C5Q;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_B6 = CLBLM_L_X8Y118_SLICE_X11Y118_CO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C1 = CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C2 = CLBLM_R_X5Y118_SLICE_X7Y118_BO5;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A1 = CLBLM_L_X10Y128_SLICE_X12Y128_CQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A2 = CLBLM_R_X11Y126_SLICE_X15Y126_DO5;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A3 = CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A5 = CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_A6 = CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_C6 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X4Y122_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D1 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D2 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D3 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D4 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B4 = CLBLL_L_X4Y122_SLICE_X5Y122_DQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D5 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X11Y116_D6 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B1 = CLBLM_L_X10Y126_SLICE_X13Y126_DQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_B3 = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C2 = CLBLM_R_X11Y123_SLICE_X14Y123_DQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C3 = CLBLM_L_X8Y126_SLICE_X11Y126_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C4 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_C6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A1 = CLBLL_L_X4Y117_SLICE_X5Y117_BQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A2 = CLBLM_R_X5Y116_SLICE_X7Y116_CQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A3 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A4 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_A5 = CLBLM_R_X7Y119_SLICE_X8Y119_DQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A1 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A2 = CLBLM_R_X5Y122_SLICE_X7Y122_BQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A3 = CLBLL_L_X4Y122_SLICE_X5Y122_AQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B2 = CLBLL_L_X4Y122_SLICE_X5Y122_BQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A4 = CLBLM_L_X10Y121_SLICE_X13Y121_B5Q;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_A5 = CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_B5 = CLBLM_R_X5Y124_SLICE_X6Y124_DO5;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B5 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_B6 = CLBLM_R_X5Y116_SLICE_X7Y116_BQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C1 = CLBLM_L_X8Y116_SLICE_X10Y116_AO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C2 = CLBLM_L_X8Y123_SLICE_X10Y123_CQ;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C3 = CLBLM_R_X3Y124_SLICE_X3Y124_DO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C4 = CLBLM_R_X3Y126_SLICE_X2Y126_BO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C5 = CLBLM_R_X7Y124_SLICE_X8Y124_B5Q;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C6 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_C6 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C1 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C3 = CLBLM_R_X5Y122_SLICE_X6Y122_AQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D1 = CLBLL_L_X4Y120_SLICE_X4Y120_C5Q;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D2 = CLBLM_R_X7Y115_SLICE_X9Y115_BO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D3 = CLBLM_R_X3Y124_SLICE_X3Y124_DO6;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D4 = 1'b1;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D5 = CLBLM_R_X7Y118_SLICE_X9Y118_BO5;
  assign CLBLM_L_X8Y116_SLICE_X10Y116_D6 = CLBLM_R_X5Y118_SLICE_X7Y118_BO5;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D1 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D2 = 1'b1;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D3 = CLBLM_L_X8Y123_SLICE_X11Y123_BQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D4 = CLBLM_R_X3Y121_SLICE_X3Y121_AQ;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y122_SLICE_X5Y122_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A1 = CLBLM_R_X11Y120_SLICE_X15Y120_AQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A2 = CLBLM_R_X5Y127_SLICE_X7Y127_BQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A4 = CLBLM_R_X11Y120_SLICE_X15Y120_BO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_A6 = CLBLM_R_X11Y122_SLICE_X14Y122_CQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D1 = CLBLM_L_X10Y125_SLICE_X12Y125_AQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B1 = CLBLM_R_X11Y121_SLICE_X15Y121_AQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B2 = CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D2 = CLBLM_R_X7Y125_SLICE_X9Y125_AQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B3 = CLBLM_R_X11Y120_SLICE_X15Y120_AQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B4 = CLBLM_R_X11Y123_SLICE_X15Y123_AQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B5 = CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_B6 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D3 = CLBLM_L_X8Y126_SLICE_X11Y126_DQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C1 = CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C2 = CLBLM_R_X11Y123_SLICE_X15Y123_AQ;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D4 = CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C3 = CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C4 = CLBLM_R_X11Y120_SLICE_X15Y120_AQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C5 = CLBLM_R_X11Y121_SLICE_X15Y121_AQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_C6 = 1'b1;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D5 = CLBLM_L_X10Y120_SLICE_X12Y120_BQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_X105Y169_IOB_X1Y170_O = CLBLM_R_X103Y171_SLICE_X163Y171_AO6;
  assign CLBLM_L_X10Y126_SLICE_X12Y126_D6 = 1'b1;
  assign RIOB33_X105Y169_IOB_X1Y169_O = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D1 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D2 = CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D3 = CLBLM_R_X11Y123_SLICE_X14Y123_CQ;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D4 = 1'b1;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D5 = CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  assign CLBLM_R_X11Y120_SLICE_X15Y120_D6 = CLBLM_R_X11Y119_SLICE_X15Y119_AO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A2 = CLBLM_R_X11Y120_SLICE_X15Y120_CO5;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A3 = CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A4 = CLBLM_R_X5Y127_SLICE_X7Y127_BQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_A6 = CLBLM_L_X8Y124_SLICE_X10Y124_AQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C3 = CLBLM_L_X10Y129_SLICE_X13Y129_CO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B2 = CLBLM_R_X11Y120_SLICE_X14Y120_BQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B4 = CLBLM_R_X11Y121_SLICE_X14Y121_AQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B5 = CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_B6 = CLBLM_R_X11Y123_SLICE_X14Y123_AQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C2 = CLBLM_R_X11Y120_SLICE_X14Y120_CQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C3 = CLBLM_R_X5Y120_SLICE_X7Y120_DO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C4 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C5 = CLBLM_L_X10Y122_SLICE_X13Y122_CQ;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_C6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C4 = CLBLM_R_X11Y129_SLICE_X15Y129_DO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D1 = CLBLM_L_X10Y121_SLICE_X13Y121_DO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D2 = CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D3 = CLBLM_R_X11Y120_SLICE_X15Y120_BO5;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D4 = CLBLM_R_X11Y120_SLICE_X15Y120_DO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D5 = CLBLM_R_X7Y120_SLICE_X9Y120_DO6;
  assign CLBLM_R_X11Y120_SLICE_X14Y120_D6 = CLBLM_L_X8Y120_SLICE_X11Y120_AO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C5 = CLBLM_R_X11Y126_SLICE_X15Y126_AQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C6 = CLBLM_R_X11Y128_SLICE_X14Y128_AO5;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A1 = CLBLM_L_X10Y127_SLICE_X13Y127_CQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A1 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A3 = CLBLL_L_X4Y123_SLICE_X4Y123_AQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A5 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A6 = CLBLM_L_X10Y129_SLICE_X12Y129_CO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A4 = CLBLM_R_X7Y129_SLICE_X8Y129_CQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A5 = CLBLM_R_X5Y124_SLICE_X6Y124_DO5;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_A6 = CLBLL_L_X4Y123_SLICE_X4Y123_CO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B2 = CLBLM_L_X10Y127_SLICE_X13Y127_BQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B3 = CLBLM_R_X11Y126_SLICE_X15Y126_CQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B4 = CLBLM_L_X8Y128_SLICE_X11Y128_AQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B5 = CLBLM_R_X11Y126_SLICE_X15Y126_DO5;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B6 = CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B1 = CLBLM_R_X5Y124_SLICE_X7Y124_CQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C1 = CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C2 = CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C3 = CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C4 = CLBLM_R_X11Y126_SLICE_X15Y126_BQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_C6 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C2 = CLBLL_L_X4Y122_SLICE_X4Y122_A5Q;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C3 = CLBLL_L_X4Y123_SLICE_X4Y123_BQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C4 = CLBLL_L_X4Y122_SLICE_X5Y122_BQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C6 = CLBLL_L_X4Y124_SLICE_X4Y124_AQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D4 = CLBLM_R_X7Y131_SLICE_X9Y131_CO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_A4 = CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_C5 = CLBLL_L_X4Y123_SLICE_X5Y123_AQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D1 = CLBLM_R_X11Y127_SLICE_X15Y127_BO6;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D2 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D3 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D4 = CLBLL_L_X4Y125_SLICE_X4Y125_CQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D5 = CLBLM_L_X10Y127_SLICE_X13Y127_CQ;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D3 = CLBLL_L_X4Y123_SLICE_X5Y123_AQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D4 = CLBLL_L_X4Y122_SLICE_X5Y122_BQ;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D1 = CLBLL_L_X4Y122_SLICE_X4Y122_CO5;
  assign CLBLL_L_X4Y123_SLICE_X4Y123_D2 = CLBLL_L_X4Y123_SLICE_X4Y123_AQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C1 = CLBLM_L_X8Y118_SLICE_X11Y118_AQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C2 = CLBLM_L_X8Y119_SLICE_X11Y119_CQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A3 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A4 = CLBLM_L_X10Y127_SLICE_X13Y127_BQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C4 = CLBLM_L_X8Y123_SLICE_X10Y123_CQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C5 = CLBLM_L_X8Y117_SLICE_X11Y117_DO6;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_C6 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D1 = CLBLL_L_X4Y120_SLICE_X4Y120_C5Q;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D2 = CLBLM_R_X7Y118_SLICE_X9Y118_AQ;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D3 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D4 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D5 = CLBLM_L_X8Y116_SLICE_X10Y116_BQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B4 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B5 = CLBLM_R_X11Y127_SLICE_X15Y127_BO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B6 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X11Y117_D6 = CLBLM_L_X10Y124_SLICE_X13Y124_D5Q;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B2 = CLBLM_L_X8Y126_SLICE_X11Y126_CQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A5 = CLBLM_R_X5Y117_SLICE_X6Y117_BQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C4 = CLBLM_L_X10Y126_SLICE_X12Y126_BO5;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A6 = CLBLM_L_X8Y116_SLICE_X10Y116_BQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C6 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C3 = CLBLM_L_X10Y127_SLICE_X12Y127_BQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_C5 = CLBLL_L_X4Y125_SLICE_X4Y125_AQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A1 = CLBLM_R_X5Y124_SLICE_X6Y124_DO5;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A2 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A3 = CLBLL_L_X4Y123_SLICE_X5Y123_AQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B4 = CLBLM_R_X5Y125_SLICE_X6Y125_BQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D2 = CLBLM_L_X10Y126_SLICE_X12Y126_A5Q;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D4 = CLBLM_L_X10Y129_SLICE_X12Y129_CO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D5 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_D6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B5 = CLBLL_L_X4Y125_SLICE_X5Y125_AQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_B6 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C1 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C2 = CLBLL_L_X4Y117_SLICE_X5Y117_BQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C3 = CLBLM_R_X5Y116_SLICE_X7Y116_CQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C4 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C5 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_C6 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_C6 = 1'b1;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D1 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D2 = CLBLL_L_X4Y117_SLICE_X5Y117_BQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D3 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D4 = CLBLM_L_X10Y119_SLICE_X12Y119_DQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D5 = CLBLM_R_X5Y116_SLICE_X7Y116_CQ;
  assign CLBLM_L_X8Y117_SLICE_X10Y117_D6 = 1'b1;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D1 = CLBLL_L_X4Y123_SLICE_X4Y123_AQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D2 = CLBLL_L_X4Y122_SLICE_X5Y122_BQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D4 = CLBLL_L_X4Y123_SLICE_X5Y123_AQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D5 = CLBLL_L_X4Y124_SLICE_X4Y124_BQ;
  assign CLBLL_L_X4Y123_SLICE_X5Y123_D6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A1 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A2 = CLBLM_R_X7Y118_SLICE_X9Y118_AQ;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1 = CLBLL_L_X2Y115_SLICE_X0Y115_AO5;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A3 = CLBLM_L_X8Y118_SLICE_X11Y118_AQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A5 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_A6 = CLBLM_R_X11Y120_SLICE_X14Y120_AQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A1 = CLBLM_R_X11Y120_SLICE_X15Y120_CO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A3 = CLBLM_R_X11Y121_SLICE_X15Y121_AQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A4 = CLBLM_R_X5Y127_SLICE_X7Y127_BQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A5 = CLBLM_R_X11Y126_SLICE_X14Y126_AQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C2 = 1'b1;
  assign RIOB33_X105Y171_IOB_X1Y171_O = CLBLM_R_X103Y171_SLICE_X163Y171_AO5;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B1 = CLBLM_R_X11Y121_SLICE_X15Y121_DO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B2 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B3 = CLBLM_R_X11Y123_SLICE_X14Y123_CQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B4 = CLBLM_R_X11Y121_SLICE_X14Y121_DO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B5 = CLBLM_L_X10Y120_SLICE_X12Y120_CQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_B6 = CLBLM_L_X10Y124_SLICE_X13Y124_BQ;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C4 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B1 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C1 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C2 = CLBLM_R_X11Y120_SLICE_X15Y120_BO5;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C3 = CLBLM_R_X7Y120_SLICE_X9Y120_DO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C4 = CLBLM_R_X11Y123_SLICE_X14Y123_CQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B2 = CLBLM_L_X8Y118_SLICE_X11Y118_BQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C5 = CLBLM_R_X11Y119_SLICE_X14Y119_AQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_C6 = CLBLM_R_X11Y121_SLICE_X15Y121_BO6;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C5 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B3 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D1 = CLBLM_R_X11Y121_SLICE_X14Y121_AQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D2 = CLBLM_L_X10Y121_SLICE_X12Y121_BQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D3 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D4 = CLBLM_R_X11Y122_SLICE_X15Y122_AQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B5 = CLBLM_R_X5Y118_SLICE_X7Y118_AQ;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D5 = 1'b1;
  assign CLBLM_R_X11Y121_SLICE_X15Y121_D6 = CLBLM_R_X11Y122_SLICE_X15Y122_BQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_T1 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_B6 = CLBLM_L_X8Y119_SLICE_X11Y119_CQ;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_D = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A1 = CLBLL_L_X4Y124_SLICE_X4Y124_DQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A2 = CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A3 = CLBLM_R_X11Y121_SLICE_X14Y121_AQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_A6 = CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B3 = CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B4 = CLBLM_R_X11Y123_SLICE_X14Y123_BQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B5 = CLBLM_R_X11Y121_SLICE_X14Y121_BQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_B6 = CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C1 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C2 = CLBLM_R_X11Y121_SLICE_X14Y121_CQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C3 = CLBLM_L_X12Y121_SLICE_X16Y121_AQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C4 = CLBLM_L_X8Y121_SLICE_X10Y121_CQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C2 = CLBLL_L_X4Y117_SLICE_X5Y117_BQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_C6 = CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C3 = CLBLM_L_X10Y119_SLICE_X13Y119_DO6;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D1 = CLBLM_R_X11Y121_SLICE_X14Y121_BQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D2 = CLBLM_R_X11Y121_SLICE_X14Y121_CQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D3 = CLBLM_L_X12Y121_SLICE_X16Y121_AQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D4 = CLBLM_R_X11Y120_SLICE_X14Y120_BQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D5 = CLBLM_R_X11Y123_SLICE_X14Y123_BQ;
  assign CLBLM_R_X11Y121_SLICE_X14Y121_D6 = CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_D = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_D = LIOB33_X0Y61_IOB_X0Y61_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_D = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_D = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A1 = CLBLM_R_X5Y123_SLICE_X6Y123_AQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A2 = CLBLL_L_X4Y122_SLICE_X4Y122_A5Q;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A3 = CLBLL_L_X4Y124_SLICE_X4Y124_AQ;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A2 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A1 = CLBLM_L_X8Y128_SLICE_X11Y128_DQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A2 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A4 = CLBLM_R_X11Y128_SLICE_X14Y128_BO6;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A5 = CLBLM_R_X11Y127_SLICE_X15Y127_BO5;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_A6 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B1 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B1 = CLBLM_R_X11Y126_SLICE_X15Y126_DO5;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B2 = CLBLM_L_X10Y128_SLICE_X13Y128_BQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B3 = CLBLM_L_X10Y126_SLICE_X13Y126_AQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B4 = CLBLM_R_X7Y125_SLICE_X8Y125_BQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_B6 = CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C1 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C1 = CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C2 = CLBLM_L_X10Y125_SLICE_X13Y125_DO5;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C3 = CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C4 = CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C5 = CLBLM_R_X11Y126_SLICE_X15Y126_BQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_C6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C3 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D1 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D1 = CLBLM_L_X10Y128_SLICE_X13Y128_CO5;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D3 = CLBLM_L_X10Y127_SLICE_X13Y127_BQ;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D5 = CLBLM_R_X11Y126_SLICE_X15Y126_DO5;
  assign CLBLM_L_X10Y128_SLICE_X13Y128_D6 = CLBLM_L_X8Y129_SLICE_X11Y129_BQ;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D5 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C4 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A3 = CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A4 = CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C5 = CLBLM_R_X5Y116_SLICE_X7Y116_CQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_C6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D1 = CLBLM_R_X7Y118_SLICE_X9Y118_AQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D2 = CLBLM_R_X5Y116_SLICE_X7Y116_BQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B1 = CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B2 = CLBLM_L_X10Y128_SLICE_X12Y128_BQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B3 = CLBLM_L_X8Y128_SLICE_X10Y128_CQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B4 = CLBLM_L_X10Y127_SLICE_X13Y127_BQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_B6 = CLBLM_R_X11Y126_SLICE_X15Y126_DO5;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D3 = CLBLM_R_X7Y118_SLICE_X8Y118_AQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D4 = CLBLM_L_X8Y119_SLICE_X11Y119_CQ;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D5 = CLBLM_L_X8Y118_SLICE_X11Y118_AQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A3 = CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A4 = CLBLL_L_X4Y120_SLICE_X5Y120_BQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A5 = CLBLL_L_X4Y123_SLICE_X4Y123_AQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A6 = CLBLL_L_X4Y125_SLICE_X4Y125_BQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C2 = CLBLM_L_X10Y128_SLICE_X12Y128_CQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B1 = CLBLL_L_X4Y122_SLICE_X4Y122_DQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C3 = CLBLM_L_X10Y126_SLICE_X13Y126_BQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B1 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C4 = CLBLM_R_X11Y126_SLICE_X15Y126_DO5;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C5 = CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_C6 = CLBLM_R_X7Y126_SLICE_X8Y126_CQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D1 = CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D2 = CLBLM_R_X11Y126_SLICE_X15Y126_BQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D3 = CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D5 = CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_D6 = CLBLM_L_X8Y129_SLICE_X11Y129_BQ;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C4 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B1 = CLBLM_R_X7Y118_SLICE_X9Y118_CO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C6 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B2 = CLBLM_L_X8Y118_SLICE_X10Y118_BQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D1 = CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D2 = CLBLL_L_X4Y123_SLICE_X5Y123_B5Q;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D3 = CLBLL_L_X4Y124_SLICE_X5Y124_DQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D4 = CLBLL_L_X4Y122_SLICE_X5Y122_DQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D5 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B4 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B5 = CLBLM_L_X8Y118_SLICE_X11Y118_AQ;
  assign RIOB33_X105Y173_IOB_X1Y173_O = CLBLM_R_X103Y171_SLICE_X163Y171_BO5;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C4 = CLBLM_L_X10Y128_SLICE_X13Y128_BQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D5 = CLBLM_L_X8Y129_SLICE_X10Y129_DO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A1 = CLBLM_R_X11Y126_SLICE_X15Y126_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A2 = CLBLM_R_X11Y122_SLICE_X15Y122_BQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A5 = CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_A6 = CLBLM_R_X11Y122_SLICE_X15Y122_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C5 = CLBLM_R_X5Y125_SLICE_X7Y125_BQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C1 = CLBLM_L_X8Y118_SLICE_X10Y118_BQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B2 = CLBLM_R_X11Y122_SLICE_X15Y122_BQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C2 = CLBLM_L_X8Y118_SLICE_X10Y118_CQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B3 = CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B4 = CLBLM_R_X7Y126_SLICE_X9Y126_BQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D6 = CLBLM_R_X7Y128_SLICE_X9Y128_DO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C3 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_B6 = CLBLM_L_X10Y124_SLICE_X13Y124_BQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C1 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C2 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C4 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C3 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C4 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C5 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_C6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C6 = CLBLM_R_X11Y126_SLICE_X15Y126_DO5;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D3 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D4 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D1 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D2 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D3 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D4 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D5 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X15Y122_D6 = 1'b1;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A1 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A3 = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A4 = CLBLM_L_X8Y122_SLICE_X11Y122_A5Q;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_A6 = CLBLM_L_X8Y122_SLICE_X11Y122_BO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B1 = CLBLM_R_X11Y122_SLICE_X14Y122_CQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B2 = CLBLM_R_X11Y122_SLICE_X14Y122_BQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B5 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_B6 = CLBLM_R_X11Y124_SLICE_X14Y124_A5Q;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A5 = CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C1 = CLBLM_L_X10Y119_SLICE_X12Y119_AQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_A6 = CLBLM_R_X5Y124_SLICE_X6Y124_DO5;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C4 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C5 = CLBLM_R_X11Y122_SLICE_X14Y122_CQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_C6 = CLBLM_R_X11Y124_SLICE_X14Y124_BQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_AX = CLBLM_R_X7Y124_SLICE_X9Y124_BO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D1 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D2 = CLBLM_L_X8Y122_SLICE_X11Y122_BO6;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D3 = CLBLM_R_X11Y122_SLICE_X14Y122_DQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D4 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D5 = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D2 = CLBLM_L_X8Y118_SLICE_X10Y118_AQ;
  assign CLBLM_R_X11Y122_SLICE_X14Y122_D6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B1 = CLBLL_L_X4Y123_SLICE_X4Y123_DO6;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D4 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B3 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D5 = CLBLM_R_X3Y123_SLICE_X2Y123_DQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B4 = CLBLM_R_X5Y124_SLICE_X6Y124_DO5;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_D6 = CLBLM_R_X3Y126_SLICE_X3Y126_AO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B5 = CLBLL_L_X4Y124_SLICE_X4Y124_BQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_B6 = CLBLM_R_X5Y120_SLICE_X6Y120_CQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C1 = CLBLL_L_X4Y124_SLICE_X4Y124_BQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C2 = CLBLL_L_X4Y124_SLICE_X4Y124_CQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C3 = CLBLM_R_X3Y123_SLICE_X3Y123_AQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A1 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A2 = CLBLM_R_X3Y122_SLICE_X3Y122_BQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C4 = CLBLM_R_X5Y124_SLICE_X6Y124_DO5;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A4 = CLBLM_L_X8Y121_SLICE_X10Y121_AO5;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_A6 = CLBLM_L_X8Y124_SLICE_X11Y124_BQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C5 = CLBLL_L_X4Y123_SLICE_X4Y123_DO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A1 = CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B1 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A3 = CLBLM_L_X10Y129_SLICE_X13Y129_AQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A4 = CLBLM_L_X10Y124_SLICE_X13Y124_DQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A6 = CLBLM_R_X11Y121_SLICE_X14Y121_BQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B2 = CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B3 = CLBLM_R_X3Y124_SLICE_X3Y124_C5Q;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B1 = CLBLM_R_X11Y126_SLICE_X15Y126_BQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B2 = CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B3 = CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B4 = CLBLM_L_X8Y129_SLICE_X11Y129_BQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B5 = CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_B6 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C1 = CLBLM_R_X3Y130_SLICE_X3Y130_BO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C2 = CLBLL_L_X2Y127_SLICE_X0Y127_CO6;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C1 = CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C2 = CLBLM_R_X11Y126_SLICE_X15Y126_BQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C3 = CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C4 = CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C5 = CLBLM_L_X10Y125_SLICE_X13Y125_DO5;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_C6 = CLBLM_L_X8Y129_SLICE_X11Y129_BQ;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A2 = CLBLM_R_X11Y120_SLICE_X14Y120_BQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A5 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_D1 = CLBLL_L_X4Y126_SLICE_X4Y126_CO5;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D1 = CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D3 = CLBLM_L_X10Y125_SLICE_X13Y125_AQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D4 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_D6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B4 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C1 = CLBLM_L_X8Y118_SLICE_X11Y118_AQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C2 = CLBLM_L_X8Y119_SLICE_X11Y119_CQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A2 = CLBLM_L_X10Y129_SLICE_X12Y129_BQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A3 = CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A4 = CLBLM_R_X11Y127_SLICE_X15Y127_CO5;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A5 = CLBLM_L_X10Y129_SLICE_X13Y129_BO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_A6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D1 = CLBLM_R_X3Y131_SLICE_X2Y131_AQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_AX = CLBLM_L_X8Y124_SLICE_X11Y124_CO6;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D2 = CLBLM_R_X5Y124_SLICE_X7Y124_CQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B5 = CLBLM_L_X10Y129_SLICE_X12Y129_CO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_B6 = CLBLM_L_X10Y129_SLICE_X12Y129_A5Q;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D3 = CLBLL_L_X4Y124_SLICE_X4Y124_DQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D3 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D4 = CLBLM_L_X8Y116_SLICE_X10Y116_AO5;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C1 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B1 = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B2 = CLBLL_L_X4Y125_SLICE_X5Y125_BQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B3 = CLBLL_L_X4Y124_SLICE_X5Y124_BQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C5 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C1 = CLBLM_R_X5Y125_SLICE_X7Y125_AQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C2 = CLBLL_L_X4Y124_SLICE_X5Y124_BQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C3 = CLBLL_L_X2Y129_SLICE_X0Y129_AO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C4 = CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C5 = CLBLM_R_X3Y130_SLICE_X3Y130_AO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_C6 = CLBLL_L_X4Y126_SLICE_X4Y126_BO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B2 = CLBLM_L_X8Y119_SLICE_X10Y119_BQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B3 = CLBLM_R_X3Y120_SLICE_X2Y120_CQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B5 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_B6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C1 = CLBLM_R_X7Y119_SLICE_X8Y119_DQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D1 = CLBLL_L_X4Y126_SLICE_X4Y126_CO5;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D2 = CLBLL_L_X2Y129_SLICE_X0Y129_AO6;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D3 = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D4 = CLBLM_R_X5Y122_SLICE_X6Y122_AQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D5 = CLBLM_R_X7Y125_SLICE_X9Y125_DQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_D6 = CLBLL_L_X4Y126_SLICE_X4Y126_BO6;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C4 = CLBLM_L_X8Y116_SLICE_X10Y116_AO5;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C5 = CLBLM_L_X8Y125_SLICE_X10Y125_DQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D1 = CLBLM_R_X5Y116_SLICE_X6Y116_AQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D2 = CLBLM_L_X10Y119_SLICE_X12Y119_CQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D3 = CLBLM_R_X7Y119_SLICE_X8Y119_CQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D4 = CLBLM_L_X10Y119_SLICE_X12Y119_DQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D5 = CLBLM_R_X7Y119_SLICE_X8Y119_DQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_D6 = CLBLM_L_X8Y119_SLICE_X11Y119_BQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D1 = CLBLM_L_X10Y125_SLICE_X13Y125_DO5;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A1 = CLBLM_R_X11Y126_SLICE_X14Y126_AO5;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A2 = CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A3 = CLBLM_R_X11Y123_SLICE_X15Y123_AQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A4 = CLBLM_R_X11Y127_SLICE_X14Y127_AQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_A6 = CLBLM_R_X11Y120_SLICE_X15Y120_BO5;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_D1 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B2 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B3 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B4 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B5 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_B6 = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_T1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C2 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C3 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C4 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C5 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_C6 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_D1 = CLBLM_R_X3Y125_SLICE_X2Y125_AQ;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_D1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_T1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D2 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D3 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D4 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D5 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X15Y123_D6 = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_T1 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_D1 = CLBLM_R_X103Y171_SLICE_X163Y171_BO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_D1 = CLBLM_L_X8Y123_SLICE_X10Y123_C5Q;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A1 = CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A2 = CLBLM_R_X11Y119_SLICE_X14Y119_BQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A3 = CLBLM_R_X11Y123_SLICE_X14Y123_AQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_A6 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_T1 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_T1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B1 = CLBLM_R_X11Y120_SLICE_X14Y120_BQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B2 = CLBLM_R_X11Y123_SLICE_X14Y123_BQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B4 = CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_B6 = CLBLM_L_X10Y126_SLICE_X13Y126_BQ;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_D1 = CLBLM_R_X103Y171_SLICE_X163Y171_AO5;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = CLBLM_L_X10Y120_SLICE_X13Y120_AQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C2 = CLBLM_R_X11Y123_SLICE_X14Y123_CQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C4 = CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C5 = CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_C6 = CLBLM_R_X11Y121_SLICE_X14Y121_BQ;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_T1 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D2 = CLBLM_R_X11Y123_SLICE_X14Y123_CQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_A2 = CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D4 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D5 = 1'b1;
  assign CLBLM_R_X11Y123_SLICE_X14Y123_D6 = CLBLM_R_X5Y124_SLICE_X6Y124_CQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B2 = CLBLL_L_X4Y124_SLICE_X5Y124_BQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B3 = CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B5 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A1 = CLBLM_R_X5Y128_SLICE_X6Y128_DQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A2 = CLBLM_R_X5Y128_SLICE_X6Y128_A5Q;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A3 = CLBLM_R_X7Y122_SLICE_X9Y122_AQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A5 = CLBLL_L_X4Y129_SLICE_X5Y129_AQ;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_A6 = CLBLL_L_X4Y119_SLICE_X4Y119_DQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_B6 = CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B2 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_B6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A1 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A2 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A3 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C2 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_C6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A4 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A5 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B1 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B2 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A1 = CLBLM_L_X8Y120_SLICE_X11Y120_DO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D1 = CLBLL_L_X2Y129_SLICE_X1Y129_CO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D2 = CLBLL_L_X2Y126_SLICE_X0Y126_BO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D3 = CLBLL_L_X4Y129_SLICE_X5Y129_DO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D4 = CLBLL_L_X4Y126_SLICE_X5Y126_DO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D5 = CLBLM_R_X3Y128_SLICE_X2Y128_DO6;
  assign CLBLL_L_X4Y126_SLICE_X4Y126_D6 = CLBLL_L_X4Y125_SLICE_X5Y125_DO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A2 = CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A3 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A4 = CLBLM_L_X10Y121_SLICE_X12Y121_BQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A5 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_A6 = CLBLM_L_X8Y120_SLICE_X11Y120_CO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B1 = CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B2 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B3 = CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B4 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B5 = CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_B6 = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C1 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C2 = CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C3 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C4 = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C5 = CLBLM_L_X10Y124_SLICE_X13Y124_BQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_C6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D3 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D4 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A1 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A2 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A3 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A4 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A5 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D1 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A1 = CLBLL_L_X4Y126_SLICE_X4Y126_CO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A2 = CLBLM_R_X3Y130_SLICE_X3Y130_AO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A3 = CLBLM_L_X10Y125_SLICE_X13Y125_AQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A4 = CLBLL_L_X4Y121_SLICE_X5Y121_BQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_A6 = CLBLM_L_X8Y126_SLICE_X11Y126_AQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D2 = CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D3 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B1 = CLBLL_L_X2Y129_SLICE_X0Y129_AO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B2 = CLBLL_L_X4Y126_SLICE_X4Y126_BO6;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B3 = CLBLL_L_X4Y124_SLICE_X5Y124_AQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B5 = CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A3 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A4 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A5 = CLBLM_L_X8Y126_SLICE_X11Y126_CQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_A6 = CLBLM_R_X5Y119_SLICE_X7Y119_CQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B4 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B1 = CLBLM_L_X10Y122_SLICE_X13Y122_CQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C5 = CLBLL_L_X4Y126_SLICE_X4Y126_CO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B2 = CLBLM_R_X5Y116_SLICE_X7Y116_CQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B3 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_B6 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C2 = CLBLM_R_X5Y120_SLICE_X7Y120_BQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C4 = CLBLM_R_X7Y126_SLICE_X9Y126_B5Q;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C1 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D1 = CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D2 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D3 = CLBLM_L_X8Y128_SLICE_X10Y128_CQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D4 = CLBLL_L_X4Y126_SLICE_X4Y126_BO5;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D5 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_D6 = CLBLM_R_X3Y130_SLICE_X3Y130_AO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C2 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C3 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C4 = CLBLM_R_X5Y119_SLICE_X7Y119_BQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C5 = CLBLM_R_X7Y120_SLICE_X8Y120_CQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_C6 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_SR = CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D1 = CLBLM_L_X8Y125_SLICE_X10Y125_AQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D2 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D3 = CLBLM_R_X7Y120_SLICE_X8Y120_CQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D4 = CLBLM_L_X12Y121_SLICE_X16Y121_AQ;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D5 = 1'b1;
  assign CLBLM_L_X8Y120_SLICE_X10Y120_D6 = CLBLM_L_X10Y120_SLICE_X12Y120_CQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D2 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A1 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A2 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A3 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A4 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A5 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_A6 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B1 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B2 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B3 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B4 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B5 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_B6 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C1 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C2 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C3 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C4 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C5 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_C6 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D1 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D2 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D3 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D4 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D5 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X15Y124_D6 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_T1 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A1 = CLBLM_R_X3Y123_SLICE_X3Y123_BQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A3 = CLBLM_R_X11Y124_SLICE_X14Y124_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A4 = CLBLM_L_X8Y119_SLICE_X10Y119_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_A6 = 1'b1;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B2 = CLBLM_R_X11Y124_SLICE_X14Y124_BQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B3 = CLBLM_R_X3Y124_SLICE_X3Y124_C5Q;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B4 = CLBLM_L_X8Y124_SLICE_X11Y124_DO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_B6 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C2 = CLBLM_R_X11Y124_SLICE_X14Y124_CQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C3 = CLBLM_R_X5Y121_SLICE_X7Y121_DO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C4 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_C6 = CLBLM_L_X12Y126_SLICE_X16Y126_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D1 = CLBLM_R_X11Y122_SLICE_X14Y122_AQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D2 = CLBLM_R_X7Y119_SLICE_X9Y119_BQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D3 = CLBLM_R_X11Y124_SLICE_X14Y124_BQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A4 = CLBLM_R_X7Y131_SLICE_X9Y131_BO6;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D4 = CLBLM_R_X11Y120_SLICE_X14Y120_CQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D5 = CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  assign CLBLM_R_X11Y124_SLICE_X14Y124_D6 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B1 = CLBLM_R_X7Y127_SLICE_X9Y127_AQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B2 = CLBLM_R_X5Y129_SLICE_X6Y129_CQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A1 = CLBLL_L_X2Y128_SLICE_X1Y128_AO5;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A2 = CLBLM_R_X3Y121_SLICE_X2Y121_AQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A3 = CLBLL_L_X2Y130_SLICE_X0Y130_CO5;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A4 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A5 = CLBLL_L_X2Y130_SLICE_X0Y130_AO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_A6 = CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B1 = CLBLM_R_X7Y126_SLICE_X9Y126_C5Q;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B2 = CLBLL_L_X2Y126_SLICE_X0Y126_AO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B3 = CLBLM_R_X5Y126_SLICE_X7Y126_BQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B4 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_B6 = CLBLM_R_X3Y127_SLICE_X3Y127_DO6;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A5 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_A6 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C1 = CLBLM_R_X3Y122_SLICE_X2Y122_DQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C2 = CLBLL_L_X2Y130_SLICE_X0Y130_BO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C3 = CLBLL_L_X2Y130_SLICE_X0Y130_CO5;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C4 = CLBLL_L_X2Y128_SLICE_X1Y128_AO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C5 = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_C6 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C1 = CLBLM_L_X8Y128_SLICE_X11Y128_CQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C2 = CLBLM_L_X8Y129_SLICE_X10Y129_AO5;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D1 = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D2 = CLBLL_L_X2Y130_SLICE_X0Y130_BO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D3 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D4 = CLBLL_L_X2Y130_SLICE_X0Y130_AO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A2 = CLBLM_R_X5Y120_SLICE_X7Y120_BQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A3 = CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A4 = CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A5 = CLBLM_R_X11Y122_SLICE_X15Y122_AQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D5 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X4Y127_D6 = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B2 = CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B3 = CLBLM_L_X8Y121_SLICE_X11Y121_AQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B5 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_B6 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_L_X10Y127_SLICE_X12Y127_B3 = CLBLM_R_X3Y121_SLICE_X2Y121_CQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C2 = CLBLM_L_X8Y121_SLICE_X11Y121_CQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C3 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C4 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_C6 = CLBLM_R_X7Y120_SLICE_X8Y120_AQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A1 = CLBLM_R_X5Y127_SLICE_X7Y127_DO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A2 = CLBLM_R_X7Y125_SLICE_X9Y125_CQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A3 = CLBLL_L_X4Y127_SLICE_X4Y127_CO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A4 = CLBLL_L_X4Y127_SLICE_X5Y127_BO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A5 = CLBLL_L_X4Y127_SLICE_X5Y127_CO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_A6 = CLBLL_L_X2Y128_SLICE_X0Y128_AO5;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D1 = CLBLM_R_X3Y123_SLICE_X2Y123_DQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D6 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B1 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B2 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B3 = CLBLL_L_X2Y130_SLICE_X1Y130_AO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B4 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B5 = CLBLL_L_X4Y124_SLICE_X5Y124_CQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_B6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A3 = CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A6 = 1'b1;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C1 = CLBLL_L_X2Y130_SLICE_X0Y130_CO5;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C5 = CLBLM_R_X3Y121_SLICE_X2Y121_C5Q;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C2 = CLBLL_L_X2Y130_SLICE_X0Y130_AO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B1 = CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B3 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B4 = CLBLM_L_X8Y126_SLICE_X11Y126_B5Q;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_B6 = CLBLL_L_X4Y119_SLICE_X4Y119_CQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C6 = CLBLL_L_X2Y130_SLICE_X0Y130_BO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D2 = CLBLL_L_X2Y128_SLICE_X1Y128_AO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D3 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C2 = CLBLM_L_X8Y121_SLICE_X10Y121_CQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C3 = CLBLM_L_X8Y118_SLICE_X10Y118_AO5;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C4 = CLBLM_L_X8Y124_SLICE_X10Y124_CO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C5 = CLBLM_R_X7Y119_SLICE_X9Y119_AQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_C6 = CLBLM_R_X7Y119_SLICE_X9Y119_CO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D4 = CLBLL_L_X2Y130_SLICE_X0Y130_BO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D5 = CLBLM_R_X5Y125_SLICE_X7Y125_BQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D6 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D1 = CLBLM_R_X3Y122_SLICE_X2Y122_A5Q;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D2 = CLBLM_L_X8Y121_SLICE_X10Y121_CQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D3 = CLBLL_L_X4Y122_SLICE_X5Y122_DQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D5 = CLBLM_L_X10Y122_SLICE_X13Y122_CQ;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_D6 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B2 = CLBLM_R_X11Y126_SLICE_X14Y126_BQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A1 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A2 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A3 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A4 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A5 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_A6 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B1 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B2 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B3 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B4 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B5 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_B6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A1 = CLBLL_L_X4Y117_SLICE_X5Y117_BQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A2 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A3 = CLBLM_R_X5Y116_SLICE_X6Y116_AQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A4 = CLBLM_R_X5Y116_SLICE_X7Y116_CQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A5 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_A6 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C1 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C2 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C3 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B1 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B2 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B3 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B4 = CLBLM_R_X5Y116_SLICE_X7Y116_CQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B5 = CLBLM_L_X10Y119_SLICE_X12Y119_CQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_B6 = CLBLL_L_X4Y117_SLICE_X5Y117_BQ;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D1 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C3 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_C6 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D3 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D4 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A1 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A2 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A3 = CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A4 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_A6 = CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D3 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X9Y115_D6 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B1 = CLBLM_L_X10Y124_SLICE_X13Y124_CQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B2 = CLBLM_R_X11Y125_SLICE_X14Y125_BQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B5 = CLBLM_L_X8Y124_SLICE_X10Y124_DO6;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A1 = CLBLL_L_X4Y117_SLICE_X5Y117_BQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A2 = CLBLM_R_X5Y116_SLICE_X7Y116_CQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A3 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A4 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A5 = CLBLM_R_X5Y119_SLICE_X6Y119_CQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_A6 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C2 = CLBLM_R_X11Y125_SLICE_X14Y125_CQ;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C4 = CLBLM_R_X11Y126_SLICE_X14Y126_CQ;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B3 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_B6 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D1 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C3 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_C6 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D3 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D4 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D5 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_D6 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D1 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D2 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D3 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D4 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D5 = 1'b1;
  assign CLBLM_R_X7Y115_SLICE_X8Y115_D6 = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_D1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A1 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A2 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C4 = CLBLM_R_X7Y131_SLICE_X9Y131_CO6;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_A3 = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_T1 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_D1 = CLBLL_L_X2Y118_SLICE_X1Y118_B5Q;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_D1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A1 = CLBLL_L_X4Y128_SLICE_X4Y128_DO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A2 = CLBLL_L_X4Y126_SLICE_X5Y126_BO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A3 = CLBLL_L_X2Y129_SLICE_X1Y129_CO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A4 = CLBLL_L_X4Y128_SLICE_X4Y128_BO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A5 = CLBLL_L_X4Y127_SLICE_X4Y127_BO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_A6 = CLBLM_R_X3Y128_SLICE_X3Y128_DO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_T1 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_D1 = CLBLM_R_X103Y173_SLICE_X163Y173_AO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B1 = CLBLM_R_X5Y128_SLICE_X7Y128_CO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B2 = CLBLL_L_X4Y128_SLICE_X5Y128_DO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B3 = CLBLL_L_X4Y127_SLICE_X4Y127_AO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B4 = CLBLM_R_X3Y130_SLICE_X2Y130_BO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B5 = CLBLL_L_X4Y119_SLICE_X4Y119_AQ;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_B6 = CLBLL_L_X4Y128_SLICE_X4Y128_CO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_D1 = CLBLL_L_X4Y126_SLICE_X4Y126_AQ;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_T1 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C1 = CLBLL_L_X2Y128_SLICE_X1Y128_AO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C2 = CLBLL_L_X2Y130_SLICE_X0Y130_CO5;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C3 = CLBLM_R_X7Y123_SLICE_X9Y123_BQ;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C4 = CLBLL_L_X2Y130_SLICE_X0Y130_BO6;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_C6 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_T1 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_D1 = CLBLM_R_X103Y171_SLICE_X163Y171_BO5;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D1 = CLBLL_L_X4Y126_SLICE_X4Y126_CO5;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D2 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D3 = CLBLL_L_X4Y119_SLICE_X5Y119_CQ;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D4 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D5 = 1'b1;
  assign CLBLL_L_X4Y128_SLICE_X4Y128_D6 = CLBLM_R_X3Y130_SLICE_X3Y130_AO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_T1 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A1 = CLBLM_R_X5Y128_SLICE_X7Y128_AQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A3 = CLBLM_R_X7Y118_SLICE_X8Y118_AQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A4 = CLBLM_L_X10Y122_SLICE_X13Y122_C5Q;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1 = CLBLM_L_X10Y123_SLICE_X13Y123_DO5;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B1 = CLBLM_L_X8Y123_SLICE_X11Y123_DO5;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B2 = CLBLL_L_X4Y128_SLICE_X4Y128_AO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B3 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B5 = CLBLM_R_X3Y123_SLICE_X2Y123_DQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_B6 = CLBLM_L_X8Y118_SLICE_X10Y118_AO5;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D3 = CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D4 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C1 = CLBLM_L_X8Y123_SLICE_X11Y123_BQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C2 = CLBLM_L_X10Y122_SLICE_X12Y122_DO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C3 = CLBLM_L_X8Y122_SLICE_X10Y122_DO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C4 = CLBLM_L_X10Y121_SLICE_X12Y121_DQ;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C5 = CLBLM_L_X8Y122_SLICE_X11Y122_DO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_C6 = CLBLL_L_X4Y123_SLICE_X5Y123_BQ;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A1 = CLBLM_R_X7Y126_SLICE_X8Y126_CQ;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A2 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A4 = CLBLL_L_X2Y130_SLICE_X0Y130_CO5;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A5 = CLBLL_L_X2Y130_SLICE_X0Y130_AO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_A6 = CLBLL_L_X2Y130_SLICE_X0Y130_BO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D1 = CLBLM_L_X10Y122_SLICE_X13Y122_C5Q;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B1 = CLBLM_R_X5Y123_SLICE_X7Y123_AQ;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B2 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D4 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D5 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D6 = CLBLM_R_X5Y125_SLICE_X6Y125_BQ;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B3 = CLBLL_L_X2Y128_SLICE_X1Y128_AO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B4 = CLBLL_L_X4Y125_SLICE_X5Y125_AQ;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B5 = CLBLL_L_X2Y130_SLICE_X0Y130_CO5;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_B6 = CLBLL_L_X2Y128_SLICE_X1Y128_AO5;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C2 = CLBLL_L_X2Y128_SLICE_X0Y128_AO5;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C3 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C5 = CLBLM_R_X3Y128_SLICE_X3Y128_AO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A5 = CLBLM_L_X8Y120_SLICE_X10Y120_BQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A6 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A2 = CLBLM_R_X5Y122_SLICE_X7Y122_AQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_A4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C4 = CLBLM_R_X5Y127_SLICE_X6Y127_DO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C6 = CLBLL_L_X4Y128_SLICE_X5Y128_BO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B1 = CLBLM_L_X8Y122_SLICE_X11Y122_CO6;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D5 = CLBLM_L_X10Y129_SLICE_X13Y129_AQ;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_D6 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B4 = CLBLL_L_X4Y122_SLICE_X4Y122_DQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B5 = CLBLM_L_X8Y122_SLICE_X11Y122_AQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B6 = CLBLM_L_X8Y122_SLICE_X10Y122_CO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_BX = CLBLM_L_X10Y122_SLICE_X13Y122_BO6;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C1 = CLBLM_L_X8Y120_SLICE_X10Y120_BQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C4 = CLBLM_L_X10Y122_SLICE_X13Y122_DQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C2 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C6 = CLBLM_L_X8Y124_SLICE_X10Y124_BQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C3 = CLBLM_R_X7Y121_SLICE_X9Y121_B5Q;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_C5 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D1 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D2 = CLBLM_L_X10Y122_SLICE_X13Y122_CQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D3 = CLBLM_L_X8Y122_SLICE_X10Y122_A5Q;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D4 = CLBLM_R_X5Y123_SLICE_X6Y123_CQ;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D5 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_D6 = CLBLM_L_X10Y122_SLICE_X12Y122_BQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A1 = CLBLM_L_X8Y119_SLICE_X11Y119_DO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A3 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_A4 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A1 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A2 = CLBLM_R_X11Y127_SLICE_X15Y127_BO5;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A3 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A4 = CLBLM_R_X11Y128_SLICE_X15Y128_BO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A5 = CLBLM_R_X11Y130_SLICE_X14Y130_BO5;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B1 = CLBLM_R_X11Y126_SLICE_X15Y126_DO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B2 = CLBLM_R_X11Y129_SLICE_X15Y129_AO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B4 = CLBLL_L_X4Y125_SLICE_X5Y125_BQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_B6 = CLBLM_R_X11Y126_SLICE_X15Y126_BQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A2 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A3 = CLBLM_R_X7Y116_SLICE_X9Y116_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A4 = CLBLM_R_X7Y118_SLICE_X8Y118_C5Q;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A5 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C2 = CLBLM_R_X11Y126_SLICE_X15Y126_CQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_C3 = CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B1 = CLBLM_R_X7Y116_SLICE_X9Y116_DO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B4 = CLBLM_L_X8Y119_SLICE_X10Y119_BQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B2 = CLBLM_L_X8Y119_SLICE_X11Y119_BQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B5 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_B6 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B3 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C1 = CLBLM_R_X7Y115_SLICE_X8Y115_AO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C2 = CLBLM_R_X7Y117_SLICE_X9Y117_AO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C3 = CLBLM_L_X10Y120_SLICE_X13Y120_A5Q;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C4 = CLBLM_R_X3Y124_SLICE_X3Y124_DO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C5 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_C6 = CLBLM_R_X3Y126_SLICE_X2Y126_BO6;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D4 = CLBLM_R_X11Y126_SLICE_X15Y126_BQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A1 = CLBLM_L_X10Y127_SLICE_X13Y127_DQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B5 = CLBLL_L_X4Y122_SLICE_X4Y122_A5Q;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C4 = CLBLL_L_X4Y128_SLICE_X4Y128_AO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A2 = CLBLM_L_X8Y128_SLICE_X11Y128_DQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_B6 = CLBLM_L_X10Y119_SLICE_X13Y119_DO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D1 = CLBLM_R_X7Y116_SLICE_X9Y116_BQ;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A3 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D2 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D3 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D4 = CLBLM_R_X7Y116_SLICE_X8Y116_BO6;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D5 = CLBLM_R_X7Y124_SLICE_X8Y124_B5Q;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y116_SLICE_X9Y116_D6 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B1 = CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_A5 = CLBLM_R_X7Y126_SLICE_X9Y126_BQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A1 = CLBLM_R_X7Y116_SLICE_X8Y116_DO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A2 = CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A3 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_A6 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C5 = CLBLM_L_X10Y125_SLICE_X12Y125_CQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C1 = CLBLM_R_X11Y130_SLICE_X14Y130_BO5;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C2 = CLBLM_R_X11Y126_SLICE_X14Y126_CQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B1 = CLBLL_L_X4Y117_SLICE_X5Y117_BQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B2 = CLBLM_L_X8Y119_SLICE_X11Y119_BQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B3 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B4 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B5 = CLBLM_R_X5Y116_SLICE_X7Y116_CQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_B6 = 1'b1;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D1 = CLBLM_R_X11Y126_SLICE_X15Y126_DO5;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C3 = CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C1 = CLBLM_R_X5Y116_SLICE_X6Y116_AQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C2 = CLBLM_R_X7Y115_SLICE_X8Y115_AO5;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C3 = CLBLM_R_X7Y117_SLICE_X8Y117_DQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C4 = CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C5 = CLBLM_R_X7Y116_SLICE_X8Y116_BO5;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_C6 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C5 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C6 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X12Y117_B1 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_C6 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D1 = CLBLM_R_X7Y118_SLICE_X8Y118_C5Q;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D2 = 1'b1;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D3 = CLBLM_R_X7Y116_SLICE_X8Y116_AQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D4 = CLBLM_R_X7Y119_SLICE_X8Y119_CQ;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D5 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X7Y116_SLICE_X8Y116_D6 = CLBLM_L_X8Y118_SLICE_X11Y118_CO6;
  assign RIOB33_X105Y183_IOB_X1Y184_O = CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  assign RIOB33_X105Y183_IOB_X1Y183_O = CLBLM_L_X10Y126_SLICE_X12Y126_DO5;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A1 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A2 = CLBLM_R_X5Y125_SLICE_X6Y125_A5Q;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A3 = CLBLL_L_X4Y129_SLICE_X4Y129_AQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A5 = CLBLL_L_X4Y125_SLICE_X4Y125_AQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A6 = CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  assign CLBLM_L_X8Y118_SLICE_X11Y118_D6 = CLBLM_L_X8Y116_SLICE_X10Y116_BQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B4 = CLBLL_L_X2Y130_SLICE_X0Y130_CO5;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D1 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C2 = CLBLL_L_X4Y130_SLICE_X4Y130_AO5;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C3 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C4 = CLBLL_L_X2Y130_SLICE_X0Y130_BO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C6 = CLBLL_L_X4Y122_SLICE_X4Y122_AQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D2 = CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D1 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D3 = CLBLL_L_X4Y127_SLICE_X4Y127_DO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D4 = CLBLL_L_X4Y120_SLICE_X5Y120_CQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D5 = CLBLL_L_X4Y129_SLICE_X4Y129_BO5;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D6 = CLBLM_R_X3Y129_SLICE_X3Y129_AO6;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D5 = CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  assign CLBLM_L_X8Y119_SLICE_X11Y119_D6 = CLBLM_L_X8Y117_SLICE_X10Y117_BQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A2 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A4 = CLBLM_L_X8Y123_SLICE_X11Y123_DO5;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A5 = CLBLM_R_X3Y120_SLICE_X2Y120_CQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_A6 = CLBLM_L_X10Y124_SLICE_X13Y124_C5Q;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B1 = CLBLM_L_X8Y123_SLICE_X11Y123_CQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B2 = CLBLM_L_X10Y126_SLICE_X12Y126_CQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B3 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B4 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C1 = CLBLM_L_X8Y123_SLICE_X11Y123_C5Q;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A1 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A2 = CLBLM_R_X7Y129_SLICE_X8Y129_A5Q;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A3 = CLBLL_L_X4Y129_SLICE_X5Y129_AQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A5 = CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C2 = CLBLM_L_X8Y123_SLICE_X10Y123_C5Q;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C4 = CLBLM_L_X10Y127_SLICE_X12Y127_DQ;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A1 = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A3 = CLBLL_L_X2Y119_SLICE_X0Y119_AO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_A6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D1 = CLBLM_L_X10Y126_SLICE_X12Y126_CQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D2 = CLBLM_L_X10Y123_SLICE_X12Y123_BQ;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_B6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A1 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A2 = CLBLL_L_X4Y123_SLICE_X5Y123_BQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A4 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_A6 = CLBLM_R_X7Y120_SLICE_X9Y120_BO6;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_C6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B1 = CLBLM_R_X11Y124_SLICE_X14Y124_CQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B2 = CLBLM_L_X8Y123_SLICE_X10Y123_BQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X0Y115_D6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B6 = CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C1 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C2 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C4 = CLBLM_L_X8Y122_SLICE_X10Y122_BQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_C6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D1 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D2 = CLBLL_L_X2Y121_SLICE_X0Y121_AQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D3 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D5 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_D6 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_A6 = 1'b1;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_D = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_B6 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_C6 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A1 = CLBLM_R_X11Y127_SLICE_X15Y127_BO5;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A2 = CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A4 = CLBLM_R_X11Y127_SLICE_X15Y127_DO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A5 = CLBLM_R_X11Y130_SLICE_X14Y130_BO5;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_A6 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D1 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D2 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D3 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D4 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D5 = 1'b1;
  assign CLBLL_L_X2Y115_SLICE_X1Y115_D6 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B1 = CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B2 = CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B3 = CLBLM_R_X11Y127_SLICE_X15Y127_CO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A1 = CLBLM_R_X7Y118_SLICE_X8Y118_DQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A2 = CLBLM_R_X5Y116_SLICE_X7Y116_CQ;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C2 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A3 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A4 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A5 = CLBLL_L_X4Y117_SLICE_X5Y117_BQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_A6 = 1'b1;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C3 = CLBLM_L_X8Y123_SLICE_X10Y123_CQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C1 = CLBLM_L_X12Y127_SLICE_X17Y127_BO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B1 = CLBLM_L_X8Y117_SLICE_X10Y117_DO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B2 = CLBLM_R_X7Y117_SLICE_X8Y117_CQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B3 = CLBLL_L_X4Y120_SLICE_X4Y120_C5Q;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A1 = CLBLM_L_X8Y118_SLICE_X10Y118_DO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B4 = CLBLM_L_X10Y119_SLICE_X12Y119_CQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B5 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_B6 = CLBLM_R_X7Y117_SLICE_X9Y117_AO5;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D3 = CLBLM_R_X11Y126_SLICE_X14Y126_DQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C1 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C2 = CLBLM_R_X7Y115_SLICE_X9Y115_AO5;
  assign CLBLM_L_X8Y119_SLICE_X10Y119_C6 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C3 = CLBLM_R_X5Y117_SLICE_X6Y117_CQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C4 = CLBLM_R_X7Y117_SLICE_X9Y117_AO5;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C5 = CLBLM_R_X7Y118_SLICE_X8Y118_DQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_C6 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D4 = CLBLM_L_X12Y127_SLICE_X16Y127_CO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A1 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A2 = CLBLM_R_X11Y127_SLICE_X15Y127_AQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A4 = CLBLL_L_X4Y123_SLICE_X5Y123_CO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A5 = CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_A6 = CLBLM_R_X11Y127_SLICE_X14Y127_CO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D1 = CLBLM_R_X5Y117_SLICE_X7Y117_CO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D2 = CLBLM_R_X7Y118_SLICE_X9Y118_DO6;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D3 = CLBLM_R_X5Y116_SLICE_X7Y116_BQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A2 = CLBLM_L_X10Y120_SLICE_X12Y120_AQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D4 = CLBLM_L_X10Y120_SLICE_X13Y120_A5Q;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D5 = CLBLM_L_X10Y121_SLICE_X12Y121_CQ;
  assign CLBLM_R_X7Y117_SLICE_X9Y117_D6 = CLBLM_L_X8Y117_SLICE_X11Y117_CO6;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D2 = CLBLL_L_X4Y122_SLICE_X4Y122_A5Q;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D4 = CLBLM_R_X11Y123_SLICE_X14Y123_DQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B1 = CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B2 = CLBLM_R_X11Y126_SLICE_X15Y126_BQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A1 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A3 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A5 = CLBLM_R_X7Y116_SLICE_X9Y116_AQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_A6 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C1 = CLBLM_L_X10Y124_SLICE_X13Y124_A5Q;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C2 = CLBLM_R_X11Y127_SLICE_X14Y127_BO5;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C3 = CLBLM_R_X11Y127_SLICE_X14Y127_AQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B1 = CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B2 = CLBLM_L_X8Y117_SLICE_X10Y117_CO5;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B4 = CLBLM_R_X7Y126_SLICE_X9Y126_BQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B5 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D5 = CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C2 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C3 = CLBLM_R_X7Y117_SLICE_X9Y117_BO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C4 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C5 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_C6 = CLBLM_R_X7Y123_SLICE_X9Y123_A5Q;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D3 = CLBLM_L_X10Y127_SLICE_X13Y127_DQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D4 = CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D6 = CLBLM_R_X11Y126_SLICE_X15Y126_BQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B5 = CLBLL_L_X4Y125_SLICE_X4Y125_C5Q;
  assign RIOB33_X105Y185_IOB_X1Y185_O = CLBLM_L_X10Y123_SLICE_X13Y123_DO5;
  assign RIOB33_X105Y185_IOB_X1Y186_O = CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_B6 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D2 = CLBLM_R_X7Y116_SLICE_X8Y116_CO6;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D3 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D4 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D5 = 1'b1;
  assign CLBLM_R_X7Y117_SLICE_X8Y117_D6 = CLBLM_R_X3Y122_SLICE_X3Y122_AQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D4 = CLBLM_L_X8Y121_SLICE_X10Y121_BQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_D6 = CLBLM_L_X10Y128_SLICE_X12Y128_BQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A2 = CLBLL_L_X4Y125_SLICE_X4Y125_C5Q;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A3 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A4 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A5 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C3 = CLBLM_R_X3Y123_SLICE_X3Y123_BQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D5 = CLBLM_L_X10Y127_SLICE_X12Y127_CQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B1 = CLBLL_L_X2Y130_SLICE_X0Y130_CO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B2 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B3 = CLBLL_L_X2Y130_SLICE_X0Y130_AO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B4 = CLBLL_L_X2Y130_SLICE_X0Y130_BO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B5 = CLBLL_L_X4Y130_SLICE_X4Y130_AO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B6 = CLBLM_R_X5Y129_SLICE_X6Y129_CQ;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C5 = CLBLM_L_X8Y117_SLICE_X10Y117_AQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C1 = CLBLM_R_X3Y130_SLICE_X3Y130_AO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C2 = CLBLL_L_X4Y130_SLICE_X5Y130_AO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C3 = CLBLM_R_X3Y123_SLICE_X2Y123_AQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C4 = CLBLL_L_X4Y131_SLICE_X4Y131_AO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C5 = CLBLL_L_X4Y127_SLICE_X4Y127_DO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C6 = CLBLL_L_X4Y130_SLICE_X4Y130_BO6;
  assign CLBLL_L_X4Y125_SLICE_X4Y125_C6 = 1'b1;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_A6 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D5 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D2 = CLBLL_L_X4Y125_SLICE_X4Y125_C5Q;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D4 = CLBLM_R_X5Y129_SLICE_X6Y129_CQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D5 = CLBLL_L_X2Y130_SLICE_X0Y130_AO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D6 = CLBLL_L_X2Y130_SLICE_X0Y130_CO6;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_D1 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A2 = CLBLM_L_X8Y126_SLICE_X11Y126_BQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A3 = CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A4 = CLBLM_R_X5Y124_SLICE_X7Y124_CQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_A6 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B2 = CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B4 = CLBLM_L_X8Y123_SLICE_X11Y123_BQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B5 = CLBLM_L_X8Y124_SLICE_X11Y124_CO5;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_B6 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A1 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A2 = CLBLL_L_X2Y130_SLICE_X0Y130_BO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A3 = CLBLL_L_X2Y130_SLICE_X0Y130_AO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A6 = CLBLL_L_X4Y120_SLICE_X5Y120_CQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C1 = CLBLM_L_X8Y123_SLICE_X10Y123_AQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C2 = CLBLM_L_X10Y124_SLICE_X13Y124_BQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C3 = CLBLM_R_X5Y124_SLICE_X6Y124_CQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C6 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_C4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A4 = CLBLL_L_X2Y130_SLICE_X0Y130_CO5;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B1 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B2 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B3 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B4 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B5 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B6 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C1 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C2 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C3 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C4 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C5 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C6 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D3 = CLBLM_R_X3Y123_SLICE_X2Y123_DQ;
  assign CLBLM_L_X8Y124_SLICE_X11Y124_D4 = CLBLM_L_X8Y121_SLICE_X10Y121_DO5;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A2 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D1 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A3 = CLBLM_L_X8Y124_SLICE_X10Y124_AQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A4 = CLBLM_R_X5Y124_SLICE_X7Y124_CQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D2 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D3 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D4 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_A6 = CLBLM_R_X7Y124_SLICE_X9Y124_AQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D6 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B1 = CLBLM_L_X8Y126_SLICE_X11Y126_B5Q;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B2 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B6 = 1'b1;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_B5 = CLBLM_L_X10Y122_SLICE_X13Y122_DQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_D1 = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C1 = CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C2 = CLBLM_R_X7Y124_SLICE_X8Y124_CO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C3 = CLBLM_R_X11Y125_SLICE_X14Y125_CQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C4 = CLBLM_R_X7Y126_SLICE_X9Y126_CQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C5 = CLBLM_L_X10Y124_SLICE_X12Y124_DO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_C6 = CLBLM_R_X7Y124_SLICE_X9Y124_CO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_T1 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_D1 = CLBLM_R_X103Y173_SLICE_X163Y173_AO5;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_D1 = CLBLM_R_X3Y123_SLICE_X3Y123_CQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D1 = CLBLM_L_X8Y124_SLICE_X10Y124_BQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D3 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D4 = CLBLL_L_X4Y124_SLICE_X4Y124_DQ;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D5 = CLBLM_L_X10Y124_SLICE_X12Y124_DO6;
  assign CLBLM_L_X8Y124_SLICE_X10Y124_D6 = CLBLM_R_X7Y124_SLICE_X9Y124_AQ;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_D1 = CLBLM_L_X10Y136_SLICE_X12Y136_BO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A1 = CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A2 = CLBLM_L_X10Y128_SLICE_X13Y128_CO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A4 = CLBLM_R_X11Y129_SLICE_X15Y129_BO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A5 = CLBLM_R_X11Y123_SLICE_X15Y123_AQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_A6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B1 = CLBLM_L_X10Y129_SLICE_X13Y129_CO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B2 = CLBLM_L_X10Y126_SLICE_X13Y126_AQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B3 = CLBLM_R_X11Y126_SLICE_X15Y126_AQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B4 = CLBLM_R_X11Y129_SLICE_X15Y129_DO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B5 = CLBLM_R_X11Y128_SLICE_X14Y128_AO5;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_B6 = CLBLM_R_X11Y129_SLICE_X15Y129_CO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A1 = CLBLM_R_X7Y125_SLICE_X9Y125_DQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A2 = CLBLM_L_X8Y116_SLICE_X10Y116_BQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A3 = CLBLM_R_X7Y118_SLICE_X9Y118_AQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A4 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_A6 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C1 = CLBLM_L_X10Y128_SLICE_X13Y128_BQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_C2 = CLBLM_R_X11Y129_SLICE_X15Y129_CO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B1 = CLBLL_L_X2Y127_SLICE_X0Y127_CO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B2 = CLBLM_R_X7Y128_SLICE_X9Y128_BO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B3 = CLBLL_L_X4Y128_SLICE_X4Y128_AO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B4 = CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B5 = CLBLM_R_X3Y127_SLICE_X2Y127_DO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_B6 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D1 = CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C1 = CLBLM_R_X3Y126_SLICE_X3Y126_AO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C2 = CLBLM_R_X7Y128_SLICE_X9Y128_BO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C3 = CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C4 = CLBLM_R_X3Y128_SLICE_X2Y128_AO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C5 = CLBLL_L_X4Y128_SLICE_X4Y128_AO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_C6 = CLBLM_R_X5Y118_SLICE_X7Y118_BO6;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D3 = CLBLM_L_X12Y127_SLICE_X16Y127_AQ;
  assign CLBLM_R_X11Y128_SLICE_X15Y128_D4 = CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  assign CLBLM_L_X8Y118_SLICE_X10Y118_B3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A1 = CLBLM_R_X11Y129_SLICE_X15Y129_AO5;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A2 = CLBLM_L_X10Y125_SLICE_X13Y125_DO5;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A3 = CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A4 = CLBLM_R_X11Y126_SLICE_X14Y126_BQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D1 = CLBLM_L_X8Y118_SLICE_X11Y118_BQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D2 = CLBLM_L_X8Y118_SLICE_X11Y118_DO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D3 = CLBLM_R_X5Y117_SLICE_X7Y117_BO6;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D4 = CLBLM_R_X3Y119_SLICE_X3Y119_BO5;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D5 = CLBLM_R_X5Y118_SLICE_X7Y118_AQ;
  assign CLBLM_R_X7Y118_SLICE_X9Y118_D6 = CLBLM_L_X10Y121_SLICE_X12Y121_CQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A5 = CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_A6 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_AX = CLBLM_L_X10Y128_SLICE_X13Y128_BQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B1 = CLBLM_L_X10Y129_SLICE_X13Y129_CO6;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B2 = CLBLM_L_X10Y128_SLICE_X12Y128_CQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_B3 = CLBLM_R_X11Y128_SLICE_X14Y128_AO5;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A1 = CLBLM_R_X7Y123_SLICE_X9Y123_A5Q;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A1 = CLBLM_R_X7Y129_SLICE_X8Y129_DQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A2 = CLBLM_R_X7Y118_SLICE_X9Y118_DO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A4 = 1'b1;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A5 = CLBLM_R_X3Y125_SLICE_X2Y125_BO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_A6 = CLBLM_R_X7Y118_SLICE_X8Y118_AQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A3 = CLBLL_L_X4Y125_SLICE_X5Y125_AQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B1 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B2 = CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B4 = CLBLM_R_X5Y119_SLICE_X7Y119_BQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A4 = CLBLM_R_X5Y128_SLICE_X6Y128_A5Q;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_B6 = CLBLL_L_X4Y118_SLICE_X4Y118_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A5 = CLBLL_L_X4Y120_SLICE_X5Y120_AQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C2 = CLBLM_R_X5Y118_SLICE_X7Y118_A5Q;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C3 = CLBLM_R_X7Y116_SLICE_X8Y116_AQ;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_A6 = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C4 = CLBLM_R_X5Y120_SLICE_X7Y120_CO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C5 = CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_C6 = 1'b1;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D3 = CLBLM_R_X11Y129_SLICE_X14Y129_BQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D4 = CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_D6 = CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  assign CLBLM_R_X11Y128_SLICE_X14Y128_SR = CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D2 = 1'b1;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D3 = CLBLM_R_X7Y118_SLICE_X8Y118_DQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D4 = CLBLM_R_X5Y118_SLICE_X7Y118_A5Q;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D5 = CLBLM_R_X7Y119_SLICE_X8Y119_DQ;
  assign CLBLM_R_X7Y118_SLICE_X8Y118_D6 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A2 = CLBLM_R_X7Y129_SLICE_X8Y129_DQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A4 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B4 = CLBLM_R_X7Y123_SLICE_X9Y123_A5Q;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B2 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B3 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B4 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B6 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y125_SLICE_X5Y125_B6 = CLBLM_R_X5Y123_SLICE_X7Y123_BQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C1 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C2 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C3 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C4 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C5 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C6 = 1'b1;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_D = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_D = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D1 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D2 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D3 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D4 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D5 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D6 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A1 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A2 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A3 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A4 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A5 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A6 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B1 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B2 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B3 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B4 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B5 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A1 = CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A3 = CLBLM_L_X8Y125_SLICE_X11Y125_AQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A4 = CLBLM_L_X10Y119_SLICE_X12Y119_BQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A5 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_A6 = CLBLM_R_X7Y126_SLICE_X9Y126_DQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C1 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C2 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C3 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B1 = CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A1 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A2 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B2 = CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B3 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_B6 = CLBLM_L_X8Y127_SLICE_X11Y127_CQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A3 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C1 = CLBLM_R_X7Y119_SLICE_X8Y119_CQ;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A3 = CLBLM_R_X3Y126_SLICE_X3Y126_AO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A4 = CLBLM_R_X3Y127_SLICE_X2Y127_DO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_A6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C2 = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y125_SLICE_X11Y125_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B2 = CLBLL_L_X4Y128_SLICE_X4Y128_AO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B3 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B4 = CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_B6 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C1 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C2 = CLBLM_R_X3Y128_SLICE_X3Y128_BO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C3 = CLBLL_L_X2Y127_SLICE_X0Y127_CO6;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C4 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C5 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_C6 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D1 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D2 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D3 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D4 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D1 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D2 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D3 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D4 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X0Y117_D6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B1 = CLBLM_L_X10Y125_SLICE_X12Y125_DQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B4 = CLBLM_L_X8Y122_SLICE_X10Y122_A5Q;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B5 = CLBLM_R_X7Y118_SLICE_X8Y118_DQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_B6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C2 = CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C3 = CLBLM_L_X10Y125_SLICE_X12Y125_CQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C4 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C5 = CLBLM_L_X8Y125_SLICE_X10Y125_BO5;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D4 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D1 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D3 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D4 = CLBLM_R_X7Y126_SLICE_X9Y126_DQ;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A1 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A2 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A3 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A4 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_A6 = 1'b1;
  assign CLBLM_L_X8Y125_SLICE_X10Y125_D6 = CLBLM_L_X8Y119_SLICE_X10Y119_CO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B1 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B2 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B3 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B4 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_B6 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C1 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C2 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C3 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C4 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_C6 = 1'b1;
  assign LIOB33_X0Y103_IOB_X0Y104_O = CLBLL_L_X2Y117_SLICE_X0Y117_AO5;
  assign LIOB33_X0Y103_IOB_X0Y103_O = CLBLL_L_X2Y125_SLICE_X1Y125_CO6;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D1 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D2 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D3 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D4 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D5 = 1'b1;
  assign CLBLL_L_X2Y117_SLICE_X1Y117_D6 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A1 = CLBLM_L_X8Y129_SLICE_X11Y129_BQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A2 = CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A3 = CLBLM_R_X11Y127_SLICE_X15Y127_CO5;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A4 = CLBLM_R_X11Y126_SLICE_X15Y126_BQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A5 = CLBLM_R_X11Y130_SLICE_X14Y130_AQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_A6 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B1 = CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B2 = CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B3 = CLBLM_R_X11Y127_SLICE_X15Y127_CO5;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B4 = CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B5 = CLBLM_R_X11Y130_SLICE_X14Y130_AQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_B6 = CLBLM_R_X11Y129_SLICE_X15Y129_AO5;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A2 = CLBLM_L_X10Y124_SLICE_X13Y124_DQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A4 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A5 = CLBLM_R_X5Y119_SLICE_X6Y119_BO5;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_A6 = CLBLL_L_X4Y119_SLICE_X5Y119_BQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C1 = CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_C2 = CLBLM_L_X12Y127_SLICE_X16Y127_AQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B1 = CLBLM_L_X8Y118_SLICE_X10Y118_CQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B2 = CLBLM_R_X7Y119_SLICE_X9Y119_BQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B4 = CLBLM_R_X5Y119_SLICE_X7Y119_DO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_B6 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D1 = CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D2 = CLBLM_L_X10Y129_SLICE_X13Y129_BO5;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C1 = CLBLM_L_X8Y118_SLICE_X10Y118_BQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C2 = CLBLM_L_X10Y122_SLICE_X12Y122_AQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C3 = CLBLL_L_X2Y127_SLICE_X0Y127_CO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C4 = CLBLM_R_X7Y128_SLICE_X9Y128_BO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C5 = CLBLM_R_X7Y119_SLICE_X9Y119_DO6;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_C6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D3 = CLBLM_L_X12Y126_SLICE_X16Y126_BQ;
  assign CLBLM_R_X11Y129_SLICE_X15Y129_D4 = CLBLM_L_X10Y128_SLICE_X13Y128_AQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A1 = CLBLM_R_X11Y127_SLICE_X15Y127_BO5;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A2 = CLBLM_R_X11Y130_SLICE_X14Y130_BO5;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A3 = CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A4 = CLBLM_L_X8Y129_SLICE_X11Y129_AQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D1 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D2 = CLBLM_L_X8Y118_SLICE_X10Y118_CQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D3 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D4 = CLBLL_L_X4Y119_SLICE_X5Y119_BQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D5 = CLBLM_R_X3Y119_SLICE_X3Y119_AQ;
  assign CLBLM_R_X7Y119_SLICE_X9Y119_D6 = 1'b1;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_A6 = CLBLM_R_X11Y129_SLICE_X14Y129_CO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B1 = CLBLM_R_X11Y127_SLICE_X15Y127_BO5;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B2 = CLBLM_R_X11Y130_SLICE_X14Y130_BO5;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_B4 = CLBLM_R_X11Y129_SLICE_X14Y129_DO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A1 = CLBLM_R_X7Y123_SLICE_X8Y123_B5Q;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A2 = CLBLM_R_X7Y119_SLICE_X8Y119_BQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A3 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_A6 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C1 = CLBLM_R_X11Y129_SLICE_X14Y129_BQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C2 = CLBLM_R_X11Y128_SLICE_X14Y128_AO5;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_C3 = CLBLM_L_X10Y126_SLICE_X13Y126_BQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B2 = CLBLM_R_X7Y119_SLICE_X8Y119_BQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B3 = CLBLM_R_X5Y119_SLICE_X6Y119_AQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B5 = CLBLM_R_X7Y116_SLICE_X9Y116_BQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_B6 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D1 = CLBLM_R_X11Y129_SLICE_X14Y129_BQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D4 = CLBLM_R_X11Y128_SLICE_X14Y128_AO5;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C1 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C2 = CLBLM_R_X7Y119_SLICE_X8Y119_CQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C4 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C5 = CLBLM_R_X7Y125_SLICE_X8Y125_DQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_C6 = CLBLM_L_X10Y119_SLICE_X12Y119_DQ;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D5 = CLBLM_L_X10Y129_SLICE_X13Y129_CO6;
  assign CLBLM_R_X11Y129_SLICE_X14Y129_D6 = CLBLM_L_X10Y129_SLICE_X13Y129_BO5;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D1 = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D2 = CLBLM_R_X7Y119_SLICE_X8Y119_CQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D3 = CLBLM_R_X7Y119_SLICE_X8Y119_DQ;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D4 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D5 = 1'b1;
  assign CLBLM_R_X7Y119_SLICE_X8Y119_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B4 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A1 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A2 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A3 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A4 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A5 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A6 = 1'b1;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A5 = CLBLM_R_X5Y127_SLICE_X7Y127_B5Q;
  assign CLBLM_L_X10Y128_SLICE_X12Y128_A6 = CLBLM_R_X11Y127_SLICE_X15Y127_CO5;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B1 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B2 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B3 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B4 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B5 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B6 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A1 = CLBLM_L_X8Y126_SLICE_X10Y126_CO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A2 = CLBLM_L_X8Y126_SLICE_X10Y126_BO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A3 = CLBLM_L_X8Y126_SLICE_X11Y126_AQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A4 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C1 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C2 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C3 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B1 = CLBLM_L_X10Y127_SLICE_X13Y127_DQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B2 = CLBLM_R_X11Y127_SLICE_X15Y127_BO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B4 = CLBLM_L_X8Y124_SLICE_X10Y124_BQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B5 = CLBLM_R_X5Y126_SLICE_X7Y126_A5Q;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_B6 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A2 = CLBLM_R_X3Y130_SLICE_X3Y130_BO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A3 = CLBLM_R_X3Y128_SLICE_X2Y128_AO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_A6 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C1 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_C2 = CLBLM_R_X11Y127_SLICE_X15Y127_BO6;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B1 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B2 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A1 = CLBLM_R_X7Y126_SLICE_X9Y126_DQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A2 = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B3 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B4 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B5 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_B6 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D1 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C1 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C2 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C3 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C4 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C5 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_C6 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D3 = CLBLM_L_X8Y126_SLICE_X11Y126_DQ;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D5 = CLBLM_L_X8Y125_SLICE_X11Y125_DO6;
  assign CLBLM_L_X8Y126_SLICE_X11Y126_D6 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A2 = CLBLM_L_X10Y125_SLICE_X12Y125_CQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A3 = CLBLM_L_X8Y125_SLICE_X10Y125_CQ;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D4 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D5 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A4 = CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A5 = CLBLM_L_X10Y124_SLICE_X13Y124_DQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_A6 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D1 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D2 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_AX = CLBLM_R_X5Y118_SLICE_X7Y118_AQ;
  assign CLBLL_L_X2Y118_SLICE_X0Y118_D3 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B1 = CLBLM_R_X7Y119_SLICE_X9Y119_AQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B2 = CLBLM_L_X8Y124_SLICE_X11Y124_BQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B3 = CLBLL_L_X4Y125_SLICE_X4Y125_AQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B4 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B5 = CLBLM_L_X8Y126_SLICE_X10Y126_AO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_B6 = CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C1 = CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C2 = CLBLM_L_X8Y127_SLICE_X10Y127_CQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C3 = CLBLM_L_X8Y127_SLICE_X11Y127_DQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C4 = CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C5 = CLBLM_L_X8Y126_SLICE_X10Y126_DO6;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_C6 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D4 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D6 = 1'b1;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D1 = CLBLM_L_X10Y125_SLICE_X13Y125_AQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D2 = CLBLM_L_X8Y127_SLICE_X10Y127_BQ;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D4 = CLBLM_R_X7Y126_SLICE_X9Y126_DQ;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A1 = CLBLL_L_X2Y118_SLICE_X1Y118_B5Q;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_D6 = CLBLM_L_X10Y127_SLICE_X12Y127_CQ;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A2 = CLBLL_L_X2Y118_SLICE_X1Y118_BQ;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A3 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y126_SLICE_X10Y126_SR = CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A5 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_A6 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B2 = CLBLL_L_X2Y118_SLICE_X1Y118_BQ;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B5 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_B6 = CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_BX = CLBLM_R_X3Y118_SLICE_X2Y118_BO5;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C2 = CLBLL_L_X2Y119_SLICE_X0Y119_CO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C3 = CLBLL_L_X2Y118_SLICE_X1Y118_BQ;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C4 = CLBLM_R_X3Y120_SLICE_X3Y120_CO6;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_C6 = 1'b1;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B6 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D1 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D2 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D3 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D4 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D5 = 1'b1;
  assign CLBLL_L_X2Y118_SLICE_X1Y118_D6 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A2 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A3 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A4 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A5 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_A6 = 1'b1;
  assign RIOB33_X105Y191_IOB_X1Y191_O = CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B2 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B3 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B4 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B5 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_B6 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A1 = CLBLM_L_X8Y122_SLICE_X11Y122_AQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A2 = CLBLM_L_X8Y121_SLICE_X11Y121_DO5;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A3 = CLBLM_R_X3Y126_SLICE_X3Y126_AO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A5 = CLBLM_R_X7Y120_SLICE_X8Y120_AQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_A6 = CLBLM_R_X7Y120_SLICE_X9Y120_CO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C2 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_C3 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B1 = CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B3 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B4 = CLBLM_L_X8Y121_SLICE_X11Y121_DO5;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B5 = CLBLM_R_X5Y124_SLICE_X6Y124_CQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_B6 = CLBLM_R_X7Y120_SLICE_X9Y120_CO6;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D2 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C2 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C3 = CLBLM_R_X3Y123_SLICE_X2Y123_DQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_C6 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D3 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X15Y130_D4 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A1 = CLBLM_R_X11Y129_SLICE_X15Y129_AO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A2 = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A3 = CLBLM_R_X11Y130_SLICE_X14Y130_AQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A4 = CLBLM_R_X11Y130_SLICE_X14Y130_BO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_A6 = CLBLM_R_X11Y127_SLICE_X15Y127_BO5;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D2 = CLBLM_R_X3Y127_SLICE_X2Y127_DO6;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D3 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D4 = CLBLM_R_X11Y122_SLICE_X14Y122_BQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D5 = CLBLM_R_X5Y119_SLICE_X7Y119_BQ;
  assign CLBLM_R_X7Y120_SLICE_X9Y120_D6 = CLBLM_R_X7Y128_SLICE_X9Y128_BO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B1 = CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B2 = CLBLM_L_X8Y129_SLICE_X11Y129_BQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B3 = CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B4 = CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_B5 = CLBLM_R_X11Y126_SLICE_X15Y126_BQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A2 = CLBLM_R_X7Y122_SLICE_X9Y122_DO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A3 = CLBLM_R_X7Y120_SLICE_X8Y120_AQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A4 = CLBLM_R_X7Y120_SLICE_X8Y120_CQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_A6 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C2 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_C3 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B1 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B2 = CLBLM_R_X7Y120_SLICE_X8Y120_BQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B4 = CLBLM_L_X8Y128_SLICE_X11Y128_BQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_B6 = CLBLM_R_X7Y122_SLICE_X8Y122_CO6;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D1 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D2 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C2 = CLBLM_R_X7Y120_SLICE_X8Y120_CQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C3 = CLBLM_R_X7Y128_SLICE_X8Y128_DQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C5 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_C6 = CLBLM_R_X7Y119_SLICE_X8Y119_BQ;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D3 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D4 = 1'b1;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D5 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y130_SLICE_X14Y130_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_T1 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D1 = CLBLM_R_X7Y118_SLICE_X8Y118_BQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D2 = CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D4 = CLBLM_R_X7Y122_SLICE_X8Y122_CO6;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D5 = 1'b1;
  assign CLBLM_R_X7Y120_SLICE_X8Y120_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C4 = CLBLM_L_X10Y125_SLICE_X12Y125_DQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C5 = CLBLM_L_X8Y130_SLICE_X10Y130_DO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C1 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C2 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A1 = CLBLM_R_X7Y123_SLICE_X9Y123_CQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A2 = CLBLM_L_X8Y127_SLICE_X11Y127_BQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A3 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A4 = CLBLM_R_X5Y130_SLICE_X7Y130_DO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_A6 = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C3 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B1 = CLBLM_R_X5Y130_SLICE_X7Y130_DO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A1 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A2 = CLBLM_R_X3Y126_SLICE_X3Y126_AO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A3 = CLBLL_L_X4Y128_SLICE_X4Y128_AO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A4 = CLBLL_L_X2Y119_SLICE_X0Y119_BO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_A6 = CLBLM_R_X5Y120_SLICE_X7Y120_A5Q;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B2 = CLBLM_L_X8Y127_SLICE_X11Y127_BQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C1 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B1 = CLBLL_L_X2Y121_SLICE_X0Y121_BO5;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B2 = CLBLM_R_X3Y119_SLICE_X2Y119_CO5;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B3 = CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B4 = CLBLM_R_X3Y128_SLICE_X2Y128_AO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B5 = CLBLM_R_X3Y128_SLICE_X3Y128_BO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_B6 = LIOB33_X0Y51_IOB_X0Y51_I;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C2 = CLBLM_R_X5Y124_SLICE_X6Y124_A5Q;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C1 = CLBLM_R_X3Y128_SLICE_X3Y128_BO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C2 = CLBLM_R_X3Y126_SLICE_X3Y126_AO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C3 = CLBLL_L_X4Y128_SLICE_X4Y128_AO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C5 = CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_C6 = CLBLL_L_X2Y119_SLICE_X0Y119_DO6;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D1 = CLBLM_R_X7Y127_SLICE_X9Y127_CQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D2 = CLBLM_R_X7Y119_SLICE_X9Y119_AQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D3 = CLBLM_L_X10Y124_SLICE_X12Y124_BO5;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D4 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D6 = CLBLM_R_X7Y127_SLICE_X9Y127_CQ;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y127_SLICE_X11Y127_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D1 = CLBLM_R_X3Y130_SLICE_X3Y130_BO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D2 = CLBLM_R_X3Y127_SLICE_X2Y127_DO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D3 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D4 = CLBLL_L_X2Y127_SLICE_X0Y127_CO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D5 = CLBLM_R_X3Y128_SLICE_X2Y128_AO6;
  assign CLBLL_L_X2Y119_SLICE_X0Y119_D6 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A1 = CLBLM_R_X5Y130_SLICE_X7Y130_DO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A2 = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A3 = CLBLM_L_X8Y127_SLICE_X10Y127_AQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A4 = CLBLM_R_X7Y127_SLICE_X9Y127_CQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_A6 = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B1 = CLBLM_R_X5Y128_SLICE_X7Y128_AQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B2 = CLBLM_L_X8Y127_SLICE_X10Y127_BQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B3 = CLBLM_L_X10Y127_SLICE_X12Y127_CQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B4 = CLBLM_L_X8Y127_SLICE_X10Y127_DO6;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C5 = 1'b1;
  assign LIOB33_X0Y107_IOB_X0Y107_O = CLBLL_L_X2Y115_SLICE_X0Y115_AO5;
  assign LIOB33_X0Y107_IOB_X0Y108_O = CLBLL_L_X2Y117_SLICE_X0Y117_BO5;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C1 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C2 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C4 = CLBLM_L_X8Y127_SLICE_X10Y127_BQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C5 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_D = LIOB33_X0Y73_IOB_X0Y74_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A1 = CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A2 = CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A3 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_A6 = CLBLL_L_X2Y119_SLICE_X1Y119_AQ;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D1 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B1 = CLBLM_R_X3Y119_SLICE_X3Y119_BO5;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B2 = CLBLM_R_X7Y117_SLICE_X9Y117_DO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B3 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B4 = CLBLM_R_X5Y120_SLICE_X7Y120_A5Q;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B5 = CLBLM_R_X3Y119_SLICE_X2Y119_CO5;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D5 = 1'b1;
  assign CLBLM_L_X8Y127_SLICE_X10Y127_D6 = CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C1 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C2 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C3 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_C6 = 1'b1;
  assign RIOB33_X105Y193_IOB_X1Y193_O = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign RIOB33_X105Y193_IOB_X1Y194_O = CLBLM_R_X11Y131_SLICE_X15Y131_AQ;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D1 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D2 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D3 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D4 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D5 = 1'b1;
  assign CLBLL_L_X2Y119_SLICE_X1Y119_D6 = 1'b1;
  assign LIOB33_X0Y119_IOB_X0Y120_O = CLBLM_L_X10Y120_SLICE_X13Y120_AQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A2 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A3 = CLBLM_R_X11Y131_SLICE_X15Y131_AQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A4 = CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A5 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A6 = 1'b1;
  assign LIOB33_X0Y119_IOB_X0Y119_O = CLBLM_L_X8Y122_SLICE_X10Y122_AQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B1 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B2 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B3 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B4 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B5 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A2 = CLBLM_R_X7Y123_SLICE_X8Y123_B5Q;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A3 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A4 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_A6 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C1 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C2 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C3 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B1 = CLBLM_R_X5Y123_SLICE_X6Y123_CQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B2 = CLBLM_R_X7Y125_SLICE_X9Y125_A5Q;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B4 = CLBLM_R_X11Y121_SLICE_X14Y121_AQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_B6 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D1 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C1 = CLBLM_L_X8Y119_SLICE_X10Y119_BQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C2 = CLBLM_R_X5Y120_SLICE_X6Y120_DQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C3 = CLBLM_R_X5Y123_SLICE_X7Y123_CQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C4 = CLBLM_R_X5Y118_SLICE_X6Y118_B5Q;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C5 = CLBLM_R_X7Y116_SLICE_X9Y116_AQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_C6 = CLBLM_L_X8Y123_SLICE_X11Y123_C5Q;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D3 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D4 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A1 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A2 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A3 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A4 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A5 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C2 = CLBLM_R_X7Y128_SLICE_X8Y128_BQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D1 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D2 = CLBLM_R_X5Y121_SLICE_X6Y121_CO5;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D3 = CLBLM_R_X3Y123_SLICE_X2Y123_DQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D4 = CLBLM_L_X8Y118_SLICE_X10Y118_AO5;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C3 = CLBLM_R_X5Y124_SLICE_X7Y124_BQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D5 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_R_X7Y121_SLICE_X9Y121_D6 = CLBLM_R_X5Y118_SLICE_X7Y118_BO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C4 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B1 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B2 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A1 = CLBLM_R_X3Y126_SLICE_X2Y126_A5Q;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A3 = CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A4 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_A6 = CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C6 = CLBLL_L_X2Y130_SLICE_X1Y130_AO6;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_AX = CLBLM_L_X8Y121_SLICE_X10Y121_AO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C1 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B1 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B2 = CLBLM_R_X7Y125_SLICE_X8Y125_BQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B4 = CLBLM_R_X11Y122_SLICE_X14Y122_BQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_B6 = CLBLM_R_X7Y121_SLICE_X8Y121_CO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B3 = CLBLM_L_X8Y123_SLICE_X11Y123_AQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B4 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D1 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C1 = CLBLM_L_X8Y124_SLICE_X10Y124_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C2 = CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C4 = CLBLM_R_X7Y124_SLICE_X8Y124_CO5;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C5 = CLBLM_L_X8Y122_SLICE_X11Y122_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_C6 = CLBLM_R_X5Y120_SLICE_X6Y120_DQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B5 = CLBLM_R_X5Y126_SLICE_X7Y126_CO5;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D6 = 1'b1;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D1 = CLBLM_L_X8Y124_SLICE_X10Y124_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D2 = CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D3 = CLBLL_L_X4Y122_SLICE_X5Y122_DQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D5 = CLBLM_R_X7Y127_SLICE_X8Y127_CQ;
  assign CLBLM_R_X7Y121_SLICE_X8Y121_D6 = CLBLM_R_X7Y124_SLICE_X8Y124_CO5;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D1 = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D2 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D3 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C4 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D5 = CLBLM_R_X7Y128_SLICE_X8Y128_CQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D6 = CLBLL_L_X2Y130_SLICE_X1Y130_AO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C6 = CLBLM_R_X5Y126_SLICE_X7Y126_CO5;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D4 = CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D5 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A1 = CLBLM_L_X8Y128_SLICE_X11Y128_AQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A2 = CLBLM_R_X5Y130_SLICE_X7Y130_DO6;
  assign CLBLM_L_X8Y120_SLICE_X11Y120_D6 = CLBLM_R_X11Y122_SLICE_X15Y122_AQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A3 = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A5 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_A6 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_A6 = CLBLM_R_X5Y128_SLICE_X6Y128_DQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_B6 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B4 = CLBLM_R_X7Y128_SLICE_X9Y128_AQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_B5 = CLBLM_R_X5Y130_SLICE_X7Y130_DO6;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_C6 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C4 = CLBLM_L_X8Y125_SLICE_X11Y125_CQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C5 = CLBLM_R_X7Y131_SLICE_X9Y131_BO6;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D2 = CLBLM_L_X8Y127_SLICE_X11Y127_DQ;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D1 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X0Y120_D6 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X11Y128_D6 = CLBLM_L_X8Y127_SLICE_X11Y127_CQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A1 = CLBLM_L_X8Y129_SLICE_X10Y129_CO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A2 = CLBLL_L_X2Y121_SLICE_X0Y121_AQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A4 = CLBLM_R_X7Y131_SLICE_X9Y131_BO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A5 = CLBLM_R_X7Y131_SLICE_X8Y131_CO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_A6 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B1 = CLBLM_L_X8Y128_SLICE_X10Y128_DO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B2 = CLBLM_R_X7Y131_SLICE_X9Y131_BO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B3 = CLBLL_L_X4Y120_SLICE_X5Y120_BQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B5 = CLBLM_R_X7Y131_SLICE_X8Y131_CO6;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_B6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOB33_X105Y195_IOB_X1Y196_O = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C2 = CLBLM_L_X8Y128_SLICE_X10Y128_CQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C4 = CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C5 = CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A1 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A3 = CLBLM_L_X10Y118_SLICE_X13Y118_AQ;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A5 = CLBLL_L_X4Y126_SLICE_X4Y126_AQ;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_A6 = CLBLL_L_X2Y121_SLICE_X0Y121_A5Q;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B1 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B3 = CLBLL_L_X4Y126_SLICE_X4Y126_AQ;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B5 = CLBLL_L_X2Y121_SLICE_X1Y121_B5Q;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_B6 = CLBLL_L_X2Y121_SLICE_X0Y121_A5Q;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D1 = CLBLM_L_X8Y127_SLICE_X11Y127_BQ;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D2 = 1'b1;
  assign CLBLM_L_X8Y128_SLICE_X10Y128_D3 = CLBLM_L_X8Y128_SLICE_X10Y128_BQ;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_C6 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C2 = CLBLL_L_X4Y124_SLICE_X5Y124_CQ;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_T1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D1 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D2 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D3 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D4 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D5 = 1'b1;
  assign CLBLL_L_X2Y120_SLICE_X1Y120_D6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C2 = CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C4 = CLBLM_R_X5Y128_SLICE_X6Y128_A5Q;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C3 = CLBLM_R_X5Y126_SLICE_X7Y126_CO5;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C5 = CLBLM_R_X7Y128_SLICE_X9Y128_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C6 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A1 = CLBLM_R_X7Y117_SLICE_X8Y117_CQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A2 = CLBLM_L_X8Y123_SLICE_X10Y123_BQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A3 = CLBLM_R_X7Y122_SLICE_X9Y122_AQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_A6 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C4 = CLBLM_R_X3Y124_SLICE_X3Y124_BQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B2 = CLBLM_L_X8Y123_SLICE_X10Y123_BQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B3 = CLBLM_R_X7Y121_SLICE_X9Y121_AQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B4 = CLBLM_L_X8Y122_SLICE_X10Y122_BO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_B6 = CLBLM_L_X10Y122_SLICE_X12Y122_AQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C2 = CLBLM_L_X8Y122_SLICE_X10Y122_BO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C3 = CLBLM_R_X5Y128_SLICE_X7Y128_B5Q;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C4 = CLBLM_L_X10Y122_SLICE_X12Y122_AQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C5 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X103Y171_SLICE_X162Y171_D3 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y171_SLICE_X162Y171_D4 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C5 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D1 = CLBLM_L_X8Y124_SLICE_X10Y124_AQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D2 = CLBLM_R_X7Y124_SLICE_X8Y124_CO6;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D4 = CLBLM_L_X10Y126_SLICE_X12Y126_CQ;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D5 = CLBLM_L_X8Y123_SLICE_X11Y123_C5Q;
  assign CLBLM_R_X7Y122_SLICE_X9Y122_D6 = CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  assign CLBLM_R_X103Y171_SLICE_X162Y171_D5 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X162Y171_D6 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A2 = CLBLM_R_X11Y122_SLICE_X15Y122_AQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A3 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A4 = CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D2 = CLBLL_L_X2Y120_SLICE_X1Y120_BO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A5 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_A6 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X5Y124_C6 = CLBLM_R_X5Y124_SLICE_X6Y124_A5Q;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B1 = CLBLM_R_X7Y123_SLICE_X8Y123_DO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B2 = CLBLM_R_X5Y125_SLICE_X6Y125_BQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B4 = 1'b1;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_B6 = CLBLM_R_X7Y119_SLICE_X9Y119_CO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D5 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C1 = CLBLM_L_X8Y124_SLICE_X10Y124_AQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C2 = CLBLM_R_X7Y124_SLICE_X8Y124_CO6;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C3 = CLBLM_R_X5Y124_SLICE_X6Y124_CQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C5 = CLBLM_R_X5Y123_SLICE_X7Y123_CQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_C6 = CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D1 = CLBLM_L_X8Y124_SLICE_X10Y124_AQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D2 = CLBLL_L_X4Y124_SLICE_X4Y124_DQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D3 = CLBLM_L_X8Y121_SLICE_X11Y121_CQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D4 = CLBLM_R_X3Y122_SLICE_X2Y122_A5Q;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D5 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign CLBLM_R_X7Y122_SLICE_X8Y122_D6 = CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_D1 = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = CLBLM_R_X3Y132_SLICE_X2Y132_BQ;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_D1 = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_D1 = CLBLM_R_X11Y124_SLICE_X14Y124_DO6;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_D1 = CLBLM_R_X3Y129_SLICE_X2Y129_AQ;
  assign LIOB33_X0Y111_IOB_X0Y112_O = CLBLM_L_X10Y121_SLICE_X13Y121_B5Q;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A1 = CLBLM_L_X8Y129_SLICE_X11Y129_DO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A1 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A2 = CLBLM_R_X5Y127_SLICE_X7Y127_BQ;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A3 = CLBLL_L_X2Y121_SLICE_X0Y121_AQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A5 = CLBLM_R_X7Y131_SLICE_X8Y131_CO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A6 = CLBLM_R_X7Y123_SLICE_X9Y123_BQ;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A4 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A2 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_AX = CLBLL_L_X2Y121_SLICE_X0Y121_BO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B4 = CLBLM_L_X10Y128_SLICE_X13Y128_DO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B5 = CLBLM_R_X5Y129_SLICE_X7Y129_BO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_B6 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B3 = CLBLL_L_X4Y126_SLICE_X4Y126_AQ;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B4 = CLBLL_L_X4Y121_SLICE_X5Y121_BQ;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B5 = CLBLL_L_X2Y121_SLICE_X0Y121_A5Q;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_B6 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_BX = CLBLL_L_X2Y121_SLICE_X1Y121_AO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C2 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C6 = CLBLM_R_X7Y131_SLICE_X9Y131_CO6;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C3 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C4 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_C6 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C3 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C4 = CLBLM_R_X7Y128_SLICE_X9Y128_DO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_C5 = CLBLM_L_X8Y129_SLICE_X10Y129_AO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D1 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D2 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D3 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D5 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D6 = CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D4 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X0Y121_D6 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D4 = CLBLM_R_X7Y131_SLICE_X9Y131_CO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A1 = CLBLM_R_X7Y130_SLICE_X9Y130_CO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A2 = CLBLM_L_X8Y128_SLICE_X10Y128_BQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A3 = CLBLM_L_X8Y128_SLICE_X10Y128_AQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A4 = CLBLM_R_X7Y129_SLICE_X9Y129_AQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A5 = CLBLM_L_X8Y129_SLICE_X11Y129_AQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1 = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_AX = CLBLM_R_X5Y124_SLICE_X6Y124_A5Q;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B1 = CLBLM_R_X7Y131_SLICE_X9Y131_CO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B2 = CLBLM_R_X7Y128_SLICE_X9Y128_DO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B3 = CLBLM_L_X8Y128_SLICE_X10Y128_AQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B4 = CLBLM_L_X8Y128_SLICE_X11Y128_AQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B5 = CLBLM_L_X8Y129_SLICE_X11Y129_AQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_B6 = CLBLM_R_X7Y130_SLICE_X9Y130_CO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C1 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A1 = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A3 = CLBLL_L_X4Y123_SLICE_X5Y123_B5Q;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C5 = CLBLM_L_X8Y128_SLICE_X10Y128_AQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C6 = CLBLM_L_X8Y129_SLICE_X11Y129_AQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A4 = CLBLL_L_X2Y121_SLICE_X0Y121_BQ;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A5 = CLBLL_L_X2Y121_SLICE_X1Y121_CO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_A6 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C2 = CLBLM_R_X7Y128_SLICE_X9Y128_DO6;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_C3 = CLBLM_R_X7Y130_SLICE_X9Y130_CO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B1 = CLBLM_R_X3Y122_SLICE_X2Y122_A5Q;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B3 = CLBLL_L_X2Y120_SLICE_X1Y120_AQ;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B4 = CLBLL_L_X2Y122_SLICE_X1Y122_BQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D2 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B5 = CLBLL_L_X4Y123_SLICE_X5Y123_AQ;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_B6 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D1 = CLBLM_L_X8Y129_SLICE_X11Y129_AQ;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C1 = CLBLM_R_X5Y127_SLICE_X7Y127_BQ;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C3 = CLBLL_L_X4Y120_SLICE_X4Y120_CQ;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C4 = CLBLM_R_X3Y123_SLICE_X3Y123_CQ;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_C6 = CLBLM_R_X3Y121_SLICE_X2Y121_CQ;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D6 = CLBLM_R_X7Y129_SLICE_X9Y129_AQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_SR = CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D1 = CLBLM_R_X5Y127_SLICE_X7Y127_BQ;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D2 = CLBLM_R_X3Y123_SLICE_X3Y123_CQ;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D4 = CLBLL_L_X4Y120_SLICE_X4Y120_CQ;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D5 = 1'b1;
  assign CLBLL_L_X2Y121_SLICE_X1Y121_D6 = CLBLM_R_X3Y121_SLICE_X2Y121_CQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A1 = CLBLM_R_X7Y123_SLICE_X9Y123_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A3 = CLBLL_L_X4Y121_SLICE_X5Y121_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A4 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_A6 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B1 = CLBLM_L_X10Y120_SLICE_X13Y120_CQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B2 = CLBLM_R_X7Y123_SLICE_X9Y123_BQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B4 = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B5 = CLBLL_L_X4Y120_SLICE_X5Y120_BQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_B6 = CLBLM_R_X7Y123_SLICE_X9Y123_A5Q;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C2 = CLBLM_R_X7Y123_SLICE_X9Y123_CQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C3 = CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C4 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C5 = CLBLM_R_X7Y121_SLICE_X9Y121_DO6;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_C6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D1 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D2 = CLBLL_L_X4Y124_SLICE_X4Y124_DQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D3 = CLBLM_L_X8Y124_SLICE_X10Y124_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D4 = CLBLM_R_X7Y123_SLICE_X9Y123_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D5 = CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  assign CLBLM_R_X7Y123_SLICE_X9Y123_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1 = CLBLM_R_X5Y118_SLICE_X6Y118_AO5;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_D = LIOB33_X0Y75_IOB_X0Y76_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A1 = CLBLM_R_X5Y122_SLICE_X6Y122_CQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A3 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A4 = CLBLM_R_X5Y124_SLICE_X7Y124_CQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_A6 = 1'b1;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_D = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A1 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B1 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B2 = CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B4 = CLBLM_R_X5Y123_SLICE_X6Y123_BQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B5 = CLBLM_R_X3Y121_SLICE_X2Y121_AQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_B6 = 1'b1;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_D = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_D = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C1 = CLBLM_L_X8Y120_SLICE_X10Y120_AQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C2 = CLBLL_L_X4Y122_SLICE_X4Y122_DQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C4 = CLBLM_R_X7Y123_SLICE_X9Y123_CQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_C6 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A2 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D1 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D2 = CLBLM_R_X5Y124_SLICE_X6Y124_A5Q;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D3 = CLBLM_R_X11Y126_SLICE_X14Y126_AQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D4 = 1'b1;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D5 = CLBLM_L_X8Y127_SLICE_X11Y127_CQ;
  assign CLBLM_R_X7Y123_SLICE_X8Y123_D6 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A3 = CLBLM_L_X10Y124_SLICE_X12Y124_AQ;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_B6 = CLBLL_L_X4Y126_SLICE_X4Y126_BO5;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A4 = 1'b1;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C1 = CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  assign LIOB33_X0Y113_IOB_X0Y114_O = CLBLL_L_X4Y118_SLICE_X5Y118_CQ;
  assign LIOB33_X0Y113_IOB_X0Y113_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_D = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLL_L_X4Y126_SLICE_X5Y126_C6 = CLBLM_R_X3Y130_SLICE_X3Y130_AO6;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A1 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A2 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A3 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A4 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A5 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_A6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A1 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A2 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B1 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B2 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B3 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B2 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B4 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B5 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_B6 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C1 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C2 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C3 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C4 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C5 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_C6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B6 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C2 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C4 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D1 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D2 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D3 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D4 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D5 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X0Y122_D6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D1 = CLBLM_L_X8Y130_SLICE_X11Y130_AO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D2 = CLBLM_R_X7Y129_SLICE_X8Y129_CQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D3 = CLBLM_L_X8Y130_SLICE_X11Y130_CO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D4 = CLBLM_L_X8Y130_SLICE_X11Y130_AO5;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D5 = CLBLM_R_X7Y125_SLICE_X8Y125_AQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D6 = CLBLM_L_X8Y130_SLICE_X11Y130_BO6;
  assign LIOB33_X0Y191_IOB_X0Y191_O = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOB33_X105Y195_IOB_X1Y195_O = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A1 = CLBLM_L_X8Y130_SLICE_X10Y130_CQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A3 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A5 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A6 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLM_L_X10Y129_SLICE_X13Y129_A2 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B1 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B2 = CLBLM_R_X7Y131_SLICE_X9Y131_BO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B4 = CLBLM_L_X10Y124_SLICE_X13Y124_A5Q;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B5 = CLBLM_R_X7Y131_SLICE_X8Y131_CO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B6 = CLBLM_L_X8Y131_SLICE_X10Y131_CO6;
  assign RIOB33_X105Y173_IOB_X1Y174_O = CLBLM_R_X103Y173_SLICE_X163Y173_AO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A1 = CLBLL_L_X4Y123_SLICE_X4Y123_BQ;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A2 = CLBLM_R_X3Y120_SLICE_X2Y120_AQ;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A3 = CLBLL_L_X2Y122_SLICE_X1Y122_AQ;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A5 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_A6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C1 = CLBLM_R_X7Y131_SLICE_X8Y131_CO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C6 = CLBLM_R_X7Y131_SLICE_X9Y131_BO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C2 = CLBLM_L_X8Y130_SLICE_X10Y130_CQ;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B2 = CLBLL_L_X2Y122_SLICE_X1Y122_BQ;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B3 = CLBLM_R_X3Y121_SLICE_X3Y121_AQ;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B4 = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B5 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_B6 = CLBLM_R_X7Y123_SLICE_X9Y123_A5Q;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C1 = CLBLL_L_X2Y122_SLICE_X1Y122_A5Q;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C2 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C3 = CLBLL_L_X4Y123_SLICE_X5Y123_B5Q;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C4 = CLBLM_R_X3Y125_SLICE_X2Y125_CO6;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C5 = CLBLM_R_X3Y126_SLICE_X2Y126_A5Q;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_C6 = CLBLM_R_X5Y125_SLICE_X6Y125_A5Q;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D1 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D2 = CLBLM_R_X7Y128_SLICE_X9Y128_DO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D3 = CLBLM_L_X8Y131_SLICE_X10Y131_BO5;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D4 = CLBLM_R_X7Y131_SLICE_X9Y131_CO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D5 = CLBLM_L_X8Y131_SLICE_X10Y131_AO5;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D1 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D2 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D3 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D4 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D5 = 1'b1;
  assign CLBLL_L_X2Y122_SLICE_X1Y122_D6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C3 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A1 = CLBLM_R_X7Y120_SLICE_X8Y120_DQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A2 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A4 = CLBLM_R_X7Y124_SLICE_X9Y124_AQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_A6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C6 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B1 = CLBLM_R_X3Y123_SLICE_X3Y123_AQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B2 = CLBLM_R_X3Y128_SLICE_X2Y128_AO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B4 = CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B5 = CLBLM_L_X10Y123_SLICE_X13Y123_AQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_B6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D2 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C1 = CLBLM_R_X7Y121_SLICE_X9Y121_CO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C2 = CLBLM_R_X7Y124_SLICE_X9Y124_AQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C3 = CLBLM_R_X7Y123_SLICE_X9Y123_AQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C4 = CLBLM_R_X7Y127_SLICE_X8Y127_CQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C5 = CLBLM_R_X7Y124_SLICE_X9Y124_DO6;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_C6 = CLBLM_R_X11Y125_SLICE_X14Y125_CQ;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D6 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D1 = CLBLM_R_X11Y124_SLICE_X14Y124_AQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D2 = CLBLM_L_X8Y121_SLICE_X11Y121_CQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D3 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D4 = CLBLM_R_X7Y129_SLICE_X9Y129_DQ;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D5 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X9Y124_D6 = CLBLM_R_X3Y120_SLICE_X2Y120_BQ;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B3 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A1 = CLBLM_R_X3Y124_SLICE_X2Y124_B5Q;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A3 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A5 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_A6 = CLBLM_R_X7Y116_SLICE_X8Y116_AQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B1 = CLBLM_L_X8Y128_SLICE_X10Y128_AQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B2 = CLBLM_R_X3Y125_SLICE_X3Y125_BQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B3 = CLBLM_L_X10Y124_SLICE_X13Y124_A5Q;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B4 = CLBLM_R_X7Y121_SLICE_X8Y121_A5Q;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_B6 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C1 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C2 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C3 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C4 = CLBLL_L_X4Y124_SLICE_X4Y124_DQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C5 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_C6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B4 = 1'b1;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D1 = CLBLM_L_X8Y124_SLICE_X10Y124_AQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D2 = CLBLM_R_X7Y129_SLICE_X9Y129_DQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D3 = CLBLM_R_X7Y124_SLICE_X8Y124_CO5;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D5 = CLBLL_L_X4Y122_SLICE_X4Y122_DQ;
  assign CLBLM_R_X7Y124_SLICE_X8Y124_D6 = CLBLM_L_X8Y124_SLICE_X11Y124_AQ;
  assign LIOB33_X0Y115_IOB_X0Y116_O = CLBLM_R_X5Y128_SLICE_X7Y128_BQ;
  assign LIOB33_X0Y115_IOB_X0Y115_O = CLBLM_L_X10Y121_SLICE_X13Y121_BQ;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A1 = CLBLM_R_X7Y131_SLICE_X9Y131_BO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A2 = CLBLM_R_X7Y131_SLICE_X8Y131_CO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A4 = CLBLM_R_X11Y130_SLICE_X14Y130_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A5 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A6 = CLBLM_L_X8Y131_SLICE_X11Y131_CO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B1 = CLBLM_L_X8Y129_SLICE_X10Y129_AO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B2 = CLBLM_L_X8Y128_SLICE_X11Y128_CQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B3 = CLBLM_R_X7Y128_SLICE_X9Y128_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B4 = CLBLM_R_X7Y131_SLICE_X9Y131_CO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B5 = CLBLM_R_X7Y128_SLICE_X9Y128_DO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B6 = CLBLM_L_X8Y129_SLICE_X10Y129_AO5;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C1 = CLBLM_R_X7Y128_SLICE_X9Y128_DO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C2 = CLBLM_L_X8Y131_SLICE_X10Y131_AO5;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C3 = CLBLM_L_X8Y131_SLICE_X10Y131_BO5;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C4 = CLBLM_L_X8Y128_SLICE_X11Y128_BQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C5 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C6 = CLBLM_R_X7Y131_SLICE_X9Y131_CO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D3 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D4 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D5 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A1 = CLBLM_L_X8Y129_SLICE_X10Y129_AO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A2 = CLBLM_L_X8Y128_SLICE_X11Y128_CQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A3 = CLBLM_L_X8Y130_SLICE_X10Y130_CQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A4 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A5 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A6 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_T1 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_AX = CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B1 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B2 = CLBLM_L_X8Y128_SLICE_X11Y128_CQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B3 = CLBLM_L_X8Y130_SLICE_X10Y130_CQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B4 = CLBLM_L_X8Y129_SLICE_X10Y129_AO5;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B5 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C1 = CLBLM_L_X8Y131_SLICE_X10Y131_AO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C2 = CLBLM_L_X8Y131_SLICE_X10Y131_BO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C3 = CLBLM_R_X7Y128_SLICE_X9Y128_DO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C4 = CLBLM_L_X8Y127_SLICE_X10Y127_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C5 = CLBLM_R_X7Y131_SLICE_X9Y131_CO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C6 = CLBLM_L_X8Y130_SLICE_X10Y130_BQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D1 = CLBLM_L_X8Y130_SLICE_X10Y130_BQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D2 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D3 = CLBLM_R_X7Y128_SLICE_X9Y128_DO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D4 = CLBLM_L_X8Y131_SLICE_X10Y131_AO5;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D5 = CLBLM_L_X8Y130_SLICE_X10Y130_CQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D6 = CLBLM_L_X8Y131_SLICE_X10Y131_BO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = CLBLL_L_X2Y125_SLICE_X1Y125_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_SR = CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_D1 = CLBLM_L_X10Y123_SLICE_X13Y123_DO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_C6 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_T1 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_D1 = CLBLM_L_X10Y126_SLICE_X12Y126_DO5;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_SING_X0Y150_IOB_X0Y150_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_T1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A3 = CLBLM_R_X7Y125_SLICE_X9Y125_AQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A4 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A5 = CLBLM_R_X7Y120_SLICE_X9Y120_BO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_A6 = CLBLM_R_X5Y126_SLICE_X7Y126_AQ;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_AX = CLBLM_L_X8Y125_SLICE_X10Y125_BO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B1 = CLBLM_R_X3Y123_SLICE_X3Y123_AQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B2 = CLBLM_R_X7Y125_SLICE_X9Y125_BQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B3 = CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B4 = CLBLM_L_X10Y126_SLICE_X12Y126_AQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_B6 = CLBLL_L_X4Y125_SLICE_X4Y125_BQ;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_BX = CLBLM_R_X7Y127_SLICE_X9Y127_DO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C1 = CLBLM_R_X7Y123_SLICE_X8Y123_AQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C2 = CLBLM_R_X7Y125_SLICE_X9Y125_CQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D2 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C3 = CLBLM_L_X10Y125_SLICE_X12Y125_CQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C4 = CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_C6 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D3 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C4 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C5 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_C6 = 1'b1;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D4 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D1 = CLBLM_L_X8Y123_SLICE_X10Y123_CQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D2 = CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D5 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D3 = CLBLM_R_X7Y125_SLICE_X9Y125_DQ;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D4 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y125_SLICE_X9Y125_D6 = CLBLM_L_X10Y127_SLICE_X12Y127_CQ;
  assign CLBLM_L_X10Y129_SLICE_X12Y129_D6 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A1 = CLBLL_L_X4Y120_SLICE_X5Y120_AQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A2 = CLBLM_R_X11Y125_SLICE_X14Y125_CQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A3 = CLBLM_R_X7Y125_SLICE_X8Y125_AQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A5 = CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_A6 = CLBLL_L_X4Y125_SLICE_X4Y125_BQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B1 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B3 = CLBLM_R_X7Y126_SLICE_X8Y126_AQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B4 = CLBLL_L_X4Y122_SLICE_X4Y122_BQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_B6 = CLBLM_R_X7Y124_SLICE_X8Y124_DO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C1 = CLBLM_R_X7Y123_SLICE_X8Y123_CO5;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C2 = CLBLM_R_X7Y125_SLICE_X9Y125_AQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C4 = 1'b1;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C5 = CLBLM_L_X8Y127_SLICE_X11Y127_DQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOB33_X0Y117_IOB_X0Y117_O = CLBLL_L_X2Y122_SLICE_X1Y122_AQ;
  assign LIOB33_X0Y117_IOB_X0Y118_O = CLBLL_L_X4Y122_SLICE_X5Y122_CQ;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D1 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D2 = CLBLM_R_X7Y127_SLICE_X8Y127_CQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D3 = CLBLM_R_X7Y125_SLICE_X8Y125_DQ;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D4 = CLBLM_R_X11Y120_SLICE_X14Y120_DO6;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y125_SLICE_X8Y125_D6 = CLBLM_R_X7Y123_SLICE_X9Y123_A5Q;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D5 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X15Y125_D6 = 1'b1;
  assign LIOB33_SING_X0Y199_IOB_X0Y199_O = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_D = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_D = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_D = RIOB33_X105Y123_IOB_X1Y124_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_D = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C4 = CLBLM_R_X5Y130_SLICE_X7Y130_DO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C5 = CLBLM_R_X7Y127_SLICE_X8Y127_DQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C6 = CLBLM_L_X8Y128_SLICE_X11Y128_BQ;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_B6 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_D = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_R_X103Y171_SLICE_X163Y171_A1 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_R_X103Y171_SLICE_X163Y171_A2 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X163Y171_A3 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X163Y171_A4 = CLBLM_L_X8Y129_SLICE_X10Y129_AQ;
  assign CLBLM_R_X103Y171_SLICE_X163Y171_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y171_SLICE_X163Y171_A6 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X163Y171_B1 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y171_SLICE_X163Y171_B2 = CLBLM_L_X12Y126_SLICE_X16Y126_AQ;
  assign CLBLM_R_X103Y171_SLICE_X163Y171_B3 = CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  assign CLBLM_R_X103Y171_SLICE_X163Y171_B4 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X163Y171_B5 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X163Y171_B6 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D2 = CLBLM_L_X8Y122_SLICE_X11Y122_AQ;
  assign CLBLM_R_X103Y171_SLICE_X163Y171_C1 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X163Y171_C2 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X163Y171_C3 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X163Y171_C4 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X163Y171_C5 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X163Y171_C6 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C5 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X163Y171_D1 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X163Y171_D2 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D6 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X163Y171_D3 = 1'b1;
  assign CLBLM_R_X11Y125_SLICE_X14Y125_C6 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X163Y171_D4 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X163Y171_D5 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X163Y171_D6 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X162Y171_A1 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X162Y171_A2 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X162Y171_A3 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X162Y171_A4 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X162Y171_A5 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X162Y171_A6 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X162Y171_B1 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X162Y171_B2 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X162Y171_B3 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X162Y171_B4 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X162Y171_B5 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X162Y171_B6 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X162Y171_C1 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X162Y171_C2 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X162Y171_C3 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A2 = CLBLM_R_X7Y129_SLICE_X9Y129_BQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A3 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A5 = CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_A6 = CLBLM_R_X7Y127_SLICE_X9Y127_DO5;
  assign CLBLM_R_X103Y171_SLICE_X162Y171_C4 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X162Y171_C5 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X162Y171_C6 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B2 = CLBLM_L_X10Y129_SLICE_X12Y129_BQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B3 = CLBLM_R_X7Y130_SLICE_X9Y130_AQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B4 = CLBLM_L_X10Y124_SLICE_X13Y124_DQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B5 = CLBLM_R_X7Y116_SLICE_X9Y116_BQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_B6 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X162Y171_D1 = 1'b1;
  assign CLBLM_R_X103Y171_SLICE_X162Y171_D2 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A1 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A2 = CLBLM_R_X7Y117_SLICE_X8Y117_CQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A3 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A4 = CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_A6 = CLBLM_R_X7Y118_SLICE_X8Y118_AQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C2 = CLBLM_R_X7Y126_SLICE_X9Y126_CQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B1 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B2 = CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B3 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B5 = CLBLL_L_X4Y123_SLICE_X5Y123_AQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_B6 = CLBLM_R_X5Y116_SLICE_X7Y116_BQ;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C1 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C1 = CLBLM_R_X5Y116_SLICE_X6Y116_AQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C2 = CLBLM_R_X5Y116_SLICE_X7Y116_CQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C4 = CLBLM_R_X7Y126_SLICE_X9Y126_BQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C5 = CLBLM_R_X5Y116_SLICE_X7Y116_DO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y126_SLICE_X9Y126_D6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A1 = CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A2 = CLBLM_L_X8Y126_SLICE_X11Y126_DQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A3 = CLBLM_R_X7Y126_SLICE_X8Y126_AQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A5 = CLBLM_R_X7Y126_SLICE_X9Y126_AQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D1 = CLBLM_L_X10Y117_SLICE_X12Y117_AQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D2 = CLBLM_R_X5Y116_SLICE_X7Y116_CQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D3 = CLBLL_L_X4Y117_SLICE_X5Y117_BQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D4 = CLBLM_R_X7Y117_SLICE_X8Y117_BQ;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D5 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X5Y116_SLICE_X7Y116_D6 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C5 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_A6 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C6 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B1 = CLBLM_R_X7Y124_SLICE_X8Y124_B5Q;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_B2 = CLBLM_R_X7Y126_SLICE_X8Y126_BQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A1 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A2 = CLBLM_R_X5Y128_SLICE_X7Y128_BQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A3 = CLBLM_R_X5Y116_SLICE_X6Y116_AQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A4 = CLBLM_L_X8Y119_SLICE_X11Y119_BQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_A6 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C1 = CLBLM_L_X8Y123_SLICE_X11Y123_AQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C2 = CLBLM_R_X7Y126_SLICE_X8Y126_CQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_C3 = CLBLM_R_X11Y126_SLICE_X14Y126_AQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B1 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B2 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B3 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B4 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B5 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_B6 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D2 = CLBLM_L_X8Y128_SLICE_X11Y128_DQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C1 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C2 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C3 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C4 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C5 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_C6 = 1'b1;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D3 = CLBLM_R_X7Y120_SLICE_X8Y120_DQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D4 = CLBLM_L_X8Y127_SLICE_X11Y127_CQ;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D5 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y126_SLICE_X8Y126_D6 = CLBLM_L_X8Y126_SLICE_X10Y126_AO5;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_A1 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_A2 = CLBLM_R_X5Y123_SLICE_X6Y123_BQ;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D3 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D4 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D5 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D6 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_A3 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_A5 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_A6 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_B1 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_B2 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_B3 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_B4 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_B5 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_B6 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D2 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_C1 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_C2 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_C3 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_C4 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_C5 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_C6 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C4 = CLBLM_R_X7Y128_SLICE_X8Y128_CQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D5 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C5 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D6 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_D1 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_D2 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_D3 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_D4 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_D5 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X54Y124_D6 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_D1 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A1 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A2 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A3 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A4 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A5 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_A6 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B1 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B2 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B3 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B4 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B5 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_B6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D2 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D3 = CLBLM_L_X8Y121_SLICE_X10Y121_DO6;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C1 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C2 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C3 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C4 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C5 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_C6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X11Y121_D4 = CLBLL_L_X4Y128_SLICE_X4Y128_AO6;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_A1 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_A2 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_A3 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_A4 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_A5 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_A6 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D1 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D2 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D3 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D4 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D5 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X0Y125_D6 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_B1 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_B2 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_B3 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_B4 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_B5 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_B6 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_C1 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_C2 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_C3 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_C4 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_C5 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_C6 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_T1 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_D1 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_D2 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_D3 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_D4 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_D5 = 1'b1;
  assign CLBLL_L_X36Y124_SLICE_X55Y124_D6 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A1 = CLBLM_R_X5Y120_SLICE_X7Y120_A5Q;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A3 = CLBLL_L_X2Y125_SLICE_X1Y125_AQ;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A4 = CLBLL_L_X2Y118_SLICE_X1Y118_AQ;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_A6 = CLBLM_R_X3Y130_SLICE_X2Y130_AO5;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A1 = CLBLM_R_X11Y122_SLICE_X14Y122_DQ;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B1 = CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B2 = CLBLL_L_X2Y125_SLICE_X1Y125_BQ;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B4 = CLBLL_L_X2Y121_SLICE_X1Y121_BQ;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B5 = CLBLM_R_X3Y123_SLICE_X2Y123_CQ;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_B6 = 1'b1;
  assign CLBLM_L_X8Y121_SLICE_X10Y121_A4 = CLBLM_L_X10Y126_SLICE_X12Y126_CQ;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C3 = CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C4 = CLBLL_L_X4Y125_SLICE_X4Y125_CQ;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_C6 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D1 = CLBLL_L_X2Y121_SLICE_X1Y121_BQ;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D2 = CLBLM_R_X3Y126_SLICE_X2Y126_A5Q;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D3 = CLBLM_R_X5Y125_SLICE_X6Y125_A5Q;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D4 = CLBLL_L_X4Y123_SLICE_X5Y123_B5Q;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D5 = 1'b1;
  assign CLBLL_L_X2Y125_SLICE_X1Y125_D6 = CLBLL_L_X2Y122_SLICE_X1Y122_A5Q;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B6 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C4 = CLBLM_R_X7Y126_SLICE_X9Y126_D5Q;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C5 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C6 = CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A2 = CLBLM_R_X7Y120_SLICE_X9Y120_AO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A3 = CLBLM_R_X7Y127_SLICE_X9Y127_AQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A4 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A5 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B4 = CLBLM_L_X10Y129_SLICE_X12Y129_CO6;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_B6 = CLBLM_R_X5Y118_SLICE_X6Y118_B5Q;
  assign LIOB33_X0Y121_IOB_X0Y121_O = CLBLM_R_X5Y128_SLICE_X7Y128_B5Q;
  assign LIOB33_X0Y121_IOB_X0Y122_O = CLBLM_R_X5Y126_SLICE_X7Y126_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A1 = CLBLM_R_X5Y117_SLICE_X6Y117_A5Q;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A2 = CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A3 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A4 = CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A5 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C2 = CLBLM_R_X7Y127_SLICE_X9Y127_CQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_C3 = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B1 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B2 = CLBLM_R_X5Y117_SLICE_X6Y117_DO5;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B3 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B4 = CLBLL_L_X4Y117_SLICE_X5Y117_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B5 = CLBLM_R_X5Y117_SLICE_X6Y117_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_B6 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C1 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C2 = CLBLM_R_X7Y124_SLICE_X8Y124_B5Q;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C3 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C4 = CLBLM_R_X7Y118_SLICE_X8Y118_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C5 = CLBLM_R_X5Y117_SLICE_X7Y117_DO6;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_C6 = CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D3 = CLBLM_R_X7Y126_SLICE_X9Y126_B5Q;
  assign CLBLM_R_X7Y127_SLICE_X9Y127_D4 = CLBLM_R_X7Y127_SLICE_X9Y127_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A1 = CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A2 = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A3 = CLBLM_R_X7Y127_SLICE_X8Y127_AQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A5 = CLBLM_R_X7Y119_SLICE_X9Y119_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D1 = CLBLM_R_X7Y124_SLICE_X8Y124_BQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D2 = CLBLM_R_X5Y117_SLICE_X6Y117_A5Q;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D3 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D4 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D5 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X7Y117_D6 = CLBLM_R_X7Y121_SLICE_X9Y121_BQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_A6 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B1 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B2 = CLBLM_R_X7Y127_SLICE_X8Y127_BQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B3 = CLBLM_R_X7Y125_SLICE_X8Y125_AQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A1 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A2 = CLBLM_R_X5Y117_SLICE_X6Y117_BQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A3 = CLBLM_R_X5Y117_SLICE_X6Y117_AQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A4 = CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_A6 = 1'b1;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C2 = CLBLM_R_X7Y127_SLICE_X8Y127_CQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_AX = CLBLM_R_X5Y117_SLICE_X6Y117_DO6;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_C3 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B1 = CLBLM_R_X3Y124_SLICE_X3Y124_CQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B2 = CLBLM_R_X5Y117_SLICE_X6Y117_BQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B4 = CLBLM_R_X5Y117_SLICE_X6Y117_CQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_B6 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D1 = CLBLM_R_X7Y130_SLICE_X9Y130_AQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D2 = CLBLM_R_X3Y124_SLICE_X2Y124_B5Q;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C1 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C2 = CLBLM_R_X7Y117_SLICE_X9Y117_CO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C4 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C5 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_C6 = CLBLM_R_X5Y126_SLICE_X6Y126_BQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D3 = CLBLM_R_X7Y127_SLICE_X8Y127_DQ;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D5 = 1'b1;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y127_SLICE_X8Y127_D6 = CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D2 = CLBLM_R_X5Y125_SLICE_X6Y125_A5Q;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D3 = CLBLM_L_X10Y119_SLICE_X13Y119_AQ;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D4 = CLBLM_R_X5Y117_SLICE_X6Y117_A5Q;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D5 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X5Y117_SLICE_X6Y117_D6 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1 = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1 = 1'b1;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_A1 = CLBLL_L_X2Y130_SLICE_X0Y130_CO6;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_A2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_A3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_A4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_A5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_A6 = 1'b1;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_B1 = CLBLL_L_X2Y128_SLICE_X0Y128_BO5;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_B2 = CLBLL_L_X2Y125_SLICE_X1Y125_BQ;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_B3 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_B4 = CLBLM_R_X5Y128_SLICE_X6Y128_A5Q;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_B5 = CLBLL_L_X2Y126_SLICE_X0Y126_AO6;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_B6 = CLBLL_L_X2Y126_SLICE_X0Y126_AO5;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_C1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_C2 = CLBLM_R_X3Y124_SLICE_X2Y124_A5Q;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_C3 = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_C4 = CLBLL_L_X2Y130_SLICE_X0Y130_BO6;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_C5 = CLBLL_L_X2Y130_SLICE_X0Y130_CO6;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_C6 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_D1 = 1'b1;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_D2 = 1'b1;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_D3 = 1'b1;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_D4 = 1'b1;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_D5 = 1'b1;
  assign CLBLL_L_X2Y126_SLICE_X0Y126_D6 = 1'b1;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_A1 = CLBLL_L_X2Y126_SLICE_X1Y126_AQ;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_A3 = CLBLL_L_X2Y121_SLICE_X1Y121_BQ;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_A4 = CLBLM_R_X3Y132_SLICE_X2Y132_CO5;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_A5 = CLBLL_L_X2Y125_SLICE_X1Y125_AQ;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_A6 = CLBLM_R_X3Y130_SLICE_X2Y130_AO5;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_B1 = CLBLL_L_X2Y130_SLICE_X0Y130_CO6;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_B2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_B3 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_B4 = CLBLL_L_X2Y130_SLICE_X0Y130_AO6;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_B5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_B6 = CLBLM_R_X3Y124_SLICE_X2Y124_BQ;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_C1 = CLBLM_R_X3Y123_SLICE_X2Y123_BQ;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_C2 = CLBLM_R_X3Y122_SLICE_X2Y122_AQ;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_C3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_C4 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_C5 = CLBLL_L_X2Y128_SLICE_X1Y128_BO5;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_C6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_A1 = CLBLM_L_X12Y121_SLICE_X16Y121_BQ;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_A2 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_A3 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_A4 = CLBLM_R_X11Y131_SLICE_X15Y131_AQ;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_A6 = 1'b1;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_D1 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_D2 = 1'b1;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_D3 = CLBLL_L_X2Y128_SLICE_X0Y128_BO5;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_D4 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_D5 = CLBLM_R_X3Y129_SLICE_X3Y129_AO5;
  assign CLBLL_L_X2Y126_SLICE_X1Y126_D6 = CLBLL_L_X2Y126_SLICE_X1Y126_BO6;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_B1 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_B2 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_B3 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_B4 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_B5 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_B6 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_C1 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_C2 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_C3 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_C4 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_C5 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_C6 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_D1 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_D2 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_D3 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_D4 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_D5 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X163Y173_D6 = 1'b1;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_D = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_A1 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_A2 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_A3 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_A4 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_A5 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_A6 = 1'b1;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_D = RIOB33_X105Y125_IOB_X1Y126_I;
  assign LIOB33_X0Y123_IOB_X0Y124_O = CLBLL_L_X4Y122_SLICE_X5Y122_C5Q;
  assign LIOB33_X0Y123_IOB_X0Y123_O = CLBLL_L_X4Y118_SLICE_X5Y118_C5Q;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_D = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_B1 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_B2 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_B3 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_B4 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_B5 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_B6 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_C1 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_C2 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_C3 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A1 = CLBLM_L_X8Y127_SLICE_X11Y127_AQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A2 = CLBLM_R_X5Y130_SLICE_X7Y130_DO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A3 = CLBLM_R_X7Y128_SLICE_X9Y128_AQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A4 = CLBLM_R_X7Y126_SLICE_X9Y126_D5Q;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_A6 = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_C4 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_C5 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_C6 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B1 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B4 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B5 = CLBLM_L_X10Y129_SLICE_X12Y129_CO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_B6 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_D1 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_D2 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A1 = CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A2 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A3 = CLBLM_R_X5Y118_SLICE_X7Y118_AQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A4 = CLBLL_L_X4Y117_SLICE_X5Y117_AQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A5 = CLBLM_L_X10Y123_SLICE_X12Y123_AQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C1 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C2 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_AX = CLBLM_R_X5Y119_SLICE_X6Y119_BO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C3 = CLBLM_L_X8Y129_SLICE_X11Y129_B5Q;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B1 = CLBLM_R_X3Y128_SLICE_X3Y128_BO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B2 = CLBLM_R_X3Y130_SLICE_X3Y130_BO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B3 = CLBLM_R_X3Y128_SLICE_X2Y128_AO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B5 = CLBLM_R_X3Y126_SLICE_X3Y126_AO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_B6 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D1 = CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C1 = CLBLL_L_X4Y128_SLICE_X4Y128_AO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C2 = CLBLM_R_X3Y127_SLICE_X2Y127_DO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C3 = CLBLL_L_X2Y127_SLICE_X0Y127_CO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C4 = CLBLM_R_X3Y124_SLICE_X3Y124_DO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C5 = CLBLM_R_X5Y118_SLICE_X7Y118_BO5;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_C6 = CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D3 = CLBLM_R_X7Y131_SLICE_X9Y131_DO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D4 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y127_SLICE_X13Y127_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A3 = CLBLM_R_X7Y128_SLICE_X8Y128_AQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A5 = CLBLM_L_X10Y126_SLICE_X13Y126_CQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A6 = CLBLM_L_X8Y127_SLICE_X11Y127_CQ;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D1 = CLBLL_L_X2Y122_SLICE_X1Y122_CO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D2 = CLBLM_R_X3Y127_SLICE_X2Y127_DO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D3 = CLBLL_L_X2Y127_SLICE_X0Y127_CO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D4 = CLBLL_L_X4Y128_SLICE_X4Y128_AO6;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D5 = CLBLM_R_X5Y118_SLICE_X7Y118_BO5;
  assign CLBLM_R_X5Y118_SLICE_X7Y118_D6 = CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B1 = CLBLM_L_X8Y128_SLICE_X11Y128_DQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B2 = CLBLM_R_X7Y128_SLICE_X8Y128_BQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B3 = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B4 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A1 = CLBLM_L_X8Y126_SLICE_X11Y126_B5Q;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A2 = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A4 = CLBLM_L_X8Y119_SLICE_X11Y119_BQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A5 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_A6 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C2 = CLBLM_R_X7Y128_SLICE_X8Y128_CQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C3 = CLBLM_R_X7Y125_SLICE_X8Y125_BQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B1 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B2 = CLBLM_R_X5Y118_SLICE_X6Y118_BQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B3 = CLBLM_R_X5Y117_SLICE_X7Y117_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B4 = CLBLM_R_X5Y118_SLICE_X7Y118_DO6;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B5 = CLBLM_R_X5Y123_SLICE_X7Y123_C5Q;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D1 = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_BX = CLBLM_R_X5Y118_SLICE_X6Y118_CO6;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C3 = CLBLM_R_X5Y119_SLICE_X6Y119_DQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C4 = CLBLM_L_X8Y123_SLICE_X11Y123_CQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C5 = CLBLM_R_X5Y118_SLICE_X6Y118_B5Q;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_C6 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D3 = CLBLM_R_X7Y128_SLICE_X8Y128_DQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D4 = CLBLM_R_X5Y126_SLICE_X7Y126_CO5;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D5 = 1'b1;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_D6 = CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D1 = CLBLM_L_X10Y118_SLICE_X12Y118_AQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D2 = CLBLM_R_X7Y120_SLICE_X8Y120_BQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D3 = CLBLM_R_X5Y118_SLICE_X6Y118_DQ;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y118_SLICE_X6Y118_D6 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_C4 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A1 = CLBLL_L_X2Y127_SLICE_X0Y127_BO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A2 = CLBLL_L_X2Y122_SLICE_X1Y122_BQ;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A3 = CLBLL_L_X2Y128_SLICE_X0Y128_AO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A4 = CLBLL_L_X4Y129_SLICE_X4Y129_BO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A5 = CLBLM_R_X3Y124_SLICE_X2Y124_DQ;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_A6 = CLBLL_L_X2Y126_SLICE_X1Y126_CO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B4 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_B6 = CLBLM_R_X5Y126_SLICE_X6Y126_BQ;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C1 = CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C2 = CLBLL_L_X2Y128_SLICE_X0Y128_AO5;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C3 = CLBLL_L_X2Y129_SLICE_X1Y129_DO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C4 = CLBLL_L_X2Y129_SLICE_X0Y129_CO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C5 = CLBLL_L_X2Y127_SLICE_X0Y127_DO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_C6 = CLBLM_R_X5Y126_SLICE_X6Y126_BQ;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D1 = CLBLL_L_X2Y128_SLICE_X0Y128_AO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D2 = CLBLL_L_X2Y126_SLICE_X1Y126_CO6;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D3 = CLBLM_R_X3Y124_SLICE_X2Y124_DQ;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D4 = CLBLL_L_X2Y122_SLICE_X1Y122_BQ;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D5 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X0Y127_D6 = CLBLL_L_X4Y129_SLICE_X4Y129_BO6;
  assign CLBLL_L_X4Y127_SLICE_X5Y127_D1 = CLBLL_L_X4Y122_SLICE_X5Y122_AQ;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A1 = CLBLL_L_X2Y127_SLICE_X1Y127_DO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A2 = CLBLM_R_X3Y127_SLICE_X2Y127_AO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A3 = CLBLM_R_X3Y129_SLICE_X3Y129_AO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A4 = CLBLL_L_X2Y127_SLICE_X1Y127_BO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A5 = CLBLM_R_X3Y126_SLICE_X2Y126_CO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_A6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B1 = CLBLL_L_X2Y128_SLICE_X1Y128_AO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B2 = CLBLL_L_X2Y130_SLICE_X0Y130_BO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B3 = CLBLM_R_X3Y125_SLICE_X3Y125_BQ;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B4 = CLBLM_R_X3Y122_SLICE_X3Y122_BQ;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B5 = CLBLL_L_X2Y130_SLICE_X0Y130_CO5;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_B6 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C1 = CLBLL_L_X2Y127_SLICE_X1Y127_AO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C2 = CLBLL_L_X2Y129_SLICE_X1Y129_BO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C3 = CLBLL_L_X4Y125_SLICE_X5Y125_CO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C4 = CLBLL_L_X2Y129_SLICE_X1Y129_AO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C5 = CLBLL_L_X2Y127_SLICE_X0Y127_AO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_C6 = CLBLM_R_X3Y126_SLICE_X3Y126_BO6;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_D = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D1 = 1'b1;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D2 = CLBLL_L_X2Y130_SLICE_X0Y130_BO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D3 = CLBLL_L_X2Y130_SLICE_X0Y130_CO6;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D4 = CLBLM_R_X7Y127_SLICE_X8Y127_DQ;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D5 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLL_L_X2Y127_SLICE_X1Y127_D6 = CLBLL_L_X2Y130_SLICE_X0Y130_AO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A6 = 1'b1;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_D = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOB33_X0Y125_IOB_X0Y126_O = CLBLM_R_X3Y125_SLICE_X2Y125_AQ;
  assign LIOB33_X0Y125_IOB_X0Y125_O = CLBLM_L_X8Y123_SLICE_X10Y123_C5Q;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B3 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B4 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B5 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A2 = CLBLM_R_X7Y131_SLICE_X9Y131_BO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A3 = CLBLM_R_X7Y129_SLICE_X9Y129_AQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A4 = CLBLM_R_X7Y131_SLICE_X8Y131_CO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A5 = CLBLM_R_X7Y129_SLICE_X9Y129_DQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A6 = CLBLM_L_X8Y129_SLICE_X10Y129_BO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B2 = CLBLM_R_X5Y129_SLICE_X6Y129_BQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B4 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C2 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B5 = CLBLM_R_X7Y131_SLICE_X9Y131_BO5;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B6 = CLBLM_R_X11Y126_SLICE_X14Y126_DQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C3 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A1 = CLBLM_R_X5Y116_SLICE_X7Y116_AQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A2 = CLBLM_R_X5Y126_SLICE_X7Y126_CO5;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A3 = CLBLM_R_X5Y119_SLICE_X7Y119_AQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A4 = CLBLL_L_X4Y122_SLICE_X4Y122_BQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C4 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_A6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C1 = CLBLM_R_X7Y131_SLICE_X9Y131_BO5;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C5 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B1 = CLBLM_R_X5Y118_SLICE_X6Y118_DQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B2 = CLBLM_R_X5Y119_SLICE_X7Y119_BQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B4 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_B6 = CLBLL_L_X2Y122_SLICE_X1Y122_A5Q;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C1 = CLBLL_L_X4Y126_SLICE_X4Y126_AQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C2 = CLBLM_R_X5Y119_SLICE_X7Y119_CQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C5 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_C6 = CLBLM_L_X8Y119_SLICE_X11Y119_AQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D3 = CLBLM_R_X7Y129_SLICE_X9Y129_DQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D4 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A1 = CLBLM_R_X7Y130_SLICE_X8Y130_DO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A2 = CLBLM_L_X8Y122_SLICE_X10Y122_BQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A4 = CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A5 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D1 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D2 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D3 = CLBLM_R_X3Y123_SLICE_X2Y123_DQ;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D5 = CLBLM_R_X3Y127_SLICE_X2Y127_DO6;
  assign CLBLM_R_X5Y119_SLICE_X7Y119_D6 = CLBLM_L_X8Y123_SLICE_X11Y123_DO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B2 = CLBLM_R_X7Y126_SLICE_X9Y126_C5Q;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B4 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A1 = CLBLM_R_X5Y120_SLICE_X6Y120_CQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A3 = CLBLM_R_X5Y117_SLICE_X6Y117_AQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A4 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_A6 = CLBLM_L_X8Y123_SLICE_X11Y123_DO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C1 = CLBLM_R_X7Y129_SLICE_X8Y129_BQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C2 = CLBLM_R_X7Y129_SLICE_X8Y129_CQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B2 = CLBLM_R_X5Y119_SLICE_X6Y119_DQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B4 = CLBLM_L_X8Y124_SLICE_X10Y124_BQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B5 = CLBLL_L_X4Y129_SLICE_X5Y129_AQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_B6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D2 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C1 = CLBLM_R_X5Y116_SLICE_X6Y116_AQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C2 = CLBLM_R_X5Y119_SLICE_X6Y119_CQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C4 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C5 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_C6 = CLBLM_R_X3Y123_SLICE_X3Y123_CQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D3 = CLBLM_R_X7Y129_SLICE_X8Y129_DQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D4 = CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D6 = CLBLM_L_X8Y127_SLICE_X11Y127_DQ;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D5 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D2 = CLBLL_L_X4Y120_SLICE_X5Y120_AQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D3 = CLBLM_R_X5Y119_SLICE_X7Y119_DO6;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D6 = 1'b1;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D5 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X5Y119_SLICE_X6Y119_D6 = CLBLM_R_X5Y119_SLICE_X6Y119_DQ;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_A1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_A2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_A3 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_A4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_A6 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_B1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_B2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_B4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_B5 = CLBLL_L_X2Y130_SLICE_X0Y130_CO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_B6 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_C1 = CLBLL_L_X2Y130_SLICE_X1Y130_AO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_C2 = CLBLL_L_X2Y128_SLICE_X1Y128_AO5;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_C3 = CLBLL_L_X2Y130_SLICE_X0Y130_CO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_C4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_C5 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_C6 = CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_D1 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_D1 = CLBLL_L_X2Y119_SLICE_X1Y119_AQ;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_D2 = CLBLL_L_X2Y130_SLICE_X0Y130_BO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_D3 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_D4 = CLBLL_L_X2Y130_SLICE_X0Y130_CO6;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_D5 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X0Y128_D6 = CLBLL_L_X2Y130_SLICE_X0Y130_AO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_T1 = 1'b1;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_D = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_D1 = CLBLM_L_X12Y126_SLICE_X16Y126_AQ;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_D1 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_AX = CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_T1 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_A1 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B1 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_A2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_A3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_A5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B2 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_A6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_T1 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_B1 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B3 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_B2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_B3 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_B4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_B5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B4 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_B6 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_T1 = 1'b1;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_C1 = CLBLL_L_X2Y128_SLICE_X1Y128_AO6;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_C2 = CLBLL_L_X2Y130_SLICE_X0Y130_CO6;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_C3 = CLBLL_L_X2Y130_SLICE_X0Y130_CO5;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_C4 = CLBLL_L_X2Y128_SLICE_X1Y128_AO5;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_C5 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_C6 = CLBLM_R_X5Y127_SLICE_X7Y127_CQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B5 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B6 = 1'b1;
  assign LIOB33_X0Y127_IOB_X0Y128_O = CLBLL_L_X2Y118_SLICE_X1Y118_B5Q;
  assign LIOB33_X0Y127_IOB_X0Y127_O = CLBLL_L_X4Y126_SLICE_X4Y126_AQ;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_D1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_D2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_D3 = CLBLL_L_X4Y130_SLICE_X4Y130_AO5;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_D4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_D5 = CLBLL_L_X2Y130_SLICE_X1Y130_AO5;
  assign CLBLL_L_X2Y128_SLICE_X1Y128_D6 = CLBLL_L_X2Y128_SLICE_X1Y128_BO6;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_A1 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_A6 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_A2 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_B1 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_B2 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_B3 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_B4 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_B5 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_B6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C1 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_C1 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_C2 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_C3 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_C4 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C2 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_C5 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_C6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C3 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C4 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_D1 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_D2 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_D3 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_D4 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C5 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_D5 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X163Y175_D6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C6 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_A1 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_A2 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_A3 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_A4 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_A5 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_A6 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_B1 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_B2 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_B3 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_B4 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_B5 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_B6 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_C1 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_C2 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_C3 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A1 = CLBLM_R_X7Y130_SLICE_X9Y130_BO5;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A2 = CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A3 = CLBLM_R_X7Y124_SLICE_X9Y124_BO5;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A4 = CLBLM_R_X7Y130_SLICE_X9Y130_DO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A5 = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_C4 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_C5 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_C6 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B1 = CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B2 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B3 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B4 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B5 = CLBLM_L_X8Y131_SLICE_X10Y131_DO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B6 = 1'b1;
  assign CLBLM_R_X103Y175_SLICE_X162Y175_D1 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A1 = CLBLM_R_X5Y122_SLICE_X7Y122_BQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A2 = CLBLM_R_X3Y119_SLICE_X3Y119_CO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A3 = CLBLM_R_X7Y118_SLICE_X9Y118_AQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A4 = CLBLM_R_X5Y126_SLICE_X7Y126_DO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_A6 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C1 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D1 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C2 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B2 = CLBLM_R_X5Y120_SLICE_X7Y120_BQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D2 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B4 = CLBLL_L_X4Y125_SLICE_X4Y125_BQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B5 = CLBLM_R_X5Y118_SLICE_X7Y118_BO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_B6 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D3 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C1 = CLBLM_R_X5Y121_SLICE_X7Y121_AQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C2 = CLBLM_L_X8Y123_SLICE_X11Y123_AQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D4 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C3 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C5 = CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_C6 = CLBLL_L_X4Y121_SLICE_X4Y121_DQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D5 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A1 = CLBLM_R_X5Y130_SLICE_X7Y130_DO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A2 = CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A3 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D6 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A4 = CLBLL_L_X4Y124_SLICE_X4Y124_CQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D1 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D3 = CLBLM_R_X5Y121_SLICE_X6Y121_CO6;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D4 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D5 = CLBLM_R_X3Y123_SLICE_X2Y123_DQ;
  assign CLBLM_R_X5Y120_SLICE_X7Y120_D6 = CLBLM_R_X3Y130_SLICE_X3Y130_BO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B2 = CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B4 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B5 = CLBLM_L_X8Y127_SLICE_X10Y127_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B6 = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B1 = CLBLM_R_X5Y130_SLICE_X7Y130_DO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A1 = CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A2 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A3 = CLBLM_R_X5Y120_SLICE_X6Y120_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A4 = CLBLM_L_X10Y120_SLICE_X13Y120_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_A6 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C1 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C2 = CLBLM_L_X8Y129_SLICE_X11Y129_B5Q;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B2 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B4 = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B5 = CLBLM_R_X7Y121_SLICE_X8Y121_DO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_B6 = CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D1 = CLBLM_L_X8Y127_SLICE_X10Y127_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C2 = CLBLM_R_X5Y125_SLICE_X6Y125_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C3 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C5 = CLBLM_R_X5Y121_SLICE_X6Y121_CO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_C6 = CLBLM_R_X3Y120_SLICE_X3Y120_BQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D3 = CLBLM_R_X5Y130_SLICE_X7Y130_DO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D4 = CLBLM_R_X7Y130_SLICE_X8Y130_CO5;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D5 = CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D2 = CLBLM_L_X8Y129_SLICE_X11Y129_BQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D3 = CLBLM_R_X11Y127_SLICE_X15Y127_CO6;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D2 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D3 = CLBLM_R_X5Y120_SLICE_X6Y120_DQ;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D5 = 1'b1;
  assign CLBLM_R_X5Y120_SLICE_X6Y120_D6 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D5 = CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  assign CLBLM_R_X11Y126_SLICE_X15Y126_D6 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A3 = CLBLL_L_X2Y130_SLICE_X0Y130_CO5;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_A6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B1 = CLBLL_L_X2Y130_SLICE_X0Y130_BO5;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B2 = CLBLL_L_X2Y130_SLICE_X0Y130_AO6;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B3 = CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B4 = CLBLL_L_X2Y130_SLICE_X0Y130_BO6;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B5 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_B6 = CLBLL_L_X2Y130_SLICE_X0Y130_CO6;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C3 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C5 = CLBLL_L_X2Y130_SLICE_X1Y130_AO5;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_C6 = CLBLL_L_X2Y118_SLICE_X1Y118_CO6;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D1 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D2 = CLBLL_L_X2Y128_SLICE_X1Y128_AO5;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D3 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D4 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D5 = CLBLL_L_X2Y130_SLICE_X1Y130_BO5;
  assign CLBLL_L_X2Y129_SLICE_X0Y129_D6 = CLBLL_L_X2Y130_SLICE_X0Y130_CO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A4 = CLBLM_R_X5Y127_SLICE_X7Y127_BQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_A6 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A1 = CLBLL_L_X2Y129_SLICE_X0Y129_AO5;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A2 = CLBLM_R_X3Y130_SLICE_X2Y130_BO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A3 = CLBLL_L_X2Y129_SLICE_X0Y129_CO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A4 = CLBLL_L_X2Y130_SLICE_X1Y130_CO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A5 = CLBLL_L_X2Y128_SLICE_X0Y128_CO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_A6 = CLBLL_L_X2Y130_SLICE_X0Y130_AO5;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C4 = CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  assign LIOB33_X0Y129_IOB_X0Y129_O = CLBLM_R_X3Y123_SLICE_X3Y123_CQ;
  assign LIOB33_X0Y129_IOB_X0Y130_O = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B1 = CLBLM_R_X3Y130_SLICE_X3Y130_AO5;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B2 = CLBLL_L_X4Y129_SLICE_X4Y129_BO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B3 = CLBLL_L_X2Y128_SLICE_X0Y128_CO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B4 = CLBLM_R_X3Y130_SLICE_X2Y130_BO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B5 = CLBLL_L_X2Y130_SLICE_X1Y130_CO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_B6 = CLBLL_L_X2Y129_SLICE_X0Y129_AO6;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C5 = CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_C6 = CLBLM_R_X5Y118_SLICE_X7Y118_BO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D6 = 1'b1;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C1 = CLBLL_L_X2Y129_SLICE_X0Y129_BO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C2 = CLBLL_L_X2Y129_SLICE_X0Y129_AO5;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C3 = CLBLM_R_X3Y129_SLICE_X3Y129_AO5;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C4 = CLBLM_R_X3Y130_SLICE_X3Y130_AO5;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C5 = CLBLL_L_X2Y128_SLICE_X1Y128_DO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_C6 = CLBLL_L_X2Y130_SLICE_X1Y130_CO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B3 = CLBLM_R_X11Y128_SLICE_X14Y128_AO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B4 = CLBLM_L_X10Y125_SLICE_X13Y125_DO5;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B5 = CLBLL_L_X2Y120_SLICE_X1Y120_AQ;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D1 = CLBLL_L_X2Y128_SLICE_X0Y128_CO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D2 = CLBLL_L_X4Y129_SLICE_X4Y129_BO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D3 = CLBLL_L_X2Y130_SLICE_X1Y130_CO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D4 = CLBLL_L_X2Y130_SLICE_X0Y130_AO5;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D5 = CLBLL_L_X2Y129_SLICE_X0Y129_AO6;
  assign CLBLL_L_X2Y129_SLICE_X1Y129_D6 = CLBLM_R_X3Y130_SLICE_X2Y130_BO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D2 = CLBLM_R_X5Y130_SLICE_X7Y130_CO5;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C3 = CLBLM_R_X11Y128_SLICE_X15Y128_CO6;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D5 = CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C5 = CLBLM_L_X10Y126_SLICE_X12Y126_CQ;
  assign CLBLM_R_X7Y128_SLICE_X9Y128_D6 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLM_R_X11Y126_SLICE_X14Y126_C6 = CLBLM_R_X11Y127_SLICE_X15Y127_BO5;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A1 = CLBLM_R_X7Y131_SLICE_X8Y131_CO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A2 = CLBLM_R_X5Y127_SLICE_X7Y127_BQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A3 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A4 = CLBLM_R_X7Y131_SLICE_X9Y131_BO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A6 = CLBLM_L_X8Y131_SLICE_X11Y131_BO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B1 = CLBLM_L_X8Y131_SLICE_X10Y131_DO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B2 = CLBLM_L_X8Y129_SLICE_X11Y129_B5Q;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B3 = CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B4 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B5 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A1 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B6 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A1 = CLBLM_L_X8Y121_SLICE_X10Y121_DO5;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A2 = CLBLM_R_X7Y121_SLICE_X9Y121_B5Q;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A4 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A5 = CLBLM_L_X8Y123_SLICE_X11Y123_AQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_A2 = CLBLM_R_X5Y126_SLICE_X7Y126_CO5;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C1 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C2 = CLBLM_L_X8Y129_SLICE_X11Y129_B5Q;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B1 = CLBLM_R_X7Y120_SLICE_X8Y120_AQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B2 = CLBLM_L_X8Y122_SLICE_X11Y122_AQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B4 = CLBLL_L_X4Y123_SLICE_X5Y123_BQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B5 = CLBLM_R_X7Y121_SLICE_X8Y121_AQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_B6 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D1 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C1 = CLBLM_R_X3Y120_SLICE_X2Y120_CQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C2 = CLBLL_L_X4Y121_SLICE_X4Y121_DQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C3 = CLBLM_L_X8Y123_SLICE_X11Y123_AQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C4 = CLBLL_L_X4Y121_SLICE_X5Y121_DO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C5 = CLBLM_R_X5Y122_SLICE_X7Y122_DO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_C6 = CLBLM_R_X7Y118_SLICE_X8Y118_CQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D3 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D4 = CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A3 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A4 = CLBLM_R_X7Y131_SLICE_X8Y131_BO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A5 = CLBLM_L_X8Y127_SLICE_X10Y127_BQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D1 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D3 = CLBLL_L_X2Y127_SLICE_X0Y127_CO6;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D4 = CLBLM_R_X7Y117_SLICE_X8Y117_AQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D5 = CLBLM_R_X3Y123_SLICE_X2Y123_DQ;
  assign CLBLM_R_X5Y121_SLICE_X7Y121_D6 = CLBLM_R_X5Y121_SLICE_X7Y121_BO5;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A6 = CLBLM_L_X8Y131_SLICE_X10Y131_DO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C4 = CLBLM_R_X5Y130_SLICE_X7Y130_BQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B1 = CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B2 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B3 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A1 = CLBLM_R_X5Y121_SLICE_X6Y121_DO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A2 = CLBLM_R_X11Y120_SLICE_X15Y120_AQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A3 = CLBLM_R_X5Y121_SLICE_X6Y121_AQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A4 = CLBLM_R_X5Y121_SLICE_X7Y121_CO6;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C5 = CLBLM_R_X7Y129_SLICE_X9Y129_CQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C6 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B2 = CLBLM_R_X5Y125_SLICE_X7Y125_AQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B4 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B5 = CLBLM_R_X5Y119_SLICE_X6Y119_AQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_B6 = CLBLM_R_X5Y121_SLICE_X7Y121_BO5;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D1 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D2 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C2 = CLBLM_R_X7Y121_SLICE_X9Y121_B5Q;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C3 = CLBLL_L_X4Y122_SLICE_X4Y122_DQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C4 = CLBLM_R_X7Y120_SLICE_X8Y120_BQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C5 = CLBLL_L_X4Y121_SLICE_X4Y121_CQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_C6 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_B6 = CLBLM_R_X5Y126_SLICE_X7Y126_CO5;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D3 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D4 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D6 = 1'b1;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D1 = CLBLM_R_X5Y119_SLICE_X6Y119_AQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D2 = CLBLM_R_X5Y120_SLICE_X6Y120_CQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D3 = CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D4 = CLBLM_L_X8Y121_SLICE_X10Y121_BQ;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y121_SLICE_X6Y121_D6 = CLBLM_R_X3Y120_SLICE_X3Y120_BQ;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_A1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_A2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_A3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_A4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_A5 = CLBLL_L_X2Y130_SLICE_X0Y130_CO5;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_A6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D2 = CLBLM_R_X7Y129_SLICE_X9Y129_CQ;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_B1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_B2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_B3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_B4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_B5 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_B6 = 1'b1;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C4 = CLBLM_R_X5Y126_SLICE_X7Y126_CO5;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_C1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_C2 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_C3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_C4 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_C5 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_C6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D5 = CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D6 = CLBLM_R_X5Y130_SLICE_X7Y130_AQ;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C5 = CLBLM_L_X8Y129_SLICE_X11Y129_B5Q;
  assign CLBLM_R_X7Y128_SLICE_X8Y128_C6 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_D1 = CLBLL_L_X2Y131_SLICE_X1Y131_AO6;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_D2 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_D3 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_D4 = CLBLL_L_X2Y130_SLICE_X0Y130_CO6;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_D5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y130_SLICE_X0Y130_D6 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D2 = CLBLM_L_X10Y119_SLICE_X12Y119_BQ;
  assign LIOB33_X0Y131_IOB_X0Y132_O = CLBLM_R_X5Y118_SLICE_X6Y118_AQ;
  assign LIOB33_X0Y131_IOB_X0Y131_O = CLBLM_R_X5Y118_SLICE_X6Y118_AO5;
  assign CLBLM_L_X8Y122_SLICE_X11Y122_D3 = CLBLM_L_X10Y126_SLICE_X13Y126_DQ;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_A1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_A2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_A3 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_A5 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_A6 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_B1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_B2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_B3 = CLBLL_L_X2Y130_SLICE_X0Y130_CO6;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_B4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_B6 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_C1 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_C2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_C3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_C4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_C5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_C6 = CLBLL_L_X2Y130_SLICE_X0Y130_CO6;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_D1 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_D2 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_D3 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_D4 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_D5 = 1'b1;
  assign CLBLL_L_X2Y130_SLICE_X1Y130_D6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A3 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A4 = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A5 = CLBLM_R_X11Y125_SLICE_X14Y125_AQ;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C4 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B5 = CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C6 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B6 = CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_D1 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A1 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B2 = CLBLM_L_X10Y126_SLICE_X12Y126_CQ;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A5 = 1'b1;
  assign CLBLM_L_X8Y122_SLICE_X10Y122_B3 = CLBLM_R_X5Y124_SLICE_X7Y124_C5Q;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_T1 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_D1 = CLBLM_L_X12Y121_SLICE_X16Y121_BQ;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_D1 = LIOB33_X0Y71_IOB_X0Y71_I;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_T1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C4 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C4 = CLBLM_R_X7Y129_SLICE_X9Y129_CQ;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_T1 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C5 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_D1 = CLBLM_L_X8Y126_SLICE_X10Y126_AQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C6 = CLBLM_R_X5Y130_SLICE_X7Y130_BQ;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D6 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_T1 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A2 = CLBLM_R_X5Y122_SLICE_X6Y122_DO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A3 = CLBLM_R_X5Y122_SLICE_X7Y122_AQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A4 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A5 = CLBLM_L_X10Y123_SLICE_X12Y123_BQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_A6 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B1 = CLBLM_L_X8Y124_SLICE_X10Y124_DO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B2 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B4 = CLBLM_R_X5Y121_SLICE_X7Y121_AQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B5 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOB33_X0Y101_IOB_X0Y102_O = CLBLL_L_X2Y117_SLICE_X0Y117_BO6;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C1 = CLBLM_R_X7Y123_SLICE_X9Y123_DO5;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C2 = CLBLM_R_X3Y120_SLICE_X2Y120_BQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C4 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C5 = CLBLL_L_X4Y124_SLICE_X4Y124_DQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_C6 = CLBLL_L_X4Y123_SLICE_X5Y123_BQ;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_D3 = 1'b1;
  assign LIOB33_X0Y101_IOB_X0Y101_O = CLBLL_L_X2Y118_SLICE_X0Y118_AO5;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_D4 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D1 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D2 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D4 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D5 = CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  assign CLBLM_R_X5Y122_SLICE_X7Y122_D6 = CLBLM_R_X5Y121_SLICE_X7Y121_AQ;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_D5 = 1'b1;
  assign CLBLM_R_X103Y173_SLICE_X162Y173_D6 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A1 = CLBLL_L_X4Y125_SLICE_X4Y125_BQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A2 = CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A3 = CLBLM_R_X5Y122_SLICE_X6Y122_AQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A4 = CLBLM_R_X7Y122_SLICE_X8Y122_AQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_A6 = CLBLM_R_X7Y121_SLICE_X8Y121_A5Q;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D3 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B1 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B2 = CLBLM_R_X7Y122_SLICE_X9Y122_DO6;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B4 = CLBLL_L_X4Y123_SLICE_X4Y123_BQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B5 = CLBLM_R_X7Y120_SLICE_X8Y120_DQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D4 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C1 = CLBLM_R_X5Y121_SLICE_X6Y121_CO5;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C3 = 1'b1;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C5 = CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_C6 = CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D1 = CLBLL_L_X4Y120_SLICE_X5Y120_BQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D2 = CLBLL_L_X4Y120_SLICE_X5Y120_AQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D3 = CLBLM_R_X5Y123_SLICE_X7Y123_BQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D4 = CLBLM_R_X3Y122_SLICE_X2Y122_CQ;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y122_SLICE_X6Y122_D6 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_A6 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_B6 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_C6 = 1'b1;
  assign LIOB33_X0Y133_IOB_X0Y133_O = CLBLM_R_X3Y132_SLICE_X2Y132_A5Q;
  assign LIOB33_X0Y133_IOB_X0Y134_O = CLBLM_R_X3Y123_SLICE_X2Y123_CQ;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X0Y131_D6 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_A6 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_B6 = 1'b1;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_D = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_D = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_C6 = 1'b1;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D1 = CLBLM_R_X7Y128_SLICE_X9Y128_DO6;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D1 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D2 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D3 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D4 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D5 = 1'b1;
  assign CLBLL_L_X2Y131_SLICE_X1Y131_D6 = 1'b1;
  assign LIOB33_X0Y195_IOB_X0Y196_O = LIOB33_X0Y69_IOB_X0Y69_I;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D2 = CLBLM_L_X8Y129_SLICE_X11Y129_AQ;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D = RIOB33_X105Y143_IOB_X1Y144_I;
  assign RIOB33_X105Y177_IOB_X1Y178_O = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D = RIOB33_X105Y143_IOB_X1Y143_I;
  assign RIOB33_X105Y177_IOB_X1Y177_O = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign CLBLM_L_X8Y129_SLICE_X11Y129_D3 = 1'b1;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_D1 = CLBLL_L_X2Y117_SLICE_X0Y117_AO6;
  assign LIOB33_X0Y191_IOB_X0Y192_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A2 = CLBLM_R_X7Y122_SLICE_X9Y122_CQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A3 = CLBLM_R_X5Y123_SLICE_X7Y123_AQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A4 = CLBLM_R_X5Y126_SLICE_X7Y126_CO5;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A5 = CLBLM_R_X5Y119_SLICE_X6Y119_AQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_A6 = 1'b1;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_T1 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B2 = CLBLM_R_X5Y123_SLICE_X7Y123_BQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B4 = CLBLM_R_X7Y119_SLICE_X8Y119_AQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B5 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_B6 = CLBLM_R_X7Y125_SLICE_X8Y125_CQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C2 = CLBLM_R_X5Y123_SLICE_X7Y123_CQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C4 = CLBLM_R_X5Y127_SLICE_X7Y127_CQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C5 = CLBLL_L_X4Y124_SLICE_X4Y124_BQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_C6 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D1 = CLBLL_L_X4Y122_SLICE_X4Y122_BQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D2 = CLBLM_R_X5Y122_SLICE_X7Y122_BQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D3 = CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D4 = CLBLM_R_X7Y125_SLICE_X8Y125_BQ;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D5 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X7Y123_D6 = CLBLM_R_X5Y120_SLICE_X6Y120_BQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A1 = CLBLM_L_X8Y126_SLICE_X11Y126_B5Q;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A3 = CLBLM_R_X5Y123_SLICE_X6Y123_AQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A4 = CLBLM_L_X8Y124_SLICE_X10Y124_B5Q;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A5 = CLBLL_L_X4Y121_SLICE_X5Y121_AQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_D = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B1 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B3 = CLBLM_R_X5Y123_SLICE_X6Y123_B5Q;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B4 = CLBLM_L_X8Y122_SLICE_X10Y122_A5Q;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B5 = CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_B6 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C2 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C3 = CLBLM_R_X5Y126_SLICE_X6Y126_DQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C4 = CLBLM_L_X8Y122_SLICE_X10Y122_A5Q;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_C6 = 1'b1;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_D = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y128_SLICE_X5Y128_C1 = CLBLL_L_X4Y128_SLICE_X5Y128_AO6;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D1 = CLBLM_R_X7Y122_SLICE_X8Y122_BQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D2 = CLBLM_R_X5Y124_SLICE_X6Y124_A5Q;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D3 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D4 = CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D5 = 1'b1;
  assign CLBLM_R_X5Y123_SLICE_X6Y123_D6 = CLBLL_L_X4Y120_SLICE_X5Y120_A5Q;
  assign LIOB33_X0Y135_IOB_X0Y135_O = CLBLM_R_X3Y129_SLICE_X2Y129_AQ;
  assign LIOB33_X0Y135_IOB_X0Y136_O = CLBLM_R_X3Y132_SLICE_X2Y132_BQ;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_A1 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_A2 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_A3 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_A4 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_A5 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_A6 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_B1 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_B2 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_B3 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_B4 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_B5 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_B6 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_C1 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_C2 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_C3 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_C4 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_C5 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_C6 = 1'b1;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_D = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_D1 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_D2 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_D3 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_D4 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_D5 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X0Y132_D6 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_A1 = CLBLM_R_X3Y132_SLICE_X2Y132_A5Q;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_A2 = CLBLM_R_X3Y123_SLICE_X2Y123_CQ;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_A3 = CLBLM_R_X3Y129_SLICE_X2Y129_AQ;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_A4 = CLBLM_R_X3Y132_SLICE_X2Y132_BQ;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_A5 = CLBLM_R_X3Y131_SLICE_X2Y131_BQ;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_A6 = CLBLM_R_X3Y131_SLICE_X2Y131_AQ;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_B1 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_B2 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_B3 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_B4 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_B5 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_B6 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_C1 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_C2 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_C3 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_C4 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_C5 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_C6 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_T1 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_D1 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_D2 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_D3 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_D4 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_D5 = 1'b1;
  assign CLBLL_L_X2Y132_SLICE_X1Y132_D6 = 1'b1;
  assign CLBLM_R_X5Y116_SLICE_X6Y116_D1 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_D1 = CLBLM_L_X10Y136_SLICE_X12Y136_AO5;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_T1 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A1 = CLBLM_R_X5Y124_SLICE_X7Y124_DO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A2 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A3 = CLBLM_R_X5Y124_SLICE_X7Y124_AQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A4 = CLBLM_R_X7Y127_SLICE_X9Y127_BQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B1 = CLBLM_L_X10Y123_SLICE_X12Y123_CQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B2 = CLBLM_R_X5Y124_SLICE_X7Y124_BQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B3 = CLBLM_R_X7Y121_SLICE_X8Y121_BQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B4 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_B6 = CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C1 = CLBLM_R_X7Y127_SLICE_X9Y127_BQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C3 = CLBLM_L_X8Y122_SLICE_X11Y122_AQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C5 = CLBLM_R_X3Y123_SLICE_X2Y123_BQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_C6 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D1 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D2 = CLBLM_R_X5Y123_SLICE_X7Y123_DO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D3 = CLBLM_R_X7Y126_SLICE_X8Y126_DO6;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D4 = CLBLM_R_X3Y124_SLICE_X3Y124_CQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D5 = CLBLM_R_X11Y126_SLICE_X14Y126_AQ;
  assign CLBLM_R_X5Y124_SLICE_X7Y124_D6 = CLBLM_R_X5Y123_SLICE_X6Y123_DO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A1 = CLBLM_R_X5Y126_SLICE_X6Y126_CQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A3 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A4 = CLBLM_R_X5Y123_SLICE_X6Y123_BQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A5 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_D = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_AX = CLBLM_R_X5Y124_SLICE_X6Y124_DO6;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B1 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B2 = CLBLM_R_X5Y124_SLICE_X6Y124_BQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B3 = CLBLM_R_X7Y124_SLICE_X8Y124_AQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B4 = CLBLL_L_X4Y124_SLICE_X5Y124_DQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_B6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign LIOB33_X0Y137_IOB_X0Y137_O = CLBLM_R_X3Y131_SLICE_X2Y131_AQ;
  assign LIOB33_X0Y137_IOB_X0Y138_O = CLBLM_R_X3Y131_SLICE_X2Y131_BQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_D1 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_D1 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C2 = CLBLM_R_X5Y124_SLICE_X7Y124_C5Q;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C3 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C4 = CLBLM_R_X5Y129_SLICE_X6Y129_AQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C5 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_T1 = 1'b1;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_D1 = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D2 = CLBLM_L_X8Y124_SLICE_X10Y124_B5Q;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D3 = CLBLM_L_X8Y126_SLICE_X11Y126_B5Q;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D4 = CLBLM_R_X3Y124_SLICE_X3Y124_CQ;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y124_SLICE_X6Y124_D6 = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_D1 = LIOB33_X0Y65_IOB_X0Y65_I;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_T1 = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_T1 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_D1 = CLBLM_R_X11Y128_SLICE_X14Y128_AQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_T1 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1 = CLBLL_L_X36Y124_SLICE_X54Y124_AO6;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_D1 = CLBLL_L_X2Y126_SLICE_X1Y126_AQ;
  assign LIOB33_X0Y105_IOB_X0Y106_O = CLBLL_L_X2Y117_SLICE_X0Y117_CO5;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C5 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_C6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_T1 = 1'b1;
  assign CLBLL_L_X4Y118_SLICE_X4Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B4 = CLBLM_R_X11Y126_SLICE_X15Y126_BQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B5 = CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_B6 = 1'b1;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_D = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_D = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A1 = CLBLL_L_X4Y125_SLICE_X4Y125_BQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A2 = CLBLM_L_X8Y130_SLICE_X10Y130_BQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A3 = CLBLM_R_X5Y125_SLICE_X7Y125_AQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A4 = CLBLM_R_X5Y123_SLICE_X7Y123_BQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_A6 = CLBLM_L_X8Y121_SLICE_X11Y121_BQ;
  assign LIOB33_X0Y105_IOB_X0Y105_O = CLBLL_L_X2Y117_SLICE_X0Y117_CO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B1 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B2 = CLBLM_R_X5Y125_SLICE_X7Y125_BQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B3 = CLBLM_R_X5Y124_SLICE_X7Y124_BQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B4 = CLBLM_R_X3Y120_SLICE_X2Y120_CQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_B6 = CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C2 = CLBLM_R_X11Y127_SLICE_X15Y127_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C3 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C1 = CLBLM_R_X3Y128_SLICE_X2Y128_AO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C2 = CLBLM_R_X3Y126_SLICE_X3Y126_AO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C3 = CLBLM_R_X5Y125_SLICE_X6Y125_DO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C4 = CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C5 = CLBLM_R_X5Y125_SLICE_X7Y125_DO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_C6 = CLBLL_L_X4Y128_SLICE_X4Y128_AO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C4 = CLBLM_R_X11Y128_SLICE_X14Y128_AO5;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C5 = CLBLM_L_X12Y127_SLICE_X16Y127_CO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y139_IOB_X0Y140_O = CLBLL_L_X2Y125_SLICE_X1Y125_AQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_C6 = 1'b1;
  assign LIOB33_X0Y139_IOB_X0Y139_O = CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D1 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D2 = CLBLM_R_X3Y128_SLICE_X3Y128_BO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D3 = CLBLM_R_X3Y130_SLICE_X3Y130_BO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D4 = CLBLM_R_X7Y123_SLICE_X8Y123_BQ;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D5 = CLBLL_L_X2Y127_SLICE_X0Y127_CO6;
  assign CLBLM_R_X5Y125_SLICE_X7Y125_D6 = CLBLM_R_X3Y127_SLICE_X2Y127_DO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A1 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A2 = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A4 = CLBLM_L_X8Y121_SLICE_X10Y121_BQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_A6 = CLBLM_R_X5Y125_SLICE_X6Y125_CO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_AX = CLBLM_R_X5Y125_SLICE_X6Y125_CO5;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B1 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B2 = CLBLM_R_X5Y130_SLICE_X7Y130_BQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B4 = CLBLM_L_X8Y124_SLICE_X10Y124_BQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_B6 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C1 = CLBLL_L_X4Y123_SLICE_X4Y123_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C3 = CLBLM_R_X11Y125_SLICE_X14Y125_BQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C4 = CLBLM_L_X8Y122_SLICE_X10Y122_A5Q;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_C6 = 1'b1;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D1 = CLBLM_L_X12Y127_SLICE_X17Y127_BO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D2 = CLBLM_R_X11Y127_SLICE_X15Y127_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D1 = CLBLL_L_X4Y120_SLICE_X5Y120_BQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D2 = CLBLM_R_X3Y122_SLICE_X3Y122_CO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D3 = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D4 = CLBLM_R_X5Y123_SLICE_X7Y123_BQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D5 = CLBLL_L_X4Y120_SLICE_X5Y120_AQ;
  assign CLBLM_R_X5Y125_SLICE_X6Y125_D6 = CLBLM_R_X3Y122_SLICE_X2Y122_CQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D3 = CLBLM_L_X10Y127_SLICE_X13Y127_BQ;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D5 = CLBLM_L_X10Y129_SLICE_X13Y129_CO6;
  assign CLBLM_R_X11Y127_SLICE_X15Y127_D6 = CLBLM_R_X11Y128_SLICE_X14Y128_AO5;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C2 = CLBLM_R_X3Y126_SLICE_X2Y126_AQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C3 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C4 = CLBLM_R_X7Y129_SLICE_X9Y129_BQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C5 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B3 = CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B4 = CLBLM_R_X11Y128_SLICE_X15Y128_AQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B5 = CLBLM_R_X11Y126_SLICE_X14Y126_BQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_B6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D2 = CLBLM_R_X7Y129_SLICE_X9Y129_CQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C4 = CLBLM_R_X11Y130_SLICE_X14Y130_AQ;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C5 = CLBLM_R_X11Y127_SLICE_X14Y127_DO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D6 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_C6 = CLBLM_R_X11Y127_SLICE_X14Y127_BO6;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D3 = CLBLM_L_X10Y127_SLICE_X12Y127_AQ;
  assign LIOB33_X0Y141_IOB_X0Y142_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOB33_X0Y141_IOB_X0Y141_O = CLBLL_L_X2Y126_SLICE_X1Y126_AQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A1 = CLBLM_R_X5Y128_SLICE_X7Y128_A5Q;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A2 = CLBLL_L_X4Y124_SLICE_X4Y124_BQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A4 = CLBLM_L_X8Y127_SLICE_X10Y127_AQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A5 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A6 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X13Y121_D6 = CLBLM_R_X11Y121_SLICE_X14Y121_CQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B1 = CLBLL_L_X2Y122_SLICE_X1Y122_A5Q;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B2 = CLBLM_R_X5Y126_SLICE_X7Y126_BQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B4 = CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B5 = CLBLM_L_X10Y128_SLICE_X13Y128_AQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B6 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C4 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C5 = CLBLM_R_X7Y122_SLICE_X9Y122_BQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C6 = 1'b1;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D1 = CLBLM_L_X10Y128_SLICE_X12Y128_AQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D2 = CLBLM_L_X8Y129_SLICE_X11Y129_BQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D1 = CLBLM_R_X5Y130_SLICE_X7Y130_CO5;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D2 = CLBLM_R_X5Y125_SLICE_X7Y125_CO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D3 = CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D4 = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D5 = CLBLM_R_X5Y120_SLICE_X7Y120_AQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D6 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLM_R_X11Y127_SLICE_X14Y127_D5 = CLBLM_L_X10Y129_SLICE_X12Y129_AQ;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1 = CLBLL_L_X2Y118_SLICE_X0Y118_AO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A1 = CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A3 = CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A4 = CLBLL_L_X4Y117_SLICE_X4Y117_AO5;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A6 = CLBLL_L_X4Y126_SLICE_X4Y126_DO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_A3 = CLBLM_L_X10Y121_SLICE_X12Y121_AQ;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B1 = CLBLM_R_X3Y124_SLICE_X2Y124_BQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B2 = CLBLM_R_X5Y126_SLICE_X6Y126_BQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B3 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B4 = CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B6 = CLBLM_L_X8Y127_SLICE_X10Y127_BQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C2 = CLBLM_R_X5Y126_SLICE_X6Y126_CQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C3 = CLBLM_R_X7Y120_SLICE_X8Y120_DQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C4 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C5 = CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C6 = CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B5 = CLBLM_R_X7Y131_SLICE_X9Y131_BO5;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D2 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D3 = CLBLM_R_X5Y126_SLICE_X6Y126_DQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D4 = CLBLM_L_X10Y128_SLICE_X12Y128_BQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D5 = CLBLM_R_X5Y123_SLICE_X7Y123_C5Q;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D6 = CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B6 = CLBLM_R_X7Y129_SLICE_X9Y129_CQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_C6 = 1'b1;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B2 = CLBLM_L_X10Y121_SLICE_X12Y121_BQ;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B3 = CLBLM_L_X8Y123_SLICE_X10Y123_DO6;
  assign CLBLM_L_X10Y121_SLICE_X12Y121_B4 = CLBLM_R_X11Y121_SLICE_X14Y121_CQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C3 = CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C4 = CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C6 = 1'b1;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D4 = CLBLM_L_X8Y125_SLICE_X11Y125_BQ;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D5 = CLBLM_L_X8Y124_SLICE_X10Y124_BQ;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_D1 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_L_X8Y123_SLICE_X11Y123_D6 = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_T1 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_D1 = CLBLM_R_X103Y175_SLICE_X163Y175_AO6;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_D1 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D2 = CLBLM_L_X10Y129_SLICE_X13Y129_DO6;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_T1 = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_T1 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_D1 = CLBLM_R_X103Y175_SLICE_X163Y175_AO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D5 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1 = CLBLM_R_X103Y171_SLICE_X163Y171_AO6;
  assign RIOB33_X105Y187_IOB_X1Y188_O = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1 = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign LIOB33_X0Y143_IOB_X0Y143_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_L_X8Y123_SLICE_X10Y123_B4 = CLBLM_R_X7Y122_SLICE_X9Y122_CQ;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A1 = CLBLL_L_X4Y122_SLICE_X5Y122_AQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A2 = CLBLM_L_X8Y125_SLICE_X10Y125_DQ;
  assign CLBLM_L_X8Y129_SLICE_X10Y129_D5 = CLBLM_L_X8Y128_SLICE_X10Y128_AQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A3 = CLBLM_R_X5Y127_SLICE_X7Y127_AQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A4 = CLBLM_R_X5Y124_SLICE_X6Y124_AQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B1 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B2 = CLBLL_L_X4Y124_SLICE_X4Y124_AQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B4 = CLBLM_L_X8Y125_SLICE_X10Y125_DQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B5 = CLBLM_L_X10Y127_SLICE_X13Y127_AQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B6 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C2 = CLBLM_R_X5Y127_SLICE_X7Y127_CQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C3 = CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C4 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C5 = CLBLM_R_X5Y127_SLICE_X7Y127_B5Q;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C6 = CLBLL_L_X2Y119_SLICE_X1Y119_BO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D2 = CLBLM_R_X7Y127_SLICE_X8Y127_BQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D4 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A1 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A2 = CLBLM_R_X5Y126_SLICE_X7Y126_CO5;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A3 = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A4 = CLBLM_L_X10Y127_SLICE_X13Y127_AQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A6 = CLBLM_R_X5Y122_SLICE_X6Y122_BQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B1 = CLBLM_R_X5Y121_SLICE_X6Y121_BQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B2 = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B3 = CLBLM_R_X5Y126_SLICE_X7Y126_CO5;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B4 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B6 = CLBLL_L_X4Y119_SLICE_X5Y119_AQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C2 = CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C3 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C4 = CLBLM_R_X5Y128_SLICE_X7Y128_A5Q;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C5 = CLBLM_R_X5Y126_SLICE_X7Y126_CO5;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C6 = CLBLM_R_X5Y120_SLICE_X6Y120_CQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D2 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D4 = CLBLM_R_X5Y126_SLICE_X6Y126_CQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign RIOB33_X105Y179_IOB_X1Y180_O = CLBLM_R_X11Y124_SLICE_X14Y124_DO6;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOB33_X105Y179_IOB_X1Y179_O = CLBLM_L_X10Y136_SLICE_X12Y136_AO5;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_D = RIOB33_X105Y135_IOB_X1Y136_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_D = RIOB33_X105Y135_IOB_X1Y135_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C1 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C4 = 1'b1;
  assign CLBLL_L_X4Y124_SLICE_X4Y124_D5 = 1'b1;
  assign CLBLM_L_X10Y117_SLICE_X13Y117_C6 = 1'b1;
  assign LIOB33_X0Y145_IOB_X0Y146_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOB33_X0Y145_IOB_X0Y145_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A1 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A2 = CLBLM_L_X8Y128_SLICE_X11Y128_CQ;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A4 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A5 = CLBLL_L_X2Y119_SLICE_X1Y119_AQ;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B1 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B2 = CLBLM_R_X11Y129_SLICE_X14Y129_AQ;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B3 = CLBLM_R_X3Y129_SLICE_X2Y129_AQ;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B4 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B6 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A1 = CLBLM_L_X8Y123_SLICE_X11Y123_CQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B2 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A3 = CLBLM_R_X3Y118_SLICE_X3Y118_AQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A4 = CLBLL_L_X2Y125_SLICE_X1Y125_BQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_A6 = CLBLM_R_X3Y118_SLICE_X3Y118_CO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C1 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B1 = CLBLM_L_X8Y123_SLICE_X11Y123_CQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B2 = CLBLM_R_X3Y118_SLICE_X3Y118_BQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B4 = CLBLM_L_X10Y125_SLICE_X13Y125_BQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B4 = CLBLL_L_X4Y118_SLICE_X5Y118_AQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B5 = CLBLM_R_X3Y118_SLICE_X3Y118_CO5;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C1 = CLBLL_L_X4Y118_SLICE_X5Y118_BQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C2 = CLBLL_L_X4Y119_SLICE_X4Y119_BQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B6 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C3 = CLBLM_R_X3Y118_SLICE_X3Y118_BQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C4 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C5 = CLBLM_R_X3Y118_SLICE_X3Y118_AQ;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_C6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A1 = CLBLM_L_X8Y129_SLICE_X11Y129_B5Q;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A2 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A3 = CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A4 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D1 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D2 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D3 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D4 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D5 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X3Y118_D6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A6 = CLBLL_L_X2Y121_SLICE_X0Y121_A5Q;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_AX = CLBLM_R_X5Y128_SLICE_X6Y128_CO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B1 = CLBLL_L_X4Y119_SLICE_X5Y119_CQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B2 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C1 = CLBLL_L_X2Y130_SLICE_X0Y130_AO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A1 = CLBLM_R_X3Y119_SLICE_X2Y119_CO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A2 = CLBLM_R_X5Y119_SLICE_X7Y119_CQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A3 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A4 = CLBLM_R_X3Y118_SLICE_X2Y118_BO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C2 = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A5 = CLBLM_R_X3Y118_SLICE_X2Y118_CO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C3 = CLBLL_L_X2Y130_SLICE_X0Y130_CO5;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B1 = CLBLL_L_X2Y119_SLICE_X1Y119_AQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B2 = CLBLM_R_X3Y119_SLICE_X2Y119_BQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B3 = CLBLM_R_X3Y118_SLICE_X2Y118_AQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C4 = CLBLL_L_X2Y128_SLICE_X1Y128_AO5;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B5 = CLBLM_R_X3Y119_SLICE_X2Y119_AQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_B6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C5 = CLBLM_R_X7Y128_SLICE_X8Y128_DQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C1 = CLBLM_R_X3Y119_SLICE_X2Y119_AQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C2 = CLBLL_L_X2Y119_SLICE_X1Y119_AQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C3 = CLBLM_R_X5Y118_SLICE_X7Y118_CO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C6 = CLBLM_R_X3Y121_SLICE_X2Y121_BQ;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C4 = CLBLM_R_X7Y117_SLICE_X9Y117_DO6;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C5 = CLBLM_R_X3Y119_SLICE_X3Y119_BO5;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_C6 = CLBLM_R_X3Y119_SLICE_X2Y119_BQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D3 = CLBLM_R_X5Y128_SLICE_X6Y128_DQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D4 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D6 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D1 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D2 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D3 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D4 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D5 = 1'b1;
  assign CLBLM_R_X3Y118_SLICE_X2Y118_D6 = 1'b1;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D1 = CLBLL_L_X4Y129_SLICE_X4Y129_BO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D2 = CLBLL_L_X4Y129_SLICE_X4Y129_CO6;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D3 = CLBLM_R_X7Y125_SLICE_X8Y125_DQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D4 = CLBLL_L_X4Y129_SLICE_X5Y129_CO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D5 = CLBLM_R_X5Y128_SLICE_X7Y128_DO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D6 = CLBLL_L_X4Y129_SLICE_X5Y129_BO6;
endmodule
