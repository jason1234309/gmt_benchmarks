module top(
  input LIOB33_SING_X0Y50_IOB_X0Y50_IPAD,
  input LIOB33_X0Y51_IOB_X0Y51_IPAD,
  input LIOB33_X0Y51_IOB_X0Y52_IPAD,
  input LIOB33_X0Y53_IOB_X0Y53_IPAD,
  input LIOB33_X0Y53_IOB_X0Y54_IPAD,
  input LIOB33_X0Y55_IOB_X0Y55_IPAD,
  input LIOB33_X0Y55_IOB_X0Y56_IPAD,
  input LIOB33_X0Y57_IOB_X0Y57_IPAD,
  input LIOB33_X0Y57_IOB_X0Y58_IPAD,
  input LIOB33_X0Y59_IOB_X0Y59_IPAD,
  input LIOB33_X0Y59_IOB_X0Y60_IPAD,
  input LIOB33_X0Y61_IOB_X0Y61_IPAD,
  input LIOB33_X0Y61_IOB_X0Y62_IPAD,
  input LIOB33_X0Y63_IOB_X0Y63_IPAD,
  input LIOB33_X0Y77_IOB_X0Y78_IPAD,
  input RIOB33_SING_X105Y100_IOB_X1Y100_IPAD,
  input RIOB33_SING_X105Y149_IOB_X1Y149_IPAD,
  input RIOB33_X105Y101_IOB_X1Y101_IPAD,
  input RIOB33_X105Y101_IOB_X1Y102_IPAD,
  input RIOB33_X105Y103_IOB_X1Y103_IPAD,
  input RIOB33_X105Y103_IOB_X1Y104_IPAD,
  input RIOB33_X105Y105_IOB_X1Y105_IPAD,
  input RIOB33_X105Y105_IOB_X1Y106_IPAD,
  input RIOB33_X105Y107_IOB_X1Y107_IPAD,
  input RIOB33_X105Y107_IOB_X1Y108_IPAD,
  input RIOB33_X105Y109_IOB_X1Y109_IPAD,
  input RIOB33_X105Y109_IOB_X1Y110_IPAD,
  input RIOB33_X105Y111_IOB_X1Y111_IPAD,
  input RIOB33_X105Y111_IOB_X1Y112_IPAD,
  input RIOB33_X105Y113_IOB_X1Y113_IPAD,
  input RIOB33_X105Y113_IOB_X1Y114_IPAD,
  input RIOB33_X105Y115_IOB_X1Y115_IPAD,
  input RIOB33_X105Y115_IOB_X1Y116_IPAD,
  input RIOB33_X105Y117_IOB_X1Y117_IPAD,
  input RIOB33_X105Y117_IOB_X1Y118_IPAD,
  input RIOB33_X105Y119_IOB_X1Y119_IPAD,
  input RIOB33_X105Y119_IOB_X1Y120_IPAD,
  input RIOB33_X105Y121_IOB_X1Y121_IPAD,
  input RIOB33_X105Y121_IOB_X1Y122_IPAD,
  input RIOB33_X105Y123_IOB_X1Y123_IPAD,
  input RIOB33_X105Y123_IOB_X1Y124_IPAD,
  input RIOB33_X105Y125_IOB_X1Y125_IPAD,
  input RIOB33_X105Y125_IOB_X1Y126_IPAD,
  input RIOB33_X105Y127_IOB_X1Y127_IPAD,
  input RIOB33_X105Y127_IOB_X1Y128_IPAD,
  input RIOB33_X105Y129_IOB_X1Y129_IPAD,
  input RIOB33_X105Y129_IOB_X1Y130_IPAD,
  input RIOB33_X105Y131_IOB_X1Y131_IPAD,
  input RIOB33_X105Y131_IOB_X1Y132_IPAD,
  input RIOB33_X105Y133_IOB_X1Y133_IPAD,
  input RIOB33_X105Y133_IOB_X1Y134_IPAD,
  input RIOB33_X105Y135_IOB_X1Y135_IPAD,
  input RIOB33_X105Y135_IOB_X1Y136_IPAD,
  input RIOB33_X105Y137_IOB_X1Y137_IPAD,
  input RIOB33_X105Y137_IOB_X1Y138_IPAD,
  input RIOB33_X105Y139_IOB_X1Y139_IPAD,
  input RIOB33_X105Y139_IOB_X1Y140_IPAD,
  input RIOB33_X105Y141_IOB_X1Y141_IPAD,
  input RIOB33_X105Y141_IOB_X1Y142_IPAD,
  input RIOB33_X105Y143_IOB_X1Y143_IPAD,
  input RIOB33_X105Y143_IOB_X1Y144_IPAD,
  input RIOB33_X105Y145_IOB_X1Y145_IPAD,
  input RIOB33_X105Y145_IOB_X1Y146_IPAD,
  input RIOB33_X105Y147_IOB_X1Y147_IPAD,
  input RIOB33_X105Y147_IOB_X1Y148_IPAD,
  output LIOB33_SING_X0Y100_IOB_X0Y100_OPAD,
  output LIOB33_SING_X0Y149_IOB_X0Y149_OPAD,
  output LIOB33_SING_X0Y150_IOB_X0Y150_OPAD,
  output LIOB33_SING_X0Y199_IOB_X0Y199_OPAD,
  output LIOB33_X0Y101_IOB_X0Y101_OPAD,
  output LIOB33_X0Y101_IOB_X0Y102_OPAD,
  output LIOB33_X0Y103_IOB_X0Y103_OPAD,
  output LIOB33_X0Y103_IOB_X0Y104_OPAD,
  output LIOB33_X0Y105_IOB_X0Y105_OPAD,
  output LIOB33_X0Y105_IOB_X0Y106_OPAD,
  output LIOB33_X0Y107_IOB_X0Y107_OPAD,
  output LIOB33_X0Y107_IOB_X0Y108_OPAD,
  output LIOB33_X0Y109_IOB_X0Y109_OPAD,
  output LIOB33_X0Y109_IOB_X0Y110_OPAD,
  output LIOB33_X0Y111_IOB_X0Y111_OPAD,
  output LIOB33_X0Y111_IOB_X0Y112_OPAD,
  output LIOB33_X0Y113_IOB_X0Y113_OPAD,
  output LIOB33_X0Y113_IOB_X0Y114_OPAD,
  output LIOB33_X0Y115_IOB_X0Y115_OPAD,
  output LIOB33_X0Y115_IOB_X0Y116_OPAD,
  output LIOB33_X0Y117_IOB_X0Y117_OPAD,
  output LIOB33_X0Y117_IOB_X0Y118_OPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD,
  output LIOB33_X0Y125_IOB_X0Y125_OPAD,
  output LIOB33_X0Y125_IOB_X0Y126_OPAD,
  output LIOB33_X0Y127_IOB_X0Y127_OPAD,
  output LIOB33_X0Y127_IOB_X0Y128_OPAD,
  output LIOB33_X0Y129_IOB_X0Y129_OPAD,
  output LIOB33_X0Y129_IOB_X0Y130_OPAD,
  output LIOB33_X0Y131_IOB_X0Y131_OPAD,
  output LIOB33_X0Y131_IOB_X0Y132_OPAD,
  output LIOB33_X0Y133_IOB_X0Y133_OPAD,
  output LIOB33_X0Y133_IOB_X0Y134_OPAD,
  output LIOB33_X0Y135_IOB_X0Y135_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output LIOB33_X0Y141_IOB_X0Y141_OPAD,
  output LIOB33_X0Y141_IOB_X0Y142_OPAD,
  output LIOB33_X0Y143_IOB_X0Y143_OPAD,
  output LIOB33_X0Y145_IOB_X0Y145_OPAD,
  output LIOB33_X0Y145_IOB_X0Y146_OPAD,
  output LIOB33_X0Y147_IOB_X0Y147_OPAD,
  output LIOB33_X0Y147_IOB_X0Y148_OPAD,
  output LIOB33_X0Y151_IOB_X0Y151_OPAD,
  output LIOB33_X0Y151_IOB_X0Y152_OPAD,
  output LIOB33_X0Y153_IOB_X0Y153_OPAD,
  output LIOB33_X0Y153_IOB_X0Y154_OPAD,
  output LIOB33_X0Y155_IOB_X0Y155_OPAD,
  output LIOB33_X0Y155_IOB_X0Y156_OPAD,
  output LIOB33_X0Y157_IOB_X0Y157_OPAD,
  output LIOB33_X0Y157_IOB_X0Y158_OPAD,
  output LIOB33_X0Y159_IOB_X0Y159_OPAD,
  output LIOB33_X0Y159_IOB_X0Y160_OPAD,
  output LIOB33_X0Y161_IOB_X0Y161_OPAD,
  output LIOB33_X0Y161_IOB_X0Y162_OPAD,
  output LIOB33_X0Y163_IOB_X0Y163_OPAD,
  output LIOB33_X0Y163_IOB_X0Y164_OPAD,
  output LIOB33_X0Y165_IOB_X0Y165_OPAD,
  output LIOB33_X0Y165_IOB_X0Y166_OPAD,
  output LIOB33_X0Y167_IOB_X0Y167_OPAD,
  output LIOB33_X0Y167_IOB_X0Y168_OPAD,
  output LIOB33_X0Y169_IOB_X0Y169_OPAD,
  output LIOB33_X0Y169_IOB_X0Y170_OPAD,
  output LIOB33_X0Y171_IOB_X0Y171_OPAD,
  output LIOB33_X0Y171_IOB_X0Y172_OPAD,
  output LIOB33_X0Y173_IOB_X0Y173_OPAD,
  output LIOB33_X0Y173_IOB_X0Y174_OPAD,
  output LIOB33_X0Y175_IOB_X0Y175_OPAD,
  output LIOB33_X0Y175_IOB_X0Y176_OPAD,
  output LIOB33_X0Y177_IOB_X0Y177_OPAD,
  output LIOB33_X0Y177_IOB_X0Y178_OPAD,
  output LIOB33_X0Y179_IOB_X0Y179_OPAD,
  output LIOB33_X0Y179_IOB_X0Y180_OPAD,
  output LIOB33_X0Y181_IOB_X0Y181_OPAD,
  output LIOB33_X0Y181_IOB_X0Y182_OPAD,
  output LIOB33_X0Y183_IOB_X0Y183_OPAD,
  output LIOB33_X0Y183_IOB_X0Y184_OPAD,
  output LIOB33_X0Y185_IOB_X0Y185_OPAD,
  output LIOB33_X0Y185_IOB_X0Y186_OPAD,
  output LIOB33_X0Y187_IOB_X0Y187_OPAD,
  output LIOB33_X0Y187_IOB_X0Y188_OPAD,
  output LIOB33_X0Y189_IOB_X0Y189_OPAD,
  output LIOB33_X0Y189_IOB_X0Y190_OPAD,
  output LIOB33_X0Y191_IOB_X0Y191_OPAD,
  output LIOB33_X0Y191_IOB_X0Y192_OPAD,
  output LIOB33_X0Y193_IOB_X0Y193_OPAD,
  output LIOB33_X0Y193_IOB_X0Y194_OPAD,
  output LIOB33_X0Y195_IOB_X0Y195_OPAD,
  output LIOB33_X0Y195_IOB_X0Y196_OPAD,
  output LIOB33_X0Y197_IOB_X0Y197_OPAD,
  output LIOB33_X0Y197_IOB_X0Y198_OPAD,
  output LIOB33_X0Y63_IOB_X0Y64_OPAD,
  output LIOB33_X0Y65_IOB_X0Y65_OPAD,
  output LIOB33_X0Y65_IOB_X0Y66_OPAD,
  output RIOB33_SING_X105Y150_IOB_X1Y150_OPAD,
  output RIOB33_SING_X105Y199_IOB_X1Y199_OPAD,
  output RIOB33_X105Y151_IOB_X1Y151_OPAD,
  output RIOB33_X105Y151_IOB_X1Y152_OPAD,
  output RIOB33_X105Y153_IOB_X1Y153_OPAD,
  output RIOB33_X105Y153_IOB_X1Y154_OPAD,
  output RIOB33_X105Y155_IOB_X1Y155_OPAD,
  output RIOB33_X105Y155_IOB_X1Y156_OPAD,
  output RIOB33_X105Y157_IOB_X1Y157_OPAD,
  output RIOB33_X105Y157_IOB_X1Y158_OPAD,
  output RIOB33_X105Y159_IOB_X1Y159_OPAD,
  output RIOB33_X105Y159_IOB_X1Y160_OPAD,
  output RIOB33_X105Y161_IOB_X1Y161_OPAD,
  output RIOB33_X105Y161_IOB_X1Y162_OPAD,
  output RIOB33_X105Y163_IOB_X1Y163_OPAD,
  output RIOB33_X105Y163_IOB_X1Y164_OPAD,
  output RIOB33_X105Y165_IOB_X1Y165_OPAD,
  output RIOB33_X105Y165_IOB_X1Y166_OPAD,
  output RIOB33_X105Y167_IOB_X1Y167_OPAD,
  output RIOB33_X105Y167_IOB_X1Y168_OPAD,
  output RIOB33_X105Y169_IOB_X1Y169_OPAD,
  output RIOB33_X105Y169_IOB_X1Y170_OPAD,
  output RIOB33_X105Y171_IOB_X1Y171_OPAD,
  output RIOB33_X105Y171_IOB_X1Y172_OPAD,
  output RIOB33_X105Y173_IOB_X1Y173_OPAD,
  output RIOB33_X105Y173_IOB_X1Y174_OPAD,
  output RIOB33_X105Y175_IOB_X1Y175_OPAD,
  output RIOB33_X105Y175_IOB_X1Y176_OPAD,
  output RIOB33_X105Y177_IOB_X1Y177_OPAD,
  output RIOB33_X105Y177_IOB_X1Y178_OPAD,
  output RIOB33_X105Y179_IOB_X1Y179_OPAD,
  output RIOB33_X105Y179_IOB_X1Y180_OPAD,
  output RIOB33_X105Y181_IOB_X1Y181_OPAD,
  output RIOB33_X105Y181_IOB_X1Y182_OPAD,
  output RIOB33_X105Y183_IOB_X1Y183_OPAD,
  output RIOB33_X105Y183_IOB_X1Y184_OPAD,
  output RIOB33_X105Y185_IOB_X1Y185_OPAD,
  output RIOB33_X105Y185_IOB_X1Y186_OPAD,
  output RIOB33_X105Y187_IOB_X1Y187_OPAD,
  output RIOB33_X105Y187_IOB_X1Y188_OPAD,
  output RIOB33_X105Y189_IOB_X1Y189_OPAD,
  output RIOB33_X105Y189_IOB_X1Y190_OPAD,
  output RIOB33_X105Y191_IOB_X1Y191_OPAD,
  output RIOB33_X105Y191_IOB_X1Y192_OPAD,
  output RIOB33_X105Y193_IOB_X1Y193_OPAD,
  output RIOB33_X105Y193_IOB_X1Y194_OPAD,
  output RIOB33_X105Y195_IOB_X1Y195_OPAD,
  output RIOB33_X105Y195_IOB_X1Y196_OPAD,
  output RIOB33_X105Y197_IOB_X1Y197_OPAD,
  output RIOB33_X105Y197_IOB_X1Y198_OPAD
  );
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_AO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_AO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_A_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_BO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_BO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_B_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_CO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_CO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_C_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_DO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_DO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X0Y133_D_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_AO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_AO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_A_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_BO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_BO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_B_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_CO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_CO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_C_XOR;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D1;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D2;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D3;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D4;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_DO5;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_DO6;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D_CY;
  wire [0:0] CLBLL_L_X2Y133_SLICE_X1Y133_D_XOR;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_A;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_A1;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_A2;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_A3;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_A4;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_A5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_A6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_AO5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_AO6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_A_CY;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_A_XOR;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_B;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_B1;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_B2;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_B3;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_B4;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_B5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_B6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_BO5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_BO6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_B_CY;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_B_XOR;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_C;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_C1;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_C2;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_C3;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_C4;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_C5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_C6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_CO5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_CO6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_C_CY;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_C_XOR;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_D;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_D1;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_D2;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_D3;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_D4;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_D5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_D6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_DO5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_DO6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_D_CY;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X0Y134_D_XOR;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_A;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_A1;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_A2;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_A3;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_A4;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_A5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_A6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_AMUX;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_AO5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_AO6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_A_CY;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_A_XOR;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_B;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_B1;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_B2;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_B3;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_B4;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_B5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_B6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_BO5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_BO6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_B_CY;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_B_XOR;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_C;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_C1;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_C2;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_C3;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_C4;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_C5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_C6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_CO5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_CO6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_C_CY;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_C_XOR;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_D;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_D1;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_D2;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_D3;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_D4;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_D5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_D6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_DO5;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_DO6;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_D_CY;
  wire [0:0] CLBLL_L_X2Y134_SLICE_X1Y134_D_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_AO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_AO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_A_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_BO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_BO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_B_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_CO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_CO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_C_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_DO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_DO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X0Y138_D_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_AMUX;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_AO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_AO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_A_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_BO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_BO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_B_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_CO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_CO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_C_XOR;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D1;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D2;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D3;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D4;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_DO5;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_DO6;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D_CY;
  wire [0:0] CLBLL_L_X2Y138_SLICE_X1Y138_D_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_AO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_AO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_A_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_BO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_BO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_B_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_CO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_CO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_C_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_DO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_DO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X0Y75_D_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_AO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_AO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_A_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_BO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_BO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_B_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_CO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_CO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_C_XOR;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D1;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D2;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D3;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D4;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_DO5;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_DO6;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D_CY;
  wire [0:0] CLBLL_L_X2Y75_SLICE_X1Y75_D_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_AO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_AO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_AQ;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_A_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_BO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_BO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_B_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_CLK;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_CO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_CO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_C_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_DO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_DO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X4Y129_D_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_AO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_AO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_A_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_BO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_BO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_B_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_CO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_CO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_C_XOR;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D1;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D2;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D3;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D4;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_DO5;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_DO6;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D_CY;
  wire [0:0] CLBLL_L_X4Y129_SLICE_X5Y129_D_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_AO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_AO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_AQ;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_A_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B5Q;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_BMUX;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_BO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_BO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_BQ;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_B_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_CLK;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_CMUX;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_CO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_CO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_C_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D5Q;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_DMUX;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_DO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_DO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_DQ;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X4Y130_D_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A5Q;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_AMUX;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_AO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_AO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_AQ;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_AX;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_A_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B5Q;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_BMUX;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_BO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_BO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_B_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_CLK;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_CMUX;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_CO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_CO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_C_XOR;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D1;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D2;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D3;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D4;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_DMUX;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_DO5;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_DO6;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D_CY;
  wire [0:0] CLBLL_L_X4Y130_SLICE_X5Y130_D_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_AO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_AO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_AQ;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_A_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_BO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_BQ;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_B_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_CLK;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_CO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_CO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_CQ;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_C_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D5Q;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_DMUX;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_DO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_DO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_DQ;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X4Y131_D_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_AO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_AO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_AQ;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_A_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B5Q;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_BMUX;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_BO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_BO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_BQ;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_B_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_CLK;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_CO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_CO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_C_XOR;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D1;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D2;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D3;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D4;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_DO5;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_DO6;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D_CY;
  wire [0:0] CLBLL_L_X4Y131_SLICE_X5Y131_D_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_AO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_AO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_AQ;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_A_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_BO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_BO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_BQ;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_B_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_CLK;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_CO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_CO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_CQ;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_C_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_DO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_DO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_DQ;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X4Y132_D_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A5Q;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_AMUX;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_AO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_AO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_A_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_BO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_BO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_BQ;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_B_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C5Q;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_CLK;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_CMUX;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_CO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_CO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_CQ;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_C_XOR;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D1;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D2;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D3;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D4;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D5Q;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_DMUX;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_DO5;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_DO6;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_DQ;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D_CY;
  wire [0:0] CLBLL_L_X4Y132_SLICE_X5Y132_D_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A5Q;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_AMUX;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_AO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_AO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_AQ;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_A_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_BMUX;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_BO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_BO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_BQ;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_B_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C5Q;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_CLK;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_CMUX;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_CO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_CO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_CQ;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_C_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D5Q;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_DMUX;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_DO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_DO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_DQ;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X4Y133_D_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_AO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_AO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_AQ;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_A_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B5Q;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_BMUX;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_BO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_BO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_BQ;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_B_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C5Q;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_CLK;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_CMUX;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_CO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_CO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_CQ;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_C_XOR;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D1;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D2;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D3;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D4;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D5Q;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_DMUX;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_DO5;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_DO6;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_DQ;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D_CY;
  wire [0:0] CLBLL_L_X4Y133_SLICE_X5Y133_D_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A5Q;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_AMUX;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_AO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_AO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_AQ;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_AX;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_A_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_BO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_BO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_BQ;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_B_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C5Q;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_CLK;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_CMUX;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_CO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_CO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_CQ;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_C_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D5Q;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_DMUX;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_DO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_DO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_DQ;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X4Y134_D_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_AO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_AO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_AQ;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_A_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_BO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_BO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_BQ;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_B_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_CLK;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_CO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_CO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_CQ;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_C_XOR;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D1;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D2;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D3;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D4;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D5Q;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_DMUX;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_DO5;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_DO6;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_DQ;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D_CY;
  wire [0:0] CLBLL_L_X4Y134_SLICE_X5Y134_D_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_AO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_AO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_AQ;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_A_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_BO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_BO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_BQ;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_B_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C5Q;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_CLK;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_CMUX;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_CO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_CO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_CQ;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_C_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D5Q;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_DMUX;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_DO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_DO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_DQ;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X4Y135_D_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_AO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_AO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_AQ;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_A_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_BO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_BO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_BQ;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_B_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C5Q;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_CLK;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_CMUX;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_CO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_CO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_CQ;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_C_XOR;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D1;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D2;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D3;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D4;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_DMUX;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_DO5;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_DO6;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D_CY;
  wire [0:0] CLBLL_L_X4Y135_SLICE_X5Y135_D_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A5Q;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_AMUX;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_AO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_AO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_AQ;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_A_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B5Q;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_BMUX;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_BO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_BO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_BQ;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_BX;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_B_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_CLK;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_CO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_CO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_CQ;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_C_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D5Q;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_DMUX;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_DO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_DO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_DQ;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X4Y136_D_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_AO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_AO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_AQ;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_A_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_BO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_BO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_BQ;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_B_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_CLK;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_CO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_CO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_CQ;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_C_XOR;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D1;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D2;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D3;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D4;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D5Q;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_DMUX;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_DO5;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_DO6;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_DQ;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D_CY;
  wire [0:0] CLBLL_L_X4Y136_SLICE_X5Y136_D_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_AO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_AO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_AQ;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_A_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_BO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_BO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_BQ;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_B_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C5Q;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_CLK;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_CMUX;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_CO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_CO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_CQ;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_C_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_DMUX;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_DO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_DO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X4Y137_D_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A5Q;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_AMUX;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_AO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_AO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_AQ;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_A_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B5Q;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_BMUX;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_BO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_BO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_BQ;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_B_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C5Q;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_CLK;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_CMUX;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_CO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_CO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_CQ;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_C_XOR;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D1;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D2;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D3;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D4;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D5Q;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_DMUX;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_DO5;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_DO6;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_DQ;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D_CY;
  wire [0:0] CLBLL_L_X4Y137_SLICE_X5Y137_D_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_AMUX;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_AO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_AO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_AQ;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_AX;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_A_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_BMUX;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_BO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_BO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_BQ;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_BX;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_B_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_CE;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_CLK;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_CO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_CO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_C_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_DO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_DO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X4Y138_D_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A5Q;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_AMUX;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_AO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_AO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_AQ;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_A_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B5Q;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_BMUX;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_BO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_BO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_BQ;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_BX;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_B_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C5Q;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_CLK;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_CMUX;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_CO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_CO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_CQ;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_CX;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_C_XOR;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D1;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D2;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D3;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D4;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D5Q;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_DMUX;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_DO5;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_DO6;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_DQ;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_DX;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D_CY;
  wire [0:0] CLBLL_L_X4Y138_SLICE_X5Y138_D_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A5Q;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_AMUX;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_AO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_AO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_A_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_BO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_BO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_BQ;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_B_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_CLK;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_CO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_CO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_CQ;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_C_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_DO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_DO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_DQ;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X4Y139_D_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_AO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_AO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_AQ;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_A_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_BO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_BO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_BQ;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_B_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C5Q;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_CLK;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_CMUX;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_CO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_CO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_CQ;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_C_XOR;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D1;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D2;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D3;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D4;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_DMUX;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_DO5;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_DO6;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D_CY;
  wire [0:0] CLBLL_L_X4Y139_SLICE_X5Y139_D_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_AMUX;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_AO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_AO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_AQ;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_AX;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_A_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_BMUX;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_BO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_BO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_B_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_CE;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_CLK;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_CMUX;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_CO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_CO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_C_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_DMUX;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_DO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_DO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X4Y140_D_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_AO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_AQ;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_A_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_BO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_BO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_BQ;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_B_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C5Q;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_CLK;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_CMUX;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_CO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_CO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_CQ;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_C_XOR;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D1;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D2;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D3;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D4;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_DO5;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_DO6;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_DQ;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D_CY;
  wire [0:0] CLBLL_L_X4Y140_SLICE_X5Y140_D_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_AO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_AO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_AQ;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_A_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_BO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_BO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_BQ;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_B_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_CLK;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_CO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_CO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_CQ;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_C_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_DO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_DO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_DQ;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X4Y141_D_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_AO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_AO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_AQ;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_A_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_BMUX;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_BO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_BO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_B_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_CLK;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_CO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_CO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_C_XOR;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D1;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D2;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D3;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D4;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_DO5;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_DO6;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D_CY;
  wire [0:0] CLBLL_L_X4Y141_SLICE_X5Y141_D_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A5Q;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_AMUX;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_AO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_AO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_AX;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_A_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_BMUX;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_BO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_BO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_B_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_CLK;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_CO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_CO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_C_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_DO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_DO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X4Y142_D_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A5Q;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_AMUX;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_AO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_AO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_AX;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_A_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_BO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_BO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_BQ;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_B_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_CLK;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_CMUX;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_CO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_CO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_C_XOR;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D1;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D2;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D3;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D4;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_DO5;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_DO6;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D_CY;
  wire [0:0] CLBLL_L_X4Y142_SLICE_X5Y142_D_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_AO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_AO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_A_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_BO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_BO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_B_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_CO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_CO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_C_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_DO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_DO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X4Y143_D_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_AO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_AO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_AQ;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_A_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_BMUX;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_BO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_BO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_B_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_CLK;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_CO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_CO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_C_XOR;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D1;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D2;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D3;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D4;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_DO5;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_DO6;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D_CY;
  wire [0:0] CLBLL_L_X4Y143_SLICE_X5Y143_D_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_AO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_AO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_A_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B5Q;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_BMUX;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_BO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_BO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_B_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C5Q;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CLK;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CMUX;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_C_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_DO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_DO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X12Y130_D_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_AO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_AO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_A_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_BO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_BO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_B_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_CO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_CO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_C_XOR;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D1;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D2;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D3;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D4;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_DO5;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_DO6;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D_CY;
  wire [0:0] CLBLM_L_X10Y130_SLICE_X13Y130_D_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_AO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_AO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_AQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_A_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_BO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_BO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_B_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C5Q;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CLK;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CMUX;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_CQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_C_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D5Q;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_DMUX;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_DO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_DO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_DQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X12Y131_D_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_AO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_AO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_AQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_A_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_BO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_BO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_BQ;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_B_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_CLK;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_CO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_CO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_C_XOR;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D1;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D2;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D3;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D4;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_DO5;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_DO6;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D_CY;
  wire [0:0] CLBLM_L_X10Y131_SLICE_X13Y131_D_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_AO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_AQ;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_A_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_BO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_BO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_BQ;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_B_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C5Q;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CLK;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CMUX;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_CQ;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_C_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_DO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X12Y132_D_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_AO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_AO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_AQ;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_A_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_BO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_B_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_CLK;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_CO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_CO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_C_XOR;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D1;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D2;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D3;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D4;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_DO5;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D_CY;
  wire [0:0] CLBLM_L_X10Y132_SLICE_X13Y132_D_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A5Q;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_AMUX;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_AO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_AO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_A_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_BO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_BO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_BQ;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_B_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_CLK;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_CO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_C_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_DO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_DO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X12Y133_D_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_AO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_AO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_AQ;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_A_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_BO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_B_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_CLK;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_CO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_CO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_C_XOR;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D1;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D2;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D3;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D4;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_DO5;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D_CY;
  wire [0:0] CLBLM_L_X10Y133_SLICE_X13Y133_D_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A5Q;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_AMUX;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_AO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_AO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_AQ;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_A_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B5Q;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_BMUX;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_BO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_BO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_BQ;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_B_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_CLK;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_CO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_CO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_C_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_DO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_DO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X12Y134_D_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A5Q;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_AMUX;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_AO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_AO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_AQ;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_A_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_BO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_BO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_B_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_CLK;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_CO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_CO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_C_XOR;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D1;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D2;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D3;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D4;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_DO5;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_DO6;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D_CY;
  wire [0:0] CLBLM_L_X10Y134_SLICE_X13Y134_D_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A5Q;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_AMUX;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_AO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_AO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_A_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B5Q;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_BMUX;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_BO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_BO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_B_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_CLK;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_CMUX;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_CO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_CO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_C_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_DO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X12Y135_D_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_AO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_AO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_AQ;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_AX;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_A_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_BO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_BO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_B_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_CLK;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_CO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_CO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_C_XOR;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D1;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D2;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D3;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D4;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_DO5;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D_CY;
  wire [0:0] CLBLM_L_X10Y135_SLICE_X13Y135_D_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_AO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_AO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_AQ;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_A_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_BO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_BO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_BQ;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_B_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C5Q;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_CLK;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_CMUX;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_CO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_CO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_CQ;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_C_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_DO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_DO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X12Y136_D_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_AO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_AO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_AQ;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_A_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_BO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_BO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_BQ;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_B_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_CLK;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_CMUX;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_CO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_CO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_C_XOR;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D1;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D2;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D3;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D4;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_DMUX;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_DO5;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_DO6;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D_CY;
  wire [0:0] CLBLM_L_X10Y136_SLICE_X13Y136_D_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_AMUX;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_AO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_AO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_AQ;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_AX;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_A_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_BO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_BO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_BQ;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_BX;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_B_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_CE;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_CLK;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_CO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_CO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_C_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_DO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_DO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X12Y137_D_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A5Q;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_AMUX;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_AO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_AO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_AQ;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_A_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_BMUX;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_BO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_BO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_B_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_CLK;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_CO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_CO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_C_XOR;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D1;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D2;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D3;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D4;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_DO5;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_DO6;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D_CY;
  wire [0:0] CLBLM_L_X10Y137_SLICE_X13Y137_D_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_AO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_AO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_A_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_BO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_BO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_BQ;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_B_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_CLK;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_CO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_CO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_C_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_DO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_DO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X12Y138_D_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_AO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_AO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_AQ;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_A_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_BO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_BO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_BQ;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_B_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_CLK;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_CO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_CO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_CQ;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_C_XOR;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D1;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D2;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D3;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D4;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_DO5;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_DO6;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_DQ;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D_CY;
  wire [0:0] CLBLM_L_X10Y138_SLICE_X13Y138_D_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_AMUX;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_AO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_AO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_AQ;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_AX;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_A_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_BO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_BO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_B_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_CE;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_CLK;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_CO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_CO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_C_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_DO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_DO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X12Y139_D_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A5Q;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_AMUX;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_AO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_AO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_AQ;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_AX;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_A_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_BO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_BO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_BQ;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_B_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_CLK;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_CO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_CO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_CQ;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_C_XOR;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D1;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D2;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D3;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D4;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_DO5;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_DO6;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D_CY;
  wire [0:0] CLBLM_L_X10Y139_SLICE_X13Y139_D_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_AO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_AO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_AQ;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_A_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_BO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_BO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_BQ;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_B_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_CLK;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_CO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_CO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_CQ;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_C_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D5Q;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_DMUX;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_DO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_DQ;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X12Y140_D_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_AO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_AO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_AQ;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_A_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B5Q;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_BMUX;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_BO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_BO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_BQ;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_B_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C5Q;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_CLK;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_CMUX;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_CO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_CO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_CQ;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_C_XOR;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D1;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D2;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D3;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D4;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D5Q;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_DMUX;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_DO5;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_DO6;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_DQ;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D_CY;
  wire [0:0] CLBLM_L_X10Y140_SLICE_X13Y140_D_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_AO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_AO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_AQ;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_A_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_BO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_BO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_BQ;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_B_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C5Q;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_CLK;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_CMUX;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_CO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_CO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_CQ;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_C_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_DMUX;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_DO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_DO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X12Y141_D_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_AO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_AO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_A_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_BO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_BO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_BQ;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_B_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_CLK;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_CO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_CO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_CQ;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_C_XOR;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D1;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D2;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D3;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D4;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_DO5;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_DQ;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D_CY;
  wire [0:0] CLBLM_L_X10Y141_SLICE_X13Y141_D_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_AO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_AO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_A_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_BMUX;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_BO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_BO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_B_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_CLK;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_CO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_CO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_C_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_DO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_DO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X12Y142_D_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_AO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_AO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_A_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_BO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_B_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_CO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_CO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_C_XOR;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D1;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D2;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D3;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D4;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_DO5;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_DO6;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D_CY;
  wire [0:0] CLBLM_L_X10Y142_SLICE_X13Y142_D_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_AO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_AO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_A_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_BO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_B_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_CO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_CO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_C_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_DO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_DO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X16Y131_D_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_AO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_AO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_A_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_BO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_B_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_CO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_CO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_C_XOR;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D1;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D2;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D3;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D4;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_DO5;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_DO6;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D_CY;
  wire [0:0] CLBLM_L_X12Y131_SLICE_X17Y131_D_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_AO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_AO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_A_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_BO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_BO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_B_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_CO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_CO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_C_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_DO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_DO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X16Y132_D_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_AO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_AO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_A_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_BO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_BO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_B_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_CO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_CO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_C_XOR;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D1;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D2;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D3;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D4;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_DO5;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_DO6;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D_CY;
  wire [0:0] CLBLM_L_X12Y132_SLICE_X17Y132_D_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_AO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_AO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_A_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_BO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_BO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_B_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_CO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_CO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_C_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_DO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_DO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X16Y133_D_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_AO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_AO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_A_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_BO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_BO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_B_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_CO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_CO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_C_XOR;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D1;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D2;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D3;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D4;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_DMUX;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_DO5;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_DO6;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D_CY;
  wire [0:0] CLBLM_L_X12Y133_SLICE_X17Y133_D_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_AMUX;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_AO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_AO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_A_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_BO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_BO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_B_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_CO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_CO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_C_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_DMUX;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_DO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_DO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X16Y134_D_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_AMUX;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_A_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_BO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_BO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_B_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_CMUX;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_CO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_CO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_C_XOR;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D1;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D2;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D3;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D4;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_DO5;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_DO6;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D_CY;
  wire [0:0] CLBLM_L_X12Y134_SLICE_X17Y134_D_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_AMUX;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_AO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_AO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_A_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_BO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_BO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_B_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_CO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_CO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_C_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_DMUX;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_DO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_DO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X16Y135_D_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_AMUX;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_AO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_AO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_A_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_BO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_BO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_B_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_CO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_CO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_C_XOR;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D1;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D2;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D3;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D4;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_DO5;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_DO6;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D_CY;
  wire [0:0] CLBLM_L_X12Y135_SLICE_X17Y135_D_XOR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A1;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A2;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A3;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A4;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A5Q;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_AMUX;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_AO5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_AO6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_AQ;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A_CY;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_A_XOR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B1;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B2;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B3;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B4;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_BO5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_BO6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B_CY;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_B_XOR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C1;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C2;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C3;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C4;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_CLK;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_CO5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_CO6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C_CY;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_C_XOR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D1;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D2;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D3;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D4;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_DO5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_DO6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D_CY;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X16Y136_D_XOR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A1;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A2;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A3;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A4;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_AMUX;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_AO5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_AO6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A_CY;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_A_XOR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B1;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B2;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B3;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B4;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_BMUX;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_BO5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_BO6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B_CY;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_B_XOR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C1;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C2;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C3;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C4;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_CMUX;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_CO5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_CO6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C_CY;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_C_XOR;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D1;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D2;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D3;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D4;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_DO5;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_DO6;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D_CY;
  wire [0:0] CLBLM_L_X12Y136_SLICE_X17Y136_D_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_AO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_AO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_A_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_BO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_BO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_B_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_CO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_CO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_C_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_DO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_DO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X16Y137_D_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_AMUX;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_AO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_AO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_A_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_BO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_BO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_B_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_CO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_CO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_C_XOR;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D1;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D2;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D3;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D4;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_DO5;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_DO6;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D_CY;
  wire [0:0] CLBLM_L_X12Y137_SLICE_X17Y137_D_XOR;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A1;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A2;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A3;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A4;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_AMUX;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_AO5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_AO6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A_CY;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_A_XOR;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B1;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B2;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B3;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B4;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_BO5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_BO6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B_CY;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_B_XOR;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C1;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C2;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C3;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C4;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_CO5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_CO6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C_CY;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_C_XOR;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D1;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D2;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D3;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D4;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_DO5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_DO6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D_CY;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X16Y138_D_XOR;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A1;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A2;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A3;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A4;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_AO5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_AO6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A_CY;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_A_XOR;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B1;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B2;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B3;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B4;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_BMUX;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_BO5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_BO6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B_CY;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_B_XOR;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C1;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C2;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C3;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C4;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_CMUX;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_CO5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_CO6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C_CY;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_C_XOR;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D1;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D2;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D3;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D4;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_DO5;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_DO6;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D_CY;
  wire [0:0] CLBLM_L_X12Y138_SLICE_X17Y138_D_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_AMUX;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_AO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_AO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_A_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_BO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_BO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_B_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_CO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_CO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_C_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_DO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_DO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X16Y139_D_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_AO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_AO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_A_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_BMUX;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_BO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_BO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_B_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_CO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_CO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_C_XOR;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D1;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D2;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D3;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D4;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_DO5;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_DO6;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D_CY;
  wire [0:0] CLBLM_L_X12Y139_SLICE_X17Y139_D_XOR;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A1;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A2;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A3;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A4;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_AMUX;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_AO5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_AO6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_AQ;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_AX;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A_CY;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_A_XOR;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B1;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B2;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B3;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B4;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_BMUX;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_BO5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_BO6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B_CY;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_B_XOR;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C1;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C2;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C3;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C4;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_CE;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_CLK;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_CMUX;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_CO5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_CO6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C_CY;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_C_XOR;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D1;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D2;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D3;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D4;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_DO5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_DO6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D_CY;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X16Y140_D_XOR;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A1;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A2;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A3;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A4;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_AO5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_AO6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A_CY;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_A_XOR;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B1;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B2;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B3;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B4;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_BO5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_BO6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B_CY;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_B_XOR;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C1;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C2;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C3;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C4;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_CO5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_CO6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C_CY;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_C_XOR;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D1;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D2;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D3;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D4;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_DO5;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_DO6;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D_CY;
  wire [0:0] CLBLM_L_X12Y140_SLICE_X17Y140_D_XOR;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A1;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A2;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A3;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A4;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_AO5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_AO6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_AQ;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A_CY;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_A_XOR;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B1;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B2;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B3;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B4;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_BMUX;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_BO5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_BO6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B_CY;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_B_XOR;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C1;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C2;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C3;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C4;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_CLK;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_CO5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_CO6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C_CY;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_C_XOR;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D1;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D2;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D3;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D4;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_DO5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_DO6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D_CY;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X16Y141_D_XOR;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A1;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A2;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A3;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A4;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_AO5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_AO6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A_CY;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_A_XOR;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B1;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B2;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B3;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B4;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_BO5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_BO6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B_CY;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_B_XOR;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C1;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C2;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C3;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C4;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_CO5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_CO6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C_CY;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_C_XOR;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D1;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D2;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D3;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D4;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_DO5;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_DO6;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D_CY;
  wire [0:0] CLBLM_L_X12Y141_SLICE_X17Y141_D_XOR;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A1;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A2;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A3;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A4;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_AMUX;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_AO5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_AO6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A_CY;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_A_XOR;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B1;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B2;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B3;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B4;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_BMUX;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_BO5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_BO6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B_CY;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_B_XOR;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C1;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C2;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C3;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C4;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_CO5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_CO6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C_CY;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_C_XOR;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D1;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D2;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D3;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D4;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_DO5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_DO6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D_CY;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X16Y142_D_XOR;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A1;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A2;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A3;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A4;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_AO5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_AO6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A_CY;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_A_XOR;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B1;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B2;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B3;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B4;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_BO5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_BO6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B_CY;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_B_XOR;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C1;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C2;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C3;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C4;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_CO5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_CO6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C_CY;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_C_XOR;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D1;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D2;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D3;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D4;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_DO5;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_DO6;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D_CY;
  wire [0:0] CLBLM_L_X12Y142_SLICE_X17Y142_D_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_AMUX;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_AO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_AO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_A_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_BO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_BO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_B_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_CO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_CO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_C_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_DO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_DO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X16Y143_D_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_AO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_AO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_A_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_BO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_BO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_B_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_CO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_CO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_C_XOR;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D1;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D2;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D3;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D4;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_DO5;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_DO6;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D_CY;
  wire [0:0] CLBLM_L_X12Y143_SLICE_X17Y143_D_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_AO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_AO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_A_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_BO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_BO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_B_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_CLK;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_CO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_CO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_C_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_DO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_DO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X10Y130_D_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_AO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_AO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_A_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_BO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_BO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_B_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_CO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_CO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_C_XOR;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D1;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D2;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D3;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D4;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_DO5;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_DO6;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D_CY;
  wire [0:0] CLBLM_L_X8Y130_SLICE_X11Y130_D_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_A_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_BO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_BO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_BQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_B_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CLK;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_CQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_C_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_DO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_DO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X10Y131_D_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_A_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_BO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_BO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_BQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_B_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C5Q;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CLK;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CMUX;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_CQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_C_XOR;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D1;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D2;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D3;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D4;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D5Q;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_DMUX;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_DO5;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_DQ;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D_CY;
  wire [0:0] CLBLM_L_X8Y131_SLICE_X11Y131_D_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A5Q;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_AMUX;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_AO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_AO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_A_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B5Q;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_BMUX;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_BO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_BO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_BQ;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_B_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_CLK;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_CO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_CO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_CQ;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_C_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_DO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_DO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X10Y132_D_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_AMUX;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_AO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_AO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_AQ;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_A_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_BO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_BO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_BQ;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_B_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_CLK;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_CO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_CO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_C_XOR;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D1;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D2;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D3;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D4;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_DMUX;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_DO5;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_DO6;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D_CY;
  wire [0:0] CLBLM_L_X8Y132_SLICE_X11Y132_D_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_AO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_AO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_AQ;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_A_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_BO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_BO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_BQ;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_B_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C5Q;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_CLK;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_CMUX;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_CO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_CO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_CQ;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_C_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_DO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_DO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X10Y133_D_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_AMUX;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_AO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_AO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_AQ;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_A_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B5Q;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_BMUX;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_BO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_BO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_BQ;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_B_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_CLK;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_CMUX;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_CO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_CO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_C_XOR;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D1;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D2;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D3;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D4;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_DO5;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_DO6;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D_CY;
  wire [0:0] CLBLM_L_X8Y133_SLICE_X11Y133_D_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A5Q;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_AMUX;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_AO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_AO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_AQ;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_A_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_BO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_BO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_B_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_CLK;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_CO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_CO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_C_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_DMUX;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_DO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_DO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X10Y134_D_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_AO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_AO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_AQ;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_A_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B5Q;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_BMUX;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_BO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_BO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_B_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_CLK;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_CO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_CO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_C_XOR;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D1;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D2;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D3;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D4;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_DO5;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_DO6;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D_CY;
  wire [0:0] CLBLM_L_X8Y134_SLICE_X11Y134_D_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_AO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_AO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_AQ;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_A_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B5Q;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_BMUX;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_BO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_BO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_BQ;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_B_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C5Q;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_CLK;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_CMUX;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_CO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_CO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_CQ;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_C_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D5Q;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_DMUX;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_DO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_DO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_DQ;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X10Y135_D_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_AO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_AO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_AQ;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_A_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_BO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_BO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_B_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_CLK;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_CO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_CO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_C_XOR;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D1;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D2;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D3;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D4;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_DO5;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_DO6;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D_CY;
  wire [0:0] CLBLM_L_X8Y135_SLICE_X11Y135_D_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_AMUX;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_AO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_AO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_AQ;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_AX;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_A_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_BO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_BO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_BQ;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_BX;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_B_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_CE;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_CLK;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_CO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_CO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_C_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_DO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_DO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X10Y136_D_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_AO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_AO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_AQ;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_A_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B5Q;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_BMUX;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_BO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_BO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_BQ;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_B_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_CLK;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_CMUX;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_CO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_CO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_C_XOR;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D1;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D2;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D3;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D4;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_DO5;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_DO6;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D_CY;
  wire [0:0] CLBLM_L_X8Y136_SLICE_X11Y136_D_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_AO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_AO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_AQ;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_A_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B5Q;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_BMUX;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_BO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_BO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_BQ;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_B_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C5Q;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_CLK;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_CMUX;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_CO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_CO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_CQ;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_C_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D5Q;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_DMUX;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_DO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_DO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_DQ;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X10Y137_D_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_AO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_AO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_AQ;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_A_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_BO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_BO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_BQ;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_B_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_CLK;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_CO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_CO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_CQ;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_C_XOR;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D1;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D2;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D3;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D4;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D5Q;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_DMUX;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_DO5;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_DO6;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_DQ;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D_CY;
  wire [0:0] CLBLM_L_X8Y137_SLICE_X11Y137_D_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A5Q;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_AMUX;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_AO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_A_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_BMUX;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_BO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_BQ;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_B_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C5Q;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_CLK;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_CMUX;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_CO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_CO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_CQ;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_C_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D5Q;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_DMUX;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_DO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_DQ;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X10Y138_D_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_AO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_AO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_AQ;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_A_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B5Q;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_BMUX;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_BO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_BO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_BQ;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_B_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C5Q;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_CLK;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_CMUX;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_CO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_CO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_CQ;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_C_XOR;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D1;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D2;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D3;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D4;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_DO5;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_DO6;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D_CY;
  wire [0:0] CLBLM_L_X8Y138_SLICE_X11Y138_D_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_AO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_AO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_AX;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_A_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_BMUX;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_BO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_BO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_B_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_CE;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_CLK;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_CO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_CO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_C_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_DO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_DO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X10Y139_D_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_AO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_AO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_A_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_BO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_BO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_BQ;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_B_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C5Q;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_CLK;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_CMUX;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_CO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_CO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_CQ;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_C_XOR;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D1;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D2;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D3;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D4;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_DO5;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D_CY;
  wire [0:0] CLBLM_L_X8Y139_SLICE_X11Y139_D_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_AO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_AO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_AQ;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_A_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_BO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_BO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_BQ;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_B_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C5Q;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_CLK;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_CMUX;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_CO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_CQ;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_C_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D5Q;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_DMUX;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_DO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X10Y140_D_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_AO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_AO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_AQ;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_A_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B5Q;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_BMUX;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_BO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_BO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_BQ;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_B_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_CLK;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_CO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_CO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_CQ;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_C_XOR;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D1;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D2;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D3;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D4;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_DO5;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_DO6;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D_CY;
  wire [0:0] CLBLM_L_X8Y140_SLICE_X11Y140_D_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_AO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_AO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_A_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_BO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_BO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_BQ;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_B_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_CLK;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_CMUX;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_CO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_CO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_C_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_DO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X10Y141_D_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_AMUX;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_AO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_AO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_AQ;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_A_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_BO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_BO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_BQ;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_B_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_CLK;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_CMUX;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_CO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_CO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_C_XOR;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D1;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D2;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D3;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D4;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_DO5;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D_CY;
  wire [0:0] CLBLM_L_X8Y141_SLICE_X11Y141_D_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A5Q;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_AMUX;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_AO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_AO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_AX;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_A_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_BMUX;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_BO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_BO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_B_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_CLK;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_CMUX;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_CO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_CO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_C_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_DO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_DO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X10Y142_D_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_AO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_AO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_AQ;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_A_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_BO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_BO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_B_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_CLK;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_CMUX;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_CO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_CO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_C_XOR;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D1;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D2;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D3;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D4;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_DO5;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_DO6;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D_CY;
  wire [0:0] CLBLM_L_X8Y142_SLICE_X11Y142_D_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_AO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_AO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_A_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_BMUX;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_BO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_BO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_B_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_CLK;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_CO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_CO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_C_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_DO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X10Y143_D_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_AO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_AO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_AQ;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_A_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_BO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_BO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_B_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_CLK;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_CO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_CO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_C_XOR;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D1;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D2;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D3;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D4;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_DO5;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_DO6;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D_CY;
  wire [0:0] CLBLM_L_X8Y143_SLICE_X11Y143_D_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_AO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_AO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_A_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_BO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_BO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_B_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_CO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_CO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_C_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_DO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_DO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X10Y144_D_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_AO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_AO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_A_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_BO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_B_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_CO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_C_XOR;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D1;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D2;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D3;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D4;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_DO5;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_DO6;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D_CY;
  wire [0:0] CLBLM_L_X8Y144_SLICE_X11Y144_D_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_AO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_AO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_A_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_BO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_BO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_B_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_CO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_CO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_C_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_DO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_DO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X162Y178_D_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_AO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_A_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_BO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_BO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_B_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_CO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_CO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_C_XOR;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D1;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D2;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D3;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D4;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_DO5;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_DO6;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D_CY;
  wire [0:0] CLBLM_R_X103Y178_SLICE_X163Y178_D_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_AMUX;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_AO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_AO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_A_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_BO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_BO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_B_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_CO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_C_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_DO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_DO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X14Y131_D_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_AO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_AO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_A_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_BO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_BO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_B_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_CO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_CO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_C_XOR;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D1;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D2;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D3;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D4;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_DO5;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_DO6;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D_CY;
  wire [0:0] CLBLM_R_X11Y131_SLICE_X15Y131_D_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_AO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_AO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_AX;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_A_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_BO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_BO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_B_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_CE;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_CLK;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_CO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_CO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_C_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_DO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_DO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X14Y132_D_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_AMUX;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_AO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_AO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_A_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_BMUX;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_BO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_BO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_B_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_CO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_CO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_C_XOR;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D1;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D2;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D3;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D4;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_DO5;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_DO6;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D_CY;
  wire [0:0] CLBLM_R_X11Y132_SLICE_X15Y132_D_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_AO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_AO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_AQ;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_A_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_BO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_BO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_BQ;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_B_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_CLK;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_CMUX;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_CO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_CO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_C_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_DMUX;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_DO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_DO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X14Y133_D_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_AO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_AO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_A_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_BO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_BO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_B_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_CO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_CO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_C_XOR;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D1;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D2;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D3;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D4;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_DO5;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_DO6;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D_CY;
  wire [0:0] CLBLM_R_X11Y133_SLICE_X15Y133_D_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_AMUX;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_AO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_AO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_A_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_BO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_BO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_B_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_CO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_CO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_C_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_DO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_DO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X14Y134_D_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_AO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_A_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_BMUX;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_BO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_B_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_CO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_CO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_C_XOR;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D1;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D2;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D3;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D4;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_DO5;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_DO6;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D_CY;
  wire [0:0] CLBLM_R_X11Y134_SLICE_X15Y134_D_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_AO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_AO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_A_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_BO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_BO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_B_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_CO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_CO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_C_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_DO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_DO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X14Y135_D_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_AO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_AO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_A_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_BO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_BO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_B_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_CO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_CO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_C_XOR;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D1;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D2;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D3;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D4;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_DO5;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_DO6;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D_CY;
  wire [0:0] CLBLM_R_X11Y135_SLICE_X15Y135_D_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_AO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_AO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_AQ;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_A_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_BO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_BO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_B_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_CLK;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_CO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_CO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_C_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_DMUX;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_DO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_DO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X14Y136_D_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_AMUX;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_AO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_AO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_AQ;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_AX;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_A_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_BO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_BO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_B_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_CE;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_CLK;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_CO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_CO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_C_XOR;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D1;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D2;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D3;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D4;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_DO5;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_DO6;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D_CY;
  wire [0:0] CLBLM_R_X11Y136_SLICE_X15Y136_D_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_AMUX;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_AO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_AO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_A_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_BO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_BO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_B_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_CO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_CO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_C_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_DO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_DO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X14Y137_D_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_AO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_AO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_A_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_BO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_BO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_B_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_CO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_CO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_C_XOR;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D1;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D2;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D3;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D4;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_DO5;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_DO6;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D_CY;
  wire [0:0] CLBLM_R_X11Y137_SLICE_X15Y137_D_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_AO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_AO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_AQ;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_AX;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_A_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_BO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_BO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_B_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_CE;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_CLK;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_CO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_CO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_C_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_DO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_DO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X14Y138_D_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_AO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_AO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_A_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_BO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_BO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_B_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_CO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_CO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_C_XOR;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D1;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D2;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D3;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D4;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_DO5;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_DO6;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D_CY;
  wire [0:0] CLBLM_R_X11Y138_SLICE_X15Y138_D_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_AMUX;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_AO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_AO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_AQ;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_AX;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_A_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_BO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_BO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_B_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_CE;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_CLK;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_CO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_CO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_C_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_DO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_DO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X14Y139_D_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_AMUX;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_AO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_AO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_A_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_BO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_BO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_B_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_CO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_CO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_C_XOR;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D1;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D2;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D3;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D4;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_DMUX;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_DO5;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_DO6;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D_CY;
  wire [0:0] CLBLM_R_X11Y139_SLICE_X15Y139_D_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_AMUX;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_AO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_AO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_AQ;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_AX;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_A_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_BMUX;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_BO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_BO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_BQ;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_BX;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_B_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_CE;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_CLK;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_CO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_CO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_CQ;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_CX;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_C_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_DO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_DO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_DQ;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_DX;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X14Y140_D_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_AO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_AO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_AQ;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_A_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B5Q;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_BMUX;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_BO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_BO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_BQ;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_B_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_CLK;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_CMUX;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_CO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_CO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_C_XOR;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D1;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D2;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D3;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D4;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_DO5;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_DO6;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D_CY;
  wire [0:0] CLBLM_R_X11Y140_SLICE_X15Y140_D_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_AO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_AO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_AQ;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_AX;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_A_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_BO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_BO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_B_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_CLK;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_CO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_CO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_C_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_DO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_DO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X14Y141_D_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_AO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_AO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_A_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_BO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_BO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_B_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_CLK;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_CO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_CO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_C_XOR;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D1;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D2;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D3;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D4;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_DO5;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_DO6;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D_CY;
  wire [0:0] CLBLM_R_X11Y141_SLICE_X15Y141_D_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_AO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_AO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_AQ;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_A_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_BO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_BO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_B_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_CLK;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_CO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_CO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_C_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_DO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_DO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X14Y142_D_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_AMUX;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_AO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_AO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_A_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_BO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_BO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_B_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_CO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_CO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_C_XOR;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D1;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D2;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D3;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D4;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_DO5;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_DO6;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D_CY;
  wire [0:0] CLBLM_R_X11Y142_SLICE_X15Y142_D_XOR;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A1;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A2;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A3;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A4;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_AO5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_AO6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A_CY;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_A_XOR;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B1;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B2;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B3;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B4;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_BO5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_BO6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B_CY;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_B_XOR;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C1;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C2;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C3;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C4;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_CO5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_CO6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C_CY;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_C_XOR;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D1;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D2;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D3;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D4;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_DMUX;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_DO5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_DO6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D_CY;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X18Y134_D_XOR;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A1;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A2;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A3;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A4;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_AO5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_AO6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A_CY;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_A_XOR;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B1;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B2;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B3;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B4;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_BO5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_BO6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B_CY;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_B_XOR;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C1;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C2;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C3;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C4;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_CO5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_CO6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C_CY;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_C_XOR;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D1;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D2;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D3;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D4;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_DO5;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_DO6;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D_CY;
  wire [0:0] CLBLM_R_X13Y134_SLICE_X19Y134_D_XOR;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_A;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_A1;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_A2;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_A3;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_A4;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_A5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_A6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_AMUX;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_AO5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_AO6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_A_CY;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_A_XOR;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_B;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_B1;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_B2;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_B3;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_B4;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_B5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_B6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_BMUX;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_BO5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_BO6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_B_CY;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_B_XOR;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_C;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_C1;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_C2;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_C3;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_C4;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_C5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_C6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_CO5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_CO6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_C_CY;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_C_XOR;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_D;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_D1;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_D2;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_D3;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_D4;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_D5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_D6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_DO5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_DO6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_D_CY;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X18Y137_D_XOR;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_A;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_A1;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_A2;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_A3;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_A4;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_A5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_A6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_AO5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_AO6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_A_CY;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_A_XOR;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_B;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_B1;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_B2;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_B3;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_B4;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_B5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_B6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_BO5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_BO6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_B_CY;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_B_XOR;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_C;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_C1;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_C2;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_C3;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_C4;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_C5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_C6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_CO5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_CO6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_C_CY;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_C_XOR;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_D;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_D1;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_D2;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_D3;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_D4;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_D5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_D6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_DO5;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_DO6;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_D_CY;
  wire [0:0] CLBLM_R_X13Y137_SLICE_X19Y137_D_XOR;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_A;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_A1;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_A2;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_A3;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_A4;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_A5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_A6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_AMUX;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_AO5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_AO6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_A_CY;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_A_XOR;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_B;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_B1;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_B2;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_B3;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_B4;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_B5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_B6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_BMUX;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_BO5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_BO6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_B_CY;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_B_XOR;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_C;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_C1;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_C2;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_C3;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_C4;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_C5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_C6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_CO5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_CO6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_C_CY;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_C_XOR;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_D;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_D1;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_D2;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_D3;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_D4;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_D5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_D6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_DO5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_DO6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_D_CY;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X18Y138_D_XOR;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_A;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_A1;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_A2;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_A3;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_A4;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_A5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_A6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_AO5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_AO6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_A_CY;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_A_XOR;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_B;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_B1;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_B2;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_B3;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_B4;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_B5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_B6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_BO5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_BO6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_B_CY;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_B_XOR;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_C;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_C1;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_C2;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_C3;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_C4;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_C5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_C6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_CO5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_CO6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_C_CY;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_C_XOR;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_D;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_D1;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_D2;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_D3;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_D4;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_D5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_D6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_DO5;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_DO6;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_D_CY;
  wire [0:0] CLBLM_R_X13Y138_SLICE_X19Y138_D_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_AO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_AO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_A_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_BO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_BO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_B_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_CO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_CO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_C_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_DO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_DO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X2Y130_D_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_AO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_AO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_A_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_BO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_BO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_B_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_CO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_CO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_C_XOR;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D1;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D2;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D3;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D4;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_DO5;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_DO6;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D_CY;
  wire [0:0] CLBLM_R_X3Y130_SLICE_X3Y130_D_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_AO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_AO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_AQ;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_A_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_BO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_BO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_BQ;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_BX;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_B_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_CLK;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_CO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_CO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_C_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_DO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_DO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X2Y131_D_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_AO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_AO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_AQ;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_A_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B5Q;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_BMUX;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_BO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_BO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_BQ;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_B_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_CLK;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_CO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_CO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_C_XOR;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D1;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D2;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D3;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D4;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_DO5;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_DO6;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D_CY;
  wire [0:0] CLBLM_R_X3Y131_SLICE_X3Y131_D_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_AO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_AO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_A_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_BO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_BO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_BQ;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_B_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_CLK;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_CMUX;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_CO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_CO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_C_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_DO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_DO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X2Y132_D_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_AO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_AO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_A_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_BO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_BO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_BQ;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_B_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_CLK;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_CO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_CO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_CQ;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_C_XOR;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D1;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D2;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D3;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D4;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D5Q;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_DMUX;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_DO5;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_DO6;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_DQ;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D_CY;
  wire [0:0] CLBLM_R_X3Y132_SLICE_X3Y132_D_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_AO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_AO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_AQ;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_A_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_BO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_BO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_BQ;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_B_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_CLK;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_CO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_CO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_C_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_DMUX;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_DO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_DO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X2Y133_D_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_AO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_AO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_A_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B5Q;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_BMUX;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_BO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_BO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_BQ;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_B_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_CLK;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_CO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_CO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_C_XOR;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D1;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D2;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D3;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D4;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_DO5;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_DO6;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D_CY;
  wire [0:0] CLBLM_R_X3Y133_SLICE_X3Y133_D_XOR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A1;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A2;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A3;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A4;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_AMUX;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_AO5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_AO6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_AQ;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_AX;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A_CY;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_A_XOR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B1;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B2;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B3;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B4;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_BO5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_BO6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B_CY;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_B_XOR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C1;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C2;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C3;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C4;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_CE;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_CLK;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_CO5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_CO6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C_CY;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_C_XOR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D1;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D2;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D3;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D4;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_DO5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_DO6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D_CY;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X2Y134_D_XOR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A1;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A2;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A3;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A4;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A5Q;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_AMUX;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_AO5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_AO6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_AQ;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A_CY;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_A_XOR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B1;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B2;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B3;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B4;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_BO5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_BO6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_BQ;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B_CY;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_B_XOR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C1;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C2;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C3;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C4;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_CLK;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_CO5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_CO6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C_CY;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_C_XOR;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D1;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D2;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D3;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D4;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_DO5;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_DO6;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D_CY;
  wire [0:0] CLBLM_R_X3Y134_SLICE_X3Y134_D_XOR;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A1;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A2;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A3;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A4;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_AO5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_AO6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_AQ;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A_CY;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_A_XOR;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B1;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B2;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B3;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B4;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_BO5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_BO6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_BQ;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B_CY;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_B_XOR;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C1;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C2;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C3;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C4;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_CLK;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_CO5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_CO6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_CQ;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C_CY;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_C_XOR;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D1;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D2;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D3;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D4;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_DO5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_DO6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_DQ;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D_CY;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X2Y135_D_XOR;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A1;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A2;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A3;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A4;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A5Q;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_AMUX;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_AO5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_AO6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_AQ;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A_CY;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_A_XOR;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B1;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B2;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B3;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B4;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_BO5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_BO6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_BQ;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B_CY;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_B_XOR;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C1;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C2;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C3;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C4;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_CLK;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_CO5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_CO6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_CQ;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C_CY;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_C_XOR;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D1;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D2;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D3;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D4;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_DO5;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_DO6;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_DQ;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D_CY;
  wire [0:0] CLBLM_R_X3Y135_SLICE_X3Y135_D_XOR;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A1;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A2;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A3;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A4;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A5Q;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_AMUX;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_AO5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_AO6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_AQ;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A_CY;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_A_XOR;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B1;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B2;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B3;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B4;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B5Q;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_BMUX;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_BO5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_BO6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_BQ;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B_CY;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_B_XOR;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C1;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C2;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C3;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C4;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_CLK;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_CO5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_CO6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_CQ;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C_CY;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_C_XOR;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D1;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D2;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D3;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D4;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_DO5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_DO6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_DQ;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D_CY;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X2Y136_D_XOR;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A1;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A2;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A3;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A4;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_AO5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_AO6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_AQ;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A_CY;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_A_XOR;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B1;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B2;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B3;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B4;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B5Q;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_BMUX;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_BO5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_BO6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B_CY;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_B_XOR;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C1;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C2;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C3;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C4;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C5Q;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_CLK;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_CMUX;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_CO5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_CO6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_CQ;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C_CY;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_C_XOR;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D1;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D2;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D3;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D4;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D5Q;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_DMUX;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_DO5;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_DO6;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_DQ;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D_CY;
  wire [0:0] CLBLM_R_X3Y136_SLICE_X3Y136_D_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_AO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_AO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_AQ;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_A_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_BO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_BO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_B_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_CLK;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_CO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_CO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_C_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_DO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_DO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X2Y137_D_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A5Q;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_AMUX;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_AO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_AO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_AQ;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_A_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B5Q;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_BMUX;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_BO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_BO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_BQ;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_B_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C5Q;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_CLK;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_CMUX;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_CO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_CO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_CQ;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_C_XOR;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D1;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D2;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D3;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D4;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D5Q;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_DMUX;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_DO5;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_DO6;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_DQ;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D_CY;
  wire [0:0] CLBLM_R_X3Y137_SLICE_X3Y137_D_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_AO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_AO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_AQ;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_A_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_BO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_BO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_BQ;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_B_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_CLK;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_CO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_CO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_CQ;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_C_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_DO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_DO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X2Y138_D_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A5Q;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_AMUX;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_AO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_AO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_AQ;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_A_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_BMUX;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_BO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_BO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_B_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_CLK;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_CO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_CO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_C_XOR;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D1;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D2;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D3;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D4;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_DO5;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_DO6;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D_CY;
  wire [0:0] CLBLM_R_X3Y138_SLICE_X3Y138_D_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_AO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_AO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_AQ;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_A_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_BO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_BO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_BQ;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_B_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C5Q;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_CLK;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_CMUX;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_CO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_CO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_CQ;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_C_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_DO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_DO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X2Y139_D_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A5Q;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_AMUX;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_AO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_AO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_AQ;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_A_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_BO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_BO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_BQ;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_BX;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_B_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_CLK;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_CO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_CO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_C_XOR;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D1;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D2;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D3;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D4;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_DO5;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_DO6;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D_CY;
  wire [0:0] CLBLM_R_X3Y139_SLICE_X3Y139_D_XOR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A1;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A2;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A3;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A4;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_AO5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_AO6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A_CY;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_A_XOR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B1;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B2;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B3;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B4;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_BO5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_BO6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B_CY;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_B_XOR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C1;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C2;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C3;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C4;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_CO5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_CO6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C_CY;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_C_XOR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D1;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D2;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D3;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D4;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_DO5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_DO6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D_CY;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X2Y140_D_XOR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A1;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A2;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A3;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A4;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_AO5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_AO6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_AQ;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A_CY;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_A_XOR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B1;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B2;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B3;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B4;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_BO5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_BO6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_BQ;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B_CY;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_B_XOR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C1;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C2;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C3;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C4;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C5Q;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_CLK;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_CMUX;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_CO5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_CO6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_CQ;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C_CY;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_C_XOR;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D1;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D2;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D3;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D4;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_DO5;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_DO6;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_DQ;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D_CY;
  wire [0:0] CLBLM_R_X3Y140_SLICE_X3Y140_D_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_AMUX;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_AO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_AO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_AQ;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_AX;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_A_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_BMUX;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_BO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_BO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_BQ;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_BX;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_B_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_CLK;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_CO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_CO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_C_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_DO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_DO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X2Y141_D_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_AMUX;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_AO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_AO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_A_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_BO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_BO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_B_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_CO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_CO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_C_XOR;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D1;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D2;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D3;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D4;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_DO5;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_DO6;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D_CY;
  wire [0:0] CLBLM_R_X3Y141_SLICE_X3Y141_D_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AMUX;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_AX;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_A_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_BO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_BO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_B_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_CLK;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_CO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_CO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_C_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_DO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_DO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X6Y126_D_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_AO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_AO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_A_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_BO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_BO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_B_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_CO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_C_XOR;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D1;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D2;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D3;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D4;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_DO5;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_DO6;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D_CY;
  wire [0:0] CLBLM_R_X5Y126_SLICE_X7Y126_D_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_AO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_AO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_A_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_BO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_BO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_B_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CLK;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_C_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_DMUX;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_DO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_DO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X6Y127_D_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_AO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_AO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_A_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_BO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_BO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_B_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_CO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_CO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_C_XOR;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D1;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D2;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D3;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D4;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_DO5;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_DO6;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D_CY;
  wire [0:0] CLBLM_R_X5Y127_SLICE_X7Y127_D_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_AO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_AO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_A_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_BO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_BO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_B_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_CLK;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_CMUX;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_CO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_CO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_C_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_DO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_DO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X6Y128_D_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_AO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_AO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_A_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_BO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_BO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_B_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_CO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_CO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_C_XOR;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D1;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D2;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D3;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D4;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_DO5;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_DO6;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D_CY;
  wire [0:0] CLBLM_R_X5Y128_SLICE_X7Y128_D_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_AO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_AO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_AQ;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_A_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_BO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_BO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_B_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_CLK;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_CO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_CO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_C_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_DO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_DO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X6Y129_D_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_AO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_AO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_A_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B5Q;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_BMUX;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_BO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_BO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_BQ;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_B_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_CLK;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_CO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_CO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_C_XOR;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D1;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D2;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D3;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D4;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_DO5;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_DO6;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D_CY;
  wire [0:0] CLBLM_R_X5Y129_SLICE_X7Y129_D_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_AO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_AO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_A_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B5Q;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_BMUX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_BO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_BO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_B_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_CLK;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_CO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_CO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_C_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_DO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_DO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X6Y130_D_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_AO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_AO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_AQ;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_A_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_BO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_BO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_BQ;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_B_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_CLK;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_CO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_CO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_CQ;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_C_XOR;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D1;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D2;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D3;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D4;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D5Q;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_DMUX;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_DO5;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_DO6;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_DQ;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D_CY;
  wire [0:0] CLBLM_R_X5Y130_SLICE_X7Y130_D_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_AO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_AO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_AQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_A_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_BO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_BO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_BQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_B_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_CLK;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_CMUX;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_CO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_CO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_C_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_DO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_DO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X6Y131_D_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_AO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_AO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_AQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_A_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_BO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_BO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_B_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_CLK;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_CO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_CO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_CQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_C_XOR;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D1;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D2;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D3;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D4;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D5Q;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_DMUX;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_DO5;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_DO6;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_DQ;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D_CY;
  wire [0:0] CLBLM_R_X5Y131_SLICE_X7Y131_D_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_AO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_AO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_AQ;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_A_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_BO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_BO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_B_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_CLK;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_CO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_CO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_C_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_DO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_DO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X6Y132_D_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_AO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_AO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_AQ;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_A_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_BO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_BO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_BQ;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_B_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C5Q;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_CLK;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_CMUX;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_CO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_CO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_CQ;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_C_XOR;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D1;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D2;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D3;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D4;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_DO5;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D_CY;
  wire [0:0] CLBLM_R_X5Y132_SLICE_X7Y132_D_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A5Q;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_AMUX;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_AO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_AO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_AQ;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_A_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B5Q;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_BMUX;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_BO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_BO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_BQ;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_B_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_CLK;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_CMUX;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_CO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_CO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_C_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_DO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_DO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X6Y133_D_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A5Q;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_AMUX;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_AO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_AO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_AQ;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_A_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B5Q;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_BMUX;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_BO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_BO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_B_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C5Q;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_CLK;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_CMUX;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_CO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_CO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_CQ;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_C_XOR;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D1;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D2;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D3;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D4;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_DO5;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_DO6;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_DQ;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D_CY;
  wire [0:0] CLBLM_R_X5Y133_SLICE_X7Y133_D_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A5Q;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_AMUX;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_AO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_AO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_AQ;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_A_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B5Q;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_BMUX;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_BO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_BO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_BQ;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_B_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C5Q;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_CLK;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_CMUX;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_CO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_CO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_CQ;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_CX;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_C_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_DO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_DO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_DQ;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X6Y134_D_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A5Q;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_AMUX;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_AO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_AO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_AQ;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_A_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_BO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_BO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_BQ;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_B_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_CLK;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_CO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_CO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_CQ;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_C_XOR;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D1;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D2;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D3;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D4;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D5Q;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_DMUX;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_DO5;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_DO6;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_DQ;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D_CY;
  wire [0:0] CLBLM_R_X5Y134_SLICE_X7Y134_D_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A5Q;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_AMUX;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_AO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_AO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_AQ;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_A_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B5Q;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_BMUX;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_BO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_BO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_BQ;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_B_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_CLK;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_CMUX;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_CO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_CO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_C_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_DO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_DO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X6Y135_D_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_AO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_AO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_AQ;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_A_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B5Q;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_BMUX;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_BO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_BO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_BQ;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_B_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_CLK;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_CO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_CO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_CQ;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_C_XOR;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D1;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D2;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D3;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D4;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D5Q;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_DMUX;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_DO5;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_DO6;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_DQ;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D_CY;
  wire [0:0] CLBLM_R_X5Y135_SLICE_X7Y135_D_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_AO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_AO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_AQ;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_A_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_BMUX;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_BO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_BO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_BQ;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_B_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_CLK;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_CO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_CO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_CQ;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_C_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_DO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_DO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_DQ;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X6Y136_D_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_AO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_AO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_AQ;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_A_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_BO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_BO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_BQ;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_B_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C5Q;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_CLK;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_CMUX;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_CO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_CO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_CQ;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_C_XOR;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D1;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D2;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D3;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D4;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D5Q;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_DMUX;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_DO5;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_DO6;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_DQ;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D_CY;
  wire [0:0] CLBLM_R_X5Y136_SLICE_X7Y136_D_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_AO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_AO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_AQ;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_A_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_BO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_BO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_BQ;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_B_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_CLK;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_CO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_CO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_CQ;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_C_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_DMUX;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_DO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_DO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X6Y137_D_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A5Q;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_AMUX;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_AO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_AO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_AQ;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_A_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B5Q;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_BMUX;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_BO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_BO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_BQ;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_B_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_CLK;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_CO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_CO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_C_XOR;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D1;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D2;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D3;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D4;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_DO5;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D_CY;
  wire [0:0] CLBLM_R_X5Y137_SLICE_X7Y137_D_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_AO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_AO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_A_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B5Q;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_BMUX;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_BO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_BQ;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_B_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_CLK;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_CO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_CO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_CQ;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_C_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_DMUX;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_DO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_DO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X6Y138_D_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_AO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_AO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_AQ;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_A_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_BMUX;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_BO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_BO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_B_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_CLK;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_CO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_CO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_C_XOR;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D1;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D2;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D3;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D4;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_DO5;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_DO6;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D_CY;
  wire [0:0] CLBLM_R_X5Y138_SLICE_X7Y138_D_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_AO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_AO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_AQ;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_A_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_BO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_B_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C5Q;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_CLK;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_CMUX;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_CO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_CO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_CQ;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_C_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_DO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_DO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X6Y139_D_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A5Q;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_AMUX;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_AO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_AO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_AQ;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_A_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B5Q;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_BMUX;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_BO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_BO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_BQ;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_B_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_CLK;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_CO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_CO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_CQ;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_C_XOR;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D1;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D2;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D3;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D4;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_DO5;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_DO6;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D_CY;
  wire [0:0] CLBLM_R_X5Y139_SLICE_X7Y139_D_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A5Q;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_AMUX;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_AO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_AO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_AQ;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_AX;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_A_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_BMUX;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_BO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_BO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_B_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_CLK;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_CO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_CO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_CQ;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_C_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_DO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_DO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X6Y140_D_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A5Q;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_AMUX;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_AO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_AO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_AQ;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_A_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B5Q;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_BMUX;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_BO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_BO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_BQ;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_B_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_CLK;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_CO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_CO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_CQ;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_C_XOR;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D1;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D2;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D3;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D4;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_DO5;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_DO6;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D_CY;
  wire [0:0] CLBLM_R_X5Y140_SLICE_X7Y140_D_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_AO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_AO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_A_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_BO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_BO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_BQ;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_B_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_CLK;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_CO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_CO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_CQ;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_C_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_DO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_DO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_DQ;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X6Y141_D_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_AMUX;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_AO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_AO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_A_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_BO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_BO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_B_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_CO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_CO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_C_XOR;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D1;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D2;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D3;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D4;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_DO5;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_DO6;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D_CY;
  wire [0:0] CLBLM_R_X5Y141_SLICE_X7Y141_D_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_AO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_AO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_AQ;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_A_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B5Q;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_BMUX;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_BO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_BO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_BQ;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_B_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_CLK;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_CO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_CO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_CQ;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_C_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_DO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_DO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X6Y142_D_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_AO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_AO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_A_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_BMUX;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_BO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_BO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_B_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_CLK;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_CO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_CO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_C_XOR;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D1;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D2;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D3;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D4;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_DO5;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_DO6;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D_CY;
  wire [0:0] CLBLM_R_X5Y142_SLICE_X7Y142_D_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_AO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_AO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_A_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_BO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_BO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_B_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_CO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_CO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_C_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_DO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_DO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X6Y143_D_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_AO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_AO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_AQ;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_A_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_BO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_BO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_B_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_CLK;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_CO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_CO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_C_XOR;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D1;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D2;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D3;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D4;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_DO5;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_DO6;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D_CY;
  wire [0:0] CLBLM_R_X5Y143_SLICE_X7Y143_D_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_AO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_AO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_AX;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_A_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_BO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_BO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_B_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_CE;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_CLK;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_CO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_CO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_C_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_DO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_DO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X8Y129_D_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_AO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_AO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_A_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_BO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_BO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_B_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_CO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_CO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_C_XOR;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D1;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D2;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D3;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D4;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_DO5;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_DO6;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D_CY;
  wire [0:0] CLBLM_R_X7Y129_SLICE_X9Y129_D_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_AO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_AO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_A_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_BO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_BO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_B_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_CLK;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_CMUX;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_CO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_C_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_DMUX;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_DO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_DO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X8Y130_D_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_AO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_AO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_AQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_A_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_BO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_BO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_B_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_CLK;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_CO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_CO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_C_XOR;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D1;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D2;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D3;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D4;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_DO5;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_DO6;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D_CY;
  wire [0:0] CLBLM_R_X7Y130_SLICE_X9Y130_D_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A5Q;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_AMUX;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_AO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_AO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_AX;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_A_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_BMUX;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_BO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_BO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_B_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C5Q;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CLK;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CMUX;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_CQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_C_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_DO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_DO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_DQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X8Y131_D_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_AO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_AO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_A_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_BO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_BO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_BQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_B_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_CLK;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_CO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_CO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_CQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_C_XOR;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D1;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D2;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D3;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D4;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D5Q;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_DMUX;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_DO5;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_DO6;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_DQ;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D_CY;
  wire [0:0] CLBLM_R_X7Y131_SLICE_X9Y131_D_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_AO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_AO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_A_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_BO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_BO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_BQ;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_B_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_CLK;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_CO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_CO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_CQ;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_C_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D5Q;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_DMUX;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_DO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_DO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_DQ;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X8Y132_D_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A5Q;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_AMUX;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_AO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_AQ;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_A_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_BO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_BO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_BQ;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_B_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_CLK;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_CO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_CO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_CQ;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_C_XOR;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D1;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D2;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D3;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D4;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D5Q;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_DMUX;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_DO5;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_DO6;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_DQ;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D_CY;
  wire [0:0] CLBLM_R_X7Y132_SLICE_X9Y132_D_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A5Q;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_AMUX;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_AO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_AO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_AQ;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_A_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_BO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_BO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_BQ;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_B_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C5Q;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_CLK;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_CMUX;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_CO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_CO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_CQ;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_C_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D5Q;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_DMUX;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_DO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_DO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_DQ;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X8Y133_D_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A5Q;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_AMUX;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_AO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_AO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_AQ;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_A_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B5Q;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_BMUX;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_BO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_BQ;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_B_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C5Q;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_CLK;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_CMUX;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_CO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_CO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_CQ;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_C_XOR;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D1;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D2;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D3;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D4;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D5Q;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_DMUX;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_DO5;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_DO6;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_DQ;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D_CY;
  wire [0:0] CLBLM_R_X7Y133_SLICE_X9Y133_D_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A5Q;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_AMUX;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_AO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_AO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_AQ;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_A_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B5Q;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_BMUX;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_BO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_BO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_BQ;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_B_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C5Q;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_CLK;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_CMUX;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_CO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_CO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_CQ;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_C_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_DMUX;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_DO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_DO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X8Y134_D_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_AO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_AO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_AQ;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_A_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_BO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_BO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_BQ;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_B_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_CLK;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_CO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_CO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_CQ;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_C_XOR;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D1;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D2;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D3;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D4;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_DO5;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_DO6;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_DQ;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D_CY;
  wire [0:0] CLBLM_R_X7Y134_SLICE_X9Y134_D_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_AO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_AO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_AQ;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_AX;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_A_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_BO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_BO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_BQ;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_BX;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_B_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_CE;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_CLK;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_CO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_CO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_C_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_DO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_DO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X8Y135_D_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A5Q;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_AMUX;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_AO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_AO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_AQ;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_A_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B5Q;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_BMUX;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_BO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_BO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_BX;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_B_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C5Q;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_CLK;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_CMUX;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_CO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_CQ;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_C_XOR;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D1;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D2;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D3;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D4;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D5Q;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_DMUX;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_DO5;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_DO6;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_DQ;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D_CY;
  wire [0:0] CLBLM_R_X7Y135_SLICE_X9Y135_D_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A5Q;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_AMUX;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_AO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_AO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_AQ;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_A_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B5Q;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_BMUX;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_BO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_BO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_BQ;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_B_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C5Q;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_CLK;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_CMUX;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_CO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_CO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_CQ;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_C_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D5Q;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_DMUX;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_DO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_DO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_DQ;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X8Y136_D_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A5Q;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_AMUX;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_AO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_AO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_A_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_BO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_BO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_BQ;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_B_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_CLK;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_CO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_CO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_CQ;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_C_XOR;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D1;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D2;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D3;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D4;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D5Q;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_DMUX;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_DO5;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_DO6;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_DQ;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D_CY;
  wire [0:0] CLBLM_R_X7Y136_SLICE_X9Y136_D_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_AO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_AO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_AQ;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_A_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B5Q;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_BMUX;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_BO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_BO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_BQ;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_B_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C5Q;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_CLK;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_CMUX;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_CO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_CO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_CQ;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_C_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D5Q;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_DMUX;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_DO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_DO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_DQ;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X8Y137_D_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_AO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_AO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_AQ;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_A_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_BO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_BO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_BQ;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_B_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_CLK;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_CO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_CO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_CQ;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_C_XOR;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D1;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D2;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D3;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D4;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D5Q;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_DMUX;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_DO5;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_DO6;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_DQ;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D_CY;
  wire [0:0] CLBLM_R_X7Y137_SLICE_X9Y137_D_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_AO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_AO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_AQ;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_A_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B5Q;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_BMUX;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_BO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_BO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_BQ;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_B_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_CLK;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_CO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_CO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_CQ;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_C_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D5Q;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_DMUX;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_DO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_DO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_DQ;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X8Y138_D_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A5Q;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_AMUX;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_AO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_AO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_AQ;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_A_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B5Q;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_BMUX;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_BO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_BQ;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_B_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C5Q;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_CLK;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_CMUX;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_CO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_CO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_CQ;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_C_XOR;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D1;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D2;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D3;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D4;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_DO5;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_DO6;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D_CY;
  wire [0:0] CLBLM_R_X7Y138_SLICE_X9Y138_D_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_AMUX;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_AO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_AO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_AQ;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_AX;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_A_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_BO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_BO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_B_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_CE;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_CLK;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_CO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_CO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_C_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_DO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_DO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X8Y139_D_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_AO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_AO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_AQ;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_A_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_BO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_BO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_BQ;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_B_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_CLK;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_CO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_CO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_C_XOR;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D1;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D2;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D3;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D4;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_DO5;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D_CY;
  wire [0:0] CLBLM_R_X7Y139_SLICE_X9Y139_D_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_AO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_AO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_AQ;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_A_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B5Q;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_BMUX;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_BO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_BO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_BQ;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_B_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C5Q;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_CLK;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_CMUX;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_CO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_CO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_CQ;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_C_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D5Q;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_DMUX;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_DO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_DO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_DQ;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X8Y140_D_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_AO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_AO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_AQ;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_A_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_BO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_BO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_BQ;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_B_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_CLK;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_CO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_CO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_CQ;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_C_XOR;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D1;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D2;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D3;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D4;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D5Q;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_DMUX;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_DO5;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_DO6;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_DQ;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D_CY;
  wire [0:0] CLBLM_R_X7Y140_SLICE_X9Y140_D_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A5Q;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_AMUX;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_AO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_AO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_AQ;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_AX;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_A_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_BMUX;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_BO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_BO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_B_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_CLK;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_CO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_CO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_C_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_DO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X8Y141_D_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A5Q;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_AMUX;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_AO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_AO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_A_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_BO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_BO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_B_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_CLK;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_CO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_CO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_C_XOR;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D1;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D2;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D3;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D4;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_DO5;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_DO6;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D_CY;
  wire [0:0] CLBLM_R_X7Y141_SLICE_X9Y141_D_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_AO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_AO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_A_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_BO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_BO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_B_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_CO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_C_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_DO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X8Y142_D_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_AO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_AO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_AQ;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_A_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_BO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_BO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_BQ;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_B_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_CLK;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_CO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_CO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_CQ;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_C_XOR;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D1;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D2;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D3;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D4;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_DMUX;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_DO5;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D_CY;
  wire [0:0] CLBLM_R_X7Y142_SLICE_X9Y142_D_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A5Q;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_AMUX;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_AO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_AO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_AX;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_A_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_BMUX;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_BO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_BO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_B_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_CLK;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_CO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_CO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_C_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_DO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_DO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X8Y143_D_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_AO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_AO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_A_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_BMUX;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_BO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_BO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_B_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_CLK;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_CO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_CO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_C_XOR;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D1;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D2;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D3;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D4;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_DO5;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_DO6;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D_CY;
  wire [0:0] CLBLM_R_X7Y143_SLICE_X9Y143_D_XOR;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_O;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_O;
  wire [0:0] LIOB33_SING_X0Y150_IOB_X0Y150_O;
  wire [0:0] LIOB33_SING_X0Y199_IOB_X0Y199_O;
  wire [0:0] LIOB33_SING_X0Y50_IOB_X0Y50_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_O;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y151_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y152_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y153_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y154_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y155_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y156_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y157_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y158_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y159_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y160_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y161_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y162_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y163_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y164_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y165_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y166_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y167_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y168_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y169_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y170_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y171_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y172_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y173_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y174_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y175_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y176_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y177_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y178_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y179_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y180_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y181_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y182_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y183_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y184_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y185_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y186_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y187_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y188_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y189_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y190_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y191_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y192_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y193_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y194_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y195_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y196_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y197_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y198_O;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y51_I;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y52_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y53_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y54_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y55_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y56_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y57_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y58_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y59_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y60_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y61_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y62_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y63_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y64_O;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y65_O;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y66_O;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y78_I;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_D;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_TQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_TQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_TQ;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_O;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_O;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y65_D1;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y65_OQ;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y65_T1;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y65_TQ;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y66_D1;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y66_OQ;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y66_T1;
  wire [0:0] LIOI3_X0Y65_OLOGIC_X0Y66_TQ;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_O;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_I;
  wire [0:0] RIOB33_SING_X105Y149_IOB_X1Y149_I;
  wire [0:0] RIOB33_SING_X105Y150_IOB_X1Y150_O;
  wire [0:0] RIOB33_SING_X105Y199_IOB_X1Y199_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y114_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y115_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y116_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y117_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y118_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y119_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y120_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y121_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y122_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y123_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y124_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y125_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y126_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y127_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y128_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y129_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y130_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y131_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y132_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y133_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y134_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y135_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y136_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y137_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y138_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y139_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y140_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y141_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y142_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y143_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y144_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y145_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y146_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y147_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y148_I;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y151_O;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y152_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y153_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y154_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y155_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y156_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y157_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y158_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y159_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y160_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y161_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y162_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y163_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y164_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y165_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y166_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y167_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y168_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y169_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y170_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y171_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y172_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y173_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y174_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y175_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y176_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y177_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y178_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y179_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y180_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y181_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y182_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y183_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y184_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y185_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y186_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y187_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y188_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y189_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y190_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y191_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y192_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y193_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y194_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y195_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y196_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y197_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y198_O;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_D;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_O;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_D;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_O;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_O;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_TQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_TQ;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X0Y75_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X0Y75_DO5),
.O6(CLBLL_L_X2Y75_SLICE_X0Y75_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X0Y75_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X0Y75_CO5),
.O6(CLBLL_L_X2Y75_SLICE_X0Y75_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X0Y75_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X0Y75_BO5),
.O6(CLBLL_L_X2Y75_SLICE_X0Y75_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0f)
  ) CLBLL_L_X2Y75_SLICE_X0Y75_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y55_IOB_X0Y56_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X0Y75_AO5),
.O6(CLBLL_L_X2Y75_SLICE_X0Y75_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X1Y75_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X1Y75_DO5),
.O6(CLBLL_L_X2Y75_SLICE_X1Y75_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X1Y75_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X1Y75_CO5),
.O6(CLBLL_L_X2Y75_SLICE_X1Y75_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X1Y75_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X1Y75_BO5),
.O6(CLBLL_L_X2Y75_SLICE_X1Y75_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y75_SLICE_X1Y75_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y75_SLICE_X1Y75_AO5),
.O6(CLBLL_L_X2Y75_SLICE_X1Y75_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y133_SLICE_X0Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X0Y133_DO5),
.O6(CLBLL_L_X2Y133_SLICE_X0Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y133_SLICE_X0Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X0Y133_CO5),
.O6(CLBLL_L_X2Y133_SLICE_X0Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y133_SLICE_X0Y133_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X0Y133_BO5),
.O6(CLBLL_L_X2Y133_SLICE_X0Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y133_SLICE_X0Y133_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X0Y133_AO5),
.O6(CLBLL_L_X2Y133_SLICE_X0Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y133_SLICE_X1Y133_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X1Y133_DO5),
.O6(CLBLL_L_X2Y133_SLICE_X1Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y133_SLICE_X1Y133_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X1Y133_CO5),
.O6(CLBLL_L_X2Y133_SLICE_X1Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800000088000000)
  ) CLBLL_L_X2Y133_SLICE_X1Y133_BLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(CLBLM_R_X7Y134_SLICE_X8Y134_CQ),
.I2(1'b1),
.I3(CLBLM_R_X3Y141_SLICE_X2Y141_CO6),
.I4(CLBLL_L_X4Y138_SLICE_X4Y138_BQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y133_SLICE_X1Y133_BO5),
.O6(CLBLL_L_X2Y133_SLICE_X1Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000008000)
  ) CLBLL_L_X2Y133_SLICE_X1Y133_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLM_R_X3Y133_SLICE_X2Y133_AQ),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLL_L_X2Y133_SLICE_X1Y133_AO5),
.O6(CLBLL_L_X2Y133_SLICE_X1Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y134_SLICE_X0Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y134_SLICE_X0Y134_DO5),
.O6(CLBLL_L_X2Y134_SLICE_X0Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y134_SLICE_X0Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y134_SLICE_X0Y134_CO5),
.O6(CLBLL_L_X2Y134_SLICE_X0Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y134_SLICE_X0Y134_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y134_SLICE_X0Y134_BO5),
.O6(CLBLL_L_X2Y134_SLICE_X0Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y134_SLICE_X0Y134_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y134_SLICE_X0Y134_AO5),
.O6(CLBLL_L_X2Y134_SLICE_X0Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y134_SLICE_X1Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y134_SLICE_X1Y134_DO5),
.O6(CLBLL_L_X2Y134_SLICE_X1Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y134_SLICE_X1Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y134_SLICE_X1Y134_CO5),
.O6(CLBLL_L_X2Y134_SLICE_X1Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y134_SLICE_X1Y134_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y134_SLICE_X1Y134_BO5),
.O6(CLBLL_L_X2Y134_SLICE_X1Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff20200000)
  ) CLBLL_L_X2Y134_SLICE_X1Y134_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(CLBLL_L_X4Y138_SLICE_X4Y138_BQ),
.I3(CLBLM_R_X3Y135_SLICE_X2Y135_AQ),
.I4(CLBLM_R_X3Y141_SLICE_X2Y141_CO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y134_SLICE_X1Y134_AO5),
.O6(CLBLL_L_X2Y134_SLICE_X1Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y138_SLICE_X0Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X0Y138_DO5),
.O6(CLBLL_L_X2Y138_SLICE_X0Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y138_SLICE_X0Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X0Y138_CO5),
.O6(CLBLL_L_X2Y138_SLICE_X0Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y138_SLICE_X0Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X0Y138_BO5),
.O6(CLBLL_L_X2Y138_SLICE_X0Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y138_SLICE_X0Y138_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X0Y138_AO5),
.O6(CLBLL_L_X2Y138_SLICE_X0Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y138_SLICE_X1Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X1Y138_DO5),
.O6(CLBLL_L_X2Y138_SLICE_X1Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y138_SLICE_X1Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X1Y138_CO5),
.O6(CLBLL_L_X2Y138_SLICE_X1Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000400000000)
  ) CLBLL_L_X2Y138_SLICE_X1Y138_BLUT (
.I0(CLBLM_R_X3Y137_SLICE_X3Y137_CQ),
.I1(CLBLM_R_X3Y139_SLICE_X3Y139_BQ),
.I2(CLBLM_R_X5Y138_SLICE_X6Y138_B5Q),
.I3(LIOB33_X0Y61_IOB_X0Y61_I),
.I4(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLL_L_X2Y138_SLICE_X1Y138_BO5),
.O6(CLBLL_L_X2Y138_SLICE_X1Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffafafffffffa)
  ) CLBLL_L_X2Y138_SLICE_X1Y138_ALUT (
.I0(CLBLM_R_X3Y137_SLICE_X3Y137_CQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y138_SLICE_X6Y138_B5Q),
.I3(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.I4(LIOB33_X0Y61_IOB_X0Y61_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y138_SLICE_X1Y138_AO5),
.O6(CLBLL_L_X2Y138_SLICE_X1Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y129_SLICE_X4Y129_AO6),
.Q(CLBLL_L_X4Y129_SLICE_X4Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y129_SLICE_X4Y129_DO5),
.O6(CLBLL_L_X4Y129_SLICE_X4Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y129_SLICE_X4Y129_CO5),
.O6(CLBLL_L_X4Y129_SLICE_X4Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y129_SLICE_X4Y129_BO5),
.O6(CLBLL_L_X4Y129_SLICE_X4Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeeeeee22222222)
  ) CLBLL_L_X4Y129_SLICE_X4Y129_ALUT (
.I0(CLBLM_R_X3Y135_SLICE_X3Y135_CQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y63_IOB_X0Y63_I),
.O5(CLBLL_L_X4Y129_SLICE_X4Y129_AO5),
.O6(CLBLL_L_X4Y129_SLICE_X4Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y129_SLICE_X5Y129_DO5),
.O6(CLBLL_L_X4Y129_SLICE_X5Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y129_SLICE_X5Y129_CO5),
.O6(CLBLL_L_X4Y129_SLICE_X5Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y129_SLICE_X5Y129_BO5),
.O6(CLBLL_L_X4Y129_SLICE_X5Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y129_SLICE_X5Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y129_SLICE_X5Y129_AO5),
.O6(CLBLL_L_X4Y129_SLICE_X5Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y130_SLICE_X4Y130_BO5),
.Q(CLBLL_L_X4Y130_SLICE_X4Y130_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y130_SLICE_X4Y130_DO5),
.Q(CLBLL_L_X4Y130_SLICE_X4Y130_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y130_SLICE_X4Y130_AO6),
.Q(CLBLL_L_X4Y130_SLICE_X4Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y130_SLICE_X4Y130_BO6),
.Q(CLBLL_L_X4Y130_SLICE_X4Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y130_SLICE_X4Y130_DO6),
.Q(CLBLL_L_X4Y130_SLICE_X4Y130_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f0f0ccccaaaa)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_DLUT (
.I0(RIOB33_X105Y121_IOB_X1Y122_I),
.I1(CLBLL_L_X4Y130_SLICE_X5Y130_A5Q),
.I2(CLBLM_R_X5Y133_SLICE_X7Y133_CQ),
.I3(CLBLM_R_X5Y133_SLICE_X7Y133_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y130_SLICE_X4Y130_DO5),
.O6(CLBLL_L_X4Y130_SLICE_X4Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00cccc08080808)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_CLUT (
.I0(CLBLM_R_X5Y129_SLICE_X6Y129_AQ),
.I1(CLBLL_L_X4Y130_SLICE_X4Y130_AQ),
.I2(CLBLM_R_X5Y130_SLICE_X6Y130_CO6),
.I3(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y130_SLICE_X4Y130_CO5),
.O6(CLBLL_L_X4Y130_SLICE_X4Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee2222e2e2e2e2)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_BLUT (
.I0(CLBLM_R_X5Y133_SLICE_X7Y133_BQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y138_SLICE_X4Y138_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y130_SLICE_X4Y130_BO5),
.O6(CLBLL_L_X4Y130_SLICE_X4Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff21ff3000210030)
  ) CLBLL_L_X4Y130_SLICE_X4Y130_ALUT (
.I0(CLBLM_R_X5Y130_SLICE_X6Y130_CO6),
.I1(CLBLM_R_X5Y130_SLICE_X6Y130_B5Q),
.I2(CLBLL_L_X4Y130_SLICE_X4Y130_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y129_SLICE_X6Y129_AQ),
.I5(CLBLM_R_X7Y131_SLICE_X8Y131_C5Q),
.O5(CLBLL_L_X4Y130_SLICE_X4Y130_AO5),
.O6(CLBLL_L_X4Y130_SLICE_X4Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y130_SLICE_X4Y130_CO6),
.Q(CLBLL_L_X4Y130_SLICE_X5Y130_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y130_SLICE_X5Y130_BO5),
.Q(CLBLL_L_X4Y130_SLICE_X5Y130_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y130_SLICE_X5Y130_AO6),
.Q(CLBLL_L_X4Y130_SLICE_X5Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y130_SLICE_X5Y130_BO6),
.Q(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f7fffffaafaaafa)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_DLUT (
.I0(CLBLL_L_X4Y130_SLICE_X4Y130_AQ),
.I1(CLBLL_L_X4Y130_SLICE_X5Y130_AQ),
.I2(CLBLM_R_X5Y129_SLICE_X6Y129_AQ),
.I3(CLBLM_R_X5Y130_SLICE_X6Y130_CO6),
.I4(CLBLL_L_X4Y131_SLICE_X4Y131_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y130_SLICE_X5Y130_DO5),
.O6(CLBLL_L_X4Y130_SLICE_X5Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffff7fff7fff)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_CLUT (
.I0(CLBLM_R_X5Y130_SLICE_X7Y130_BQ),
.I1(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I2(CLBLL_L_X4Y134_SLICE_X4Y134_CQ),
.I3(CLBLM_R_X7Y131_SLICE_X8Y131_A5Q),
.I4(CLBLM_R_X3Y131_SLICE_X3Y131_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y130_SLICE_X5Y130_CO5),
.O6(CLBLL_L_X4Y130_SLICE_X5Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa00aaccaaccaa)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_BLUT (
.I0(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y141_SLICE_X4Y141_DQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y130_SLICE_X5Y130_BO5),
.O6(CLBLL_L_X4Y130_SLICE_X5Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfff5ccccff5f)
  ) CLBLL_L_X4Y130_SLICE_X5Y130_ALUT (
.I0(CLBLL_L_X4Y130_SLICE_X5Y130_DO6),
.I1(CLBLM_R_X3Y137_SLICE_X3Y137_D5Q),
.I2(CLBLL_L_X4Y130_SLICE_X5Y130_AQ),
.I3(CLBLM_R_X5Y130_SLICE_X6Y130_B5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X4Y130_SLICE_X5Y130_CO6),
.O5(CLBLL_L_X4Y130_SLICE_X5Y130_AO5),
.O6(CLBLL_L_X4Y130_SLICE_X5Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X4Y131_DO5),
.Q(CLBLL_L_X4Y131_SLICE_X4Y131_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X4Y131_AO6),
.Q(CLBLL_L_X4Y131_SLICE_X4Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X4Y131_BO6),
.Q(CLBLL_L_X4Y131_SLICE_X4Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X4Y131_CO6),
.Q(CLBLL_L_X4Y131_SLICE_X4Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X4Y131_DO6),
.Q(CLBLL_L_X4Y131_SLICE_X4Y131_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55aa00e4e4e4e4)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y132_SLICE_X5Y132_A5Q),
.I2(CLBLL_L_X4Y131_SLICE_X4Y131_DQ),
.I3(CLBLM_R_X3Y132_SLICE_X3Y132_D5Q),
.I4(CLBLM_R_X3Y135_SLICE_X3Y135_DQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X4Y131_DO5),
.O6(CLBLL_L_X4Y131_SLICE_X4Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaeaffee50405544)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y131_SLICE_X4Y131_CQ),
.I2(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I3(CLBLM_R_X3Y131_SLICE_X3Y131_B5Q),
.I4(CLBLL_L_X4Y135_SLICE_X5Y135_CQ),
.I5(CLBLM_R_X5Y130_SLICE_X7Y130_D5Q),
.O5(CLBLL_L_X4Y131_SLICE_X4Y131_CO5),
.O6(CLBLL_L_X4Y131_SLICE_X4Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0003030c0c)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y131_SLICE_X4Y131_BQ),
.I2(CLBLM_R_X5Y130_SLICE_X6Y130_B5Q),
.I3(CLBLL_L_X4Y132_SLICE_X4Y132_BQ),
.I4(CLBLL_L_X4Y130_SLICE_X4Y130_CO5),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y131_SLICE_X4Y131_BO5),
.O6(CLBLL_L_X4Y131_SLICE_X4Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbb88888bbb8bbb8)
  ) CLBLL_L_X4Y131_SLICE_X4Y131_ALUT (
.I0(CLBLM_R_X5Y141_SLICE_X6Y141_CQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y131_SLICE_X4Y131_AQ),
.I3(CLBLM_R_X3Y132_SLICE_X3Y132_D5Q),
.I4(CLBLM_R_X5Y133_SLICE_X7Y133_AQ),
.I5(CLBLL_L_X4Y135_SLICE_X4Y135_D5Q),
.O5(CLBLL_L_X4Y131_SLICE_X4Y131_AO5),
.O6(CLBLL_L_X4Y131_SLICE_X4Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X5Y131_BO5),
.Q(CLBLL_L_X4Y131_SLICE_X5Y131_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X5Y131_AO6),
.Q(CLBLL_L_X4Y131_SLICE_X5Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y131_SLICE_X5Y131_BO6),
.Q(CLBLL_L_X4Y131_SLICE_X5Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5ff55ff5affaaffa)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_DLUT (
.I0(CLBLM_L_X8Y134_SLICE_X10Y134_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I3(CLBLM_L_X8Y139_SLICE_X11Y139_C5Q),
.I4(1'b1),
.I5(CLBLL_L_X4Y131_SLICE_X4Y131_BQ),
.O5(CLBLL_L_X4Y131_SLICE_X5Y131_DO5),
.O6(CLBLL_L_X4Y131_SLICE_X5Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7d7d7d7dbebebebe)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_CLUT (
.I0(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.I1(CLBLM_R_X3Y137_SLICE_X3Y137_C5Q),
.I2(CLBLL_L_X4Y130_SLICE_X4Y130_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X3Y131_SLICE_X3Y131_AQ),
.O5(CLBLL_L_X4Y131_SLICE_X5Y131_CO5),
.O6(CLBLL_L_X4Y131_SLICE_X5Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc3300fc30fc30)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X11Y135_SLICE_X14Y135_AO6),
.I3(CLBLL_L_X4Y131_SLICE_X4Y131_BQ),
.I4(CLBLM_R_X5Y138_SLICE_X7Y138_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y131_SLICE_X5Y131_BO5),
.O6(CLBLL_L_X4Y131_SLICE_X5Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf5cca0ccf0ccf0)
  ) CLBLL_L_X4Y131_SLICE_X5Y131_ALUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_C5Q),
.I1(CLBLL_L_X4Y133_SLICE_X5Y133_D5Q),
.I2(CLBLL_L_X4Y131_SLICE_X5Y131_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y131_SLICE_X5Y131_BQ),
.I5(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.O5(CLBLL_L_X4Y131_SLICE_X5Y131_AO5),
.O6(CLBLL_L_X4Y131_SLICE_X5Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y132_SLICE_X4Y132_AO6),
.Q(CLBLL_L_X4Y132_SLICE_X4Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y132_SLICE_X4Y132_BO6),
.Q(CLBLL_L_X4Y132_SLICE_X4Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y132_SLICE_X4Y132_CO6),
.Q(CLBLL_L_X4Y132_SLICE_X4Y132_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y132_SLICE_X4Y132_DO6),
.Q(CLBLL_L_X4Y132_SLICE_X4Y132_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff3cff00003c0000)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y132_SLICE_X11Y132_CO6),
.I2(CLBLL_L_X4Y132_SLICE_X4Y132_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.I5(CLBLM_R_X5Y133_SLICE_X6Y133_BQ),
.O5(CLBLL_L_X4Y132_SLICE_X4Y132_DO5),
.O6(CLBLL_L_X4Y132_SLICE_X4Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff340034)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_CLUT (
.I0(CLBLL_L_X4Y132_SLICE_X4Y132_BQ),
.I1(CLBLL_L_X4Y132_SLICE_X4Y132_CQ),
.I2(CLBLL_L_X4Y132_SLICE_X4Y132_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y132_SLICE_X3Y132_CQ),
.I5(CLBLL_L_X4Y133_SLICE_X4Y133_AQ),
.O5(CLBLL_L_X4Y132_SLICE_X4Y132_CO5),
.O6(CLBLL_L_X4Y132_SLICE_X4Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff640064)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_BLUT (
.I0(CLBLL_L_X4Y132_SLICE_X4Y132_CQ),
.I1(CLBLL_L_X4Y132_SLICE_X4Y132_BQ),
.I2(CLBLL_L_X4Y132_SLICE_X4Y132_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y133_SLICE_X4Y133_C5Q),
.I5(CLBLL_L_X4Y133_SLICE_X4Y133_AQ),
.O5(CLBLL_L_X4Y132_SLICE_X4Y132_BO5),
.O6(CLBLL_L_X4Y132_SLICE_X4Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccffccafcc0f)
  ) CLBLL_L_X4Y132_SLICE_X4Y132_ALUT (
.I0(CLBLL_L_X4Y132_SLICE_X4Y132_CQ),
.I1(CLBLL_L_X4Y136_SLICE_X5Y136_D5Q),
.I2(CLBLL_L_X4Y132_SLICE_X4Y132_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y132_SLICE_X4Y132_BQ),
.I5(CLBLL_L_X4Y133_SLICE_X4Y133_AQ),
.O5(CLBLL_L_X4Y132_SLICE_X4Y132_AO5),
.O6(CLBLL_L_X4Y132_SLICE_X4Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y132_SLICE_X5Y132_AO5),
.Q(CLBLL_L_X4Y132_SLICE_X5Y132_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y132_SLICE_X5Y132_CO5),
.Q(CLBLL_L_X4Y132_SLICE_X5Y132_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y132_SLICE_X5Y132_DO5),
.Q(CLBLL_L_X4Y132_SLICE_X5Y132_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y132_SLICE_X5Y132_AO6),
.Q(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y132_SLICE_X5Y132_BO6),
.Q(CLBLL_L_X4Y132_SLICE_X5Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y132_SLICE_X5Y132_CO6),
.Q(CLBLL_L_X4Y132_SLICE_X5Y132_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y132_SLICE_X5Y132_DO6),
.Q(CLBLL_L_X4Y132_SLICE_X5Y132_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d8fafa5050)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y133_SLICE_X4Y133_AQ),
.I2(CLBLM_L_X10Y140_SLICE_X13Y140_B5Q),
.I3(1'b1),
.I4(CLBLM_R_X5Y128_SLICE_X6Y128_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y132_SLICE_X5Y132_DO5),
.O6(CLBLL_L_X4Y132_SLICE_X5Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1b1e4e4fa50fa50)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_DO6),
.I2(CLBLM_R_X7Y140_SLICE_X9Y140_BQ),
.I3(CLBLM_R_X5Y134_SLICE_X7Y134_DQ),
.I4(CLBLL_L_X4Y132_SLICE_X5Y132_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y132_SLICE_X5Y132_CO5),
.O6(CLBLL_L_X4Y132_SLICE_X5Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ccccff005f5f)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_BLUT (
.I0(CLBLL_L_X4Y136_SLICE_X5Y136_CQ),
.I1(CLBLL_L_X4Y132_SLICE_X5Y132_BQ),
.I2(CLBLM_R_X5Y141_SLICE_X6Y141_CQ),
.I3(CLBLL_L_X4Y131_SLICE_X5Y131_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y134_SLICE_X7Y134_BQ),
.O5(CLBLL_L_X4Y132_SLICE_X5Y132_BO5),
.O6(CLBLL_L_X4Y132_SLICE_X5Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ccffaaccaacc)
  ) CLBLL_L_X4Y132_SLICE_X5Y132_ALUT (
.I0(CLBLL_L_X4Y136_SLICE_X5Y136_CQ),
.I1(CLBLL_L_X4Y130_SLICE_X4Y130_DQ),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y140_SLICE_X13Y140_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y132_SLICE_X5Y132_AO5),
.O6(CLBLL_L_X4Y132_SLICE_X5Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X4Y133_AO5),
.Q(CLBLL_L_X4Y133_SLICE_X4Y133_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X4Y133_CO5),
.Q(CLBLL_L_X4Y133_SLICE_X4Y133_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X4Y133_DO5),
.Q(CLBLL_L_X4Y133_SLICE_X4Y133_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X4Y133_AO6),
.Q(CLBLL_L_X4Y133_SLICE_X4Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X4Y133_BO6),
.Q(CLBLL_L_X4Y133_SLICE_X4Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X4Y133_CO6),
.Q(CLBLL_L_X4Y133_SLICE_X4Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X4Y133_DO6),
.Q(CLBLL_L_X4Y133_SLICE_X4Y133_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaccf0fff000)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_DLUT (
.I0(CLBLM_R_X5Y132_SLICE_X7Y132_AQ),
.I1(CLBLM_R_X5Y137_SLICE_X7Y137_BQ),
.I2(CLBLL_L_X4Y133_SLICE_X4Y133_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y130_SLICE_X4Y130_DQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y133_SLICE_X4Y133_DO5),
.O6(CLBLL_L_X4Y133_SLICE_X4Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55aa008d8dd8d8)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y132_SLICE_X5Y132_D5Q),
.I2(CLBLM_R_X3Y137_SLICE_X3Y137_DQ),
.I3(CLBLL_L_X4Y132_SLICE_X4Y132_DQ),
.I4(CLBLM_R_X7Y138_SLICE_X9Y138_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y133_SLICE_X4Y133_CO5),
.O6(CLBLL_L_X4Y133_SLICE_X4Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f066cc00ff00ff)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_BLUT (
.I0(CLBLM_R_X5Y134_SLICE_X6Y134_C5Q),
.I1(CLBLL_L_X4Y133_SLICE_X4Y133_BQ),
.I2(CLBLM_R_X5Y135_SLICE_X7Y135_B5Q),
.I3(LIOB33_X0Y59_IOB_X0Y60_I),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y133_SLICE_X4Y133_BO5),
.O6(CLBLL_L_X4Y133_SLICE_X4Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff005555f0f0cccc)
  ) CLBLL_L_X4Y133_SLICE_X4Y133_ALUT (
.I0(CLBLM_R_X5Y140_SLICE_X7Y140_B5Q),
.I1(CLBLM_R_X5Y133_SLICE_X6Y133_BQ),
.I2(CLBLL_L_X4Y134_SLICE_X4Y134_CQ),
.I3(CLBLM_R_X3Y133_SLICE_X2Y133_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y133_SLICE_X4Y133_AO5),
.O6(CLBLL_L_X4Y133_SLICE_X4Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X5Y133_BO5),
.Q(CLBLL_L_X4Y133_SLICE_X5Y133_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X5Y133_CO5),
.Q(CLBLL_L_X4Y133_SLICE_X5Y133_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X5Y133_DO5),
.Q(CLBLL_L_X4Y133_SLICE_X5Y133_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X5Y133_AO6),
.Q(CLBLL_L_X4Y133_SLICE_X5Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X5Y133_BO6),
.Q(CLBLL_L_X4Y133_SLICE_X5Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X5Y133_CO6),
.Q(CLBLL_L_X4Y133_SLICE_X5Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y133_SLICE_X5Y133_DO6),
.Q(CLBLL_L_X4Y133_SLICE_X5Y133_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f033ccaaaaff00)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_DLUT (
.I0(CLBLL_L_X4Y133_SLICE_X4Y133_D5Q),
.I1(CLBLM_R_X7Y140_SLICE_X8Y140_D5Q),
.I2(CLBLM_R_X5Y134_SLICE_X6Y134_C5Q),
.I3(CLBLM_R_X5Y132_SLICE_X6Y132_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y133_SLICE_X5Y133_DO5),
.O6(CLBLL_L_X4Y133_SLICE_X5Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000aaffaa00)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_CLUT (
.I0(CLBLM_L_X8Y134_SLICE_X10Y134_AQ),
.I1(1'b1),
.I2(CLBLM_R_X3Y136_SLICE_X3Y136_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y132_SLICE_X6Y132_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y133_SLICE_X5Y133_CO5),
.O6(CLBLL_L_X4Y133_SLICE_X5Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0a0fc0cfc0c)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_BLUT (
.I0(CLBLM_R_X7Y131_SLICE_X8Y131_DQ),
.I1(CLBLM_R_X5Y130_SLICE_X7Y130_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I4(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y133_SLICE_X5Y133_BO5),
.O6(CLBLL_L_X4Y133_SLICE_X5Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ea40ff55fa50)
  ) CLBLL_L_X4Y133_SLICE_X5Y133_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y140_SLICE_X13Y140_D5Q),
.I2(CLBLL_L_X4Y133_SLICE_X5Y133_AQ),
.I3(CLBLM_R_X5Y132_SLICE_X7Y132_BQ),
.I4(CLBLL_L_X4Y133_SLICE_X5Y133_C5Q),
.I5(CLBLM_R_X7Y131_SLICE_X9Y131_D5Q),
.O5(CLBLL_L_X4Y133_SLICE_X5Y133_AO5),
.O6(CLBLL_L_X4Y133_SLICE_X5Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y140_SLICE_X4Y140_AO6),
.Q(CLBLL_L_X4Y134_SLICE_X4Y134_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y134_SLICE_X4Y134_CO5),
.Q(CLBLL_L_X4Y134_SLICE_X4Y134_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y134_SLICE_X4Y134_DO5),
.Q(CLBLL_L_X4Y134_SLICE_X4Y134_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y134_SLICE_X4Y134_AO6),
.Q(CLBLL_L_X4Y134_SLICE_X4Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y134_SLICE_X4Y134_BO6),
.Q(CLBLL_L_X4Y134_SLICE_X4Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y134_SLICE_X4Y134_CO6),
.Q(CLBLL_L_X4Y134_SLICE_X4Y134_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y134_SLICE_X4Y134_DO6),
.Q(CLBLL_L_X4Y134_SLICE_X4Y134_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0caa0cfff000f0)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_DLUT (
.I0(CLBLL_L_X4Y129_SLICE_X4Y129_AQ),
.I1(CLBLM_R_X7Y136_SLICE_X8Y136_AQ),
.I2(CLBLM_R_X3Y135_SLICE_X2Y135_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y136_SLICE_X3Y136_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y134_SLICE_X4Y134_DO5),
.O6(CLBLL_L_X4Y134_SLICE_X4Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0fcc0ff0aaf0aa)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_CLUT (
.I0(CLBLM_L_X12Y133_SLICE_X16Y133_AO6),
.I1(CLBLL_L_X4Y134_SLICE_X4Y134_D5Q),
.I2(CLBLM_R_X5Y140_SLICE_X7Y140_B5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y134_SLICE_X4Y134_CO5),
.O6(CLBLL_L_X4Y134_SLICE_X4Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0aca0afafacac)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_BLUT (
.I0(CLBLM_R_X3Y135_SLICE_X3Y135_DQ),
.I1(CLBLL_L_X4Y134_SLICE_X4Y134_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_CQ),
.I4(CLBLL_L_X4Y133_SLICE_X5Y133_D5Q),
.I5(CLBLL_L_X4Y136_SLICE_X4Y136_D5Q),
.O5(CLBLL_L_X4Y134_SLICE_X4Y134_BO5),
.O6(CLBLL_L_X4Y134_SLICE_X4Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcdddc33301110)
  ) CLBLL_L_X4Y134_SLICE_X4Y134_ALUT (
.I0(CLBLM_R_X7Y131_SLICE_X9Y131_D5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y134_SLICE_X4Y134_AQ),
.I3(CLBLL_L_X4Y137_SLICE_X5Y137_D5Q),
.I4(CLBLM_L_X10Y140_SLICE_X13Y140_D5Q),
.I5(CLBLM_R_X5Y134_SLICE_X7Y134_D5Q),
.O5(CLBLL_L_X4Y134_SLICE_X4Y134_AO5),
.O6(CLBLL_L_X4Y134_SLICE_X4Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y134_SLICE_X5Y134_DO5),
.Q(CLBLL_L_X4Y134_SLICE_X5Y134_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y134_SLICE_X5Y134_AO6),
.Q(CLBLL_L_X4Y134_SLICE_X5Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y134_SLICE_X5Y134_BO6),
.Q(CLBLL_L_X4Y134_SLICE_X5Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y134_SLICE_X5Y134_CO6),
.Q(CLBLL_L_X4Y134_SLICE_X5Y134_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y134_SLICE_X5Y134_DO6),
.Q(CLBLL_L_X4Y134_SLICE_X5Y134_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0eeee4444)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y134_SLICE_X6Y134_BQ),
.I2(CLBLM_R_X5Y138_SLICE_X6Y138_B5Q),
.I3(CLBLM_R_X3Y137_SLICE_X3Y137_D5Q),
.I4(CLBLM_R_X7Y140_SLICE_X9Y140_DQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y134_SLICE_X5Y134_DO5),
.O6(CLBLL_L_X4Y134_SLICE_X5Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff002200000022)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_CLUT (
.I0(CLBLM_R_X5Y134_SLICE_X7Y134_BQ),
.I1(CLBLL_L_X4Y134_SLICE_X5Y134_CQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y139_SLICE_X5Y139_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X3Y139_SLICE_X2Y139_BQ),
.O5(CLBLL_L_X4Y134_SLICE_X5Y134_CO5),
.O6(CLBLL_L_X4Y134_SLICE_X5Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaf8c0000af8c)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_BLUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_CQ),
.I1(CLBLL_L_X4Y134_SLICE_X5Y134_BQ),
.I2(CLBLL_L_X4Y136_SLICE_X4Y136_D5Q),
.I3(CLBLM_R_X5Y135_SLICE_X6Y135_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y134_SLICE_X6Y134_BQ),
.O5(CLBLL_L_X4Y134_SLICE_X5Y134_BO5),
.O6(CLBLL_L_X4Y134_SLICE_X5Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000cccc5a5a)
  ) CLBLL_L_X4Y134_SLICE_X5Y134_ALUT (
.I0(CLBLL_L_X4Y135_SLICE_X5Y135_BQ),
.I1(CLBLM_R_X5Y135_SLICE_X6Y135_BQ),
.I2(CLBLL_L_X4Y134_SLICE_X5Y134_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLL_L_X4Y134_SLICE_X5Y134_AO5),
.O6(CLBLL_L_X4Y134_SLICE_X5Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y135_SLICE_X4Y135_CO5),
.Q(CLBLL_L_X4Y135_SLICE_X4Y135_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y135_SLICE_X4Y135_DO5),
.Q(CLBLL_L_X4Y135_SLICE_X4Y135_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y135_SLICE_X4Y135_AO6),
.Q(CLBLL_L_X4Y135_SLICE_X4Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y135_SLICE_X4Y135_BO6),
.Q(CLBLL_L_X4Y135_SLICE_X4Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y135_SLICE_X4Y135_CO6),
.Q(CLBLL_L_X4Y135_SLICE_X4Y135_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y135_SLICE_X4Y135_DO6),
.Q(CLBLL_L_X4Y135_SLICE_X4Y135_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc00f0aaf0aa)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_DLUT (
.I0(CLBLM_R_X5Y133_SLICE_X7Y133_AQ),
.I1(CLBLL_L_X4Y135_SLICE_X5Y135_C5Q),
.I2(CLBLM_R_X5Y136_SLICE_X7Y136_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y135_SLICE_X3Y135_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y135_SLICE_X4Y135_DO5),
.O6(CLBLL_L_X4Y135_SLICE_X4Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaff660066)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_CLUT (
.I0(CLBLM_R_X3Y135_SLICE_X3Y135_BQ),
.I1(CLBLM_R_X5Y135_SLICE_X7Y135_B5Q),
.I2(CLBLL_L_X4Y141_SLICE_X4Y141_CQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y134_SLICE_X4Y134_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y135_SLICE_X4Y135_CO5),
.O6(CLBLL_L_X4Y135_SLICE_X4Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0fff0ccf000)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y135_SLICE_X4Y135_BQ),
.I2(CLBLM_R_X3Y132_SLICE_X3Y132_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.I5(CLBLM_R_X5Y136_SLICE_X7Y136_BQ),
.O5(CLBLL_L_X4Y135_SLICE_X4Y135_BO5),
.O6(CLBLL_L_X4Y135_SLICE_X4Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8bbbbbbb88888888)
  ) CLBLL_L_X4Y135_SLICE_X4Y135_ALUT (
.I0(CLBLM_R_X5Y135_SLICE_X7Y135_CQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(LIOB33_X0Y59_IOB_X0Y60_I),
.I3(CLBLL_L_X4Y133_SLICE_X4Y133_BQ),
.I4(CLBLM_R_X5Y134_SLICE_X6Y134_C5Q),
.I5(CLBLL_L_X4Y138_SLICE_X4Y138_AO5),
.O5(CLBLL_L_X4Y135_SLICE_X4Y135_AO5),
.O6(CLBLL_L_X4Y135_SLICE_X4Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y135_SLICE_X5Y135_CO5),
.Q(CLBLL_L_X4Y135_SLICE_X5Y135_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y135_SLICE_X5Y135_AO6),
.Q(CLBLL_L_X4Y135_SLICE_X5Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y135_SLICE_X5Y135_BO6),
.Q(CLBLL_L_X4Y135_SLICE_X5Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y135_SLICE_X5Y135_CO6),
.Q(CLBLL_L_X4Y135_SLICE_X5Y135_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfbfbfbccffcc00)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_DLUT (
.I0(CLBLL_L_X4Y134_SLICE_X5Y134_AQ),
.I1(CLBLL_L_X4Y135_SLICE_X5Y135_AQ),
.I2(CLBLL_L_X4Y135_SLICE_X5Y135_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y134_SLICE_X5Y134_D5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y135_SLICE_X5Y135_DO5),
.O6(CLBLL_L_X4Y135_SLICE_X5Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88ff55aa00)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y129_SLICE_X7Y129_B5Q),
.I2(1'b1),
.I3(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I4(CLBLM_R_X5Y134_SLICE_X6Y134_DQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y135_SLICE_X5Y135_CO5),
.O6(CLBLL_L_X4Y135_SLICE_X5Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h888888888d8d888d)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y137_SLICE_X5Y137_D5Q),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLL_L_X4Y135_SLICE_X5Y135_AQ),
.I4(CLBLL_L_X4Y134_SLICE_X5Y134_AQ),
.I5(CLBLL_L_X4Y135_SLICE_X5Y135_BQ),
.O5(CLBLL_L_X4Y135_SLICE_X5Y135_BO5),
.O6(CLBLL_L_X4Y135_SLICE_X5Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h888b8b888b888b88)
  ) CLBLL_L_X4Y135_SLICE_X5Y135_ALUT (
.I0(CLBLM_R_X5Y137_SLICE_X7Y137_B5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLL_L_X4Y135_SLICE_X5Y135_AQ),
.I4(CLBLL_L_X4Y134_SLICE_X5Y134_AQ),
.I5(CLBLL_L_X4Y135_SLICE_X5Y135_BQ),
.O5(CLBLL_L_X4Y135_SLICE_X5Y135_AO5),
.O6(CLBLL_L_X4Y135_SLICE_X5Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X4Y136_AO5),
.Q(CLBLL_L_X4Y136_SLICE_X4Y136_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y138_SLICE_X4Y138_BO6),
.Q(CLBLL_L_X4Y136_SLICE_X4Y136_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X4Y136_DO5),
.Q(CLBLL_L_X4Y136_SLICE_X4Y136_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X4Y136_AO6),
.Q(CLBLL_L_X4Y136_SLICE_X4Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X4Y136_BO6),
.Q(CLBLL_L_X4Y136_SLICE_X4Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X4Y136_CO6),
.Q(CLBLL_L_X4Y136_SLICE_X4Y136_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X4Y136_DO6),
.Q(CLBLL_L_X4Y136_SLICE_X4Y136_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee2222bb88bb88)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_DLUT (
.I0(CLBLM_R_X5Y129_SLICE_X6Y129_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_CQ),
.I4(CLBLM_L_X8Y137_SLICE_X10Y137_DQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y136_SLICE_X4Y136_DO5),
.O6(CLBLL_L_X4Y136_SLICE_X4Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff19ff0c0019000c)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_CLUT (
.I0(CLBLM_R_X11Y140_SLICE_X15Y140_CO6),
.I1(CLBLL_L_X4Y136_SLICE_X4Y136_CQ),
.I2(CLBLL_L_X4Y136_SLICE_X4Y136_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y136_SLICE_X3Y136_C5Q),
.I5(CLBLL_L_X4Y136_SLICE_X4Y136_D5Q),
.O5(CLBLL_L_X4Y136_SLICE_X4Y136_CO5),
.O6(CLBLL_L_X4Y136_SLICE_X4Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffa8fc0000a8fc)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_BLUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_CQ),
.I1(CLBLL_L_X4Y136_SLICE_X4Y136_BQ),
.I2(CLBLL_L_X4Y135_SLICE_X5Y135_C5Q),
.I3(CLBLL_L_X4Y136_SLICE_X4Y136_D5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X3Y136_SLICE_X3Y136_DQ),
.O5(CLBLL_L_X4Y136_SLICE_X4Y136_BO5),
.O6(CLBLL_L_X4Y136_SLICE_X4Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0a0afc0cfc0c)
  ) CLBLL_L_X4Y136_SLICE_X4Y136_ALUT (
.I0(CLBLM_L_X8Y140_SLICE_X11Y140_DO6),
.I1(CLBLM_L_X10Y137_SLICE_X13Y137_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X3Y136_SLICE_X2Y136_A5Q),
.I4(CLBLL_L_X4Y133_SLICE_X5Y133_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y136_SLICE_X4Y136_AO5),
.O6(CLBLL_L_X4Y136_SLICE_X4Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X5Y136_DO5),
.Q(CLBLL_L_X4Y136_SLICE_X5Y136_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X5Y136_AO6),
.Q(CLBLL_L_X4Y136_SLICE_X5Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X5Y136_BO6),
.Q(CLBLL_L_X4Y136_SLICE_X5Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X5Y136_CO6),
.Q(CLBLL_L_X4Y136_SLICE_X5Y136_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y136_SLICE_X5Y136_DO6),
.Q(CLBLL_L_X4Y136_SLICE_X5Y136_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ff338888bbbb)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_DLUT (
.I0(CLBLL_L_X4Y140_SLICE_X5Y140_DQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLL_L_X4Y140_SLICE_X5Y140_CQ),
.I4(CLBLL_L_X4Y131_SLICE_X5Y131_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y136_SLICE_X5Y136_DO5),
.O6(CLBLL_L_X4Y136_SLICE_X5Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaabaf00000105)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y136_SLICE_X5Y136_CQ),
.I2(CLBLM_L_X8Y137_SLICE_X10Y137_DQ),
.I3(CLBLL_L_X4Y136_SLICE_X5Y136_BQ),
.I4(CLBLL_L_X4Y137_SLICE_X5Y137_DQ),
.I5(CLBLM_R_X7Y137_SLICE_X8Y137_D5Q),
.O5(CLBLL_L_X4Y136_SLICE_X5Y136_CO5),
.O6(CLBLL_L_X4Y136_SLICE_X5Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fffff0f0ffaa)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_BLUT (
.I0(CLBLL_L_X4Y137_SLICE_X5Y137_DQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y130_SLICE_X5Y130_B5Q),
.I3(CLBLL_L_X4Y136_SLICE_X5Y136_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X8Y137_SLICE_X10Y137_DQ),
.O5(CLBLL_L_X4Y136_SLICE_X5Y136_BO5),
.O6(CLBLL_L_X4Y136_SLICE_X5Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff78ff0000780000)
  ) CLBLL_L_X4Y136_SLICE_X5Y136_ALUT (
.I0(CLBLM_R_X3Y136_SLICE_X3Y136_AQ),
.I1(CLBLM_L_X8Y139_SLICE_X11Y139_BQ),
.I2(CLBLL_L_X4Y136_SLICE_X5Y136_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.I5(CLBLL_L_X4Y136_SLICE_X5Y136_BQ),
.O5(CLBLL_L_X4Y136_SLICE_X5Y136_AO5),
.O6(CLBLL_L_X4Y136_SLICE_X5Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y137_SLICE_X4Y137_CO5),
.Q(CLBLL_L_X4Y137_SLICE_X4Y137_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y137_SLICE_X4Y137_AO6),
.Q(CLBLL_L_X4Y137_SLICE_X4Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y137_SLICE_X4Y137_BO6),
.Q(CLBLL_L_X4Y137_SLICE_X4Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y137_SLICE_X4Y137_CO6),
.Q(CLBLL_L_X4Y137_SLICE_X4Y137_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffcc4cffff0080)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_DLUT (
.I0(CLBLM_R_X3Y135_SLICE_X3Y135_DQ),
.I1(CLBLM_R_X5Y138_SLICE_X7Y138_AQ),
.I2(CLBLM_R_X7Y138_SLICE_X9Y138_B5Q),
.I3(CLBLM_R_X5Y138_SLICE_X7Y138_CO6),
.I4(CLBLM_R_X5Y130_SLICE_X7Y130_DQ),
.I5(CLBLM_R_X5Y137_SLICE_X7Y137_BQ),
.O5(CLBLL_L_X4Y137_SLICE_X4Y137_DO5),
.O6(CLBLL_L_X4Y137_SLICE_X4Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3aca3acfafa0a0a)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_CLUT (
.I0(CLBLM_R_X3Y137_SLICE_X3Y137_AQ),
.I1(CLBLM_R_X3Y135_SLICE_X3Y135_DQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y134_SLICE_X6Y134_A5Q),
.I4(CLBLL_L_X4Y138_SLICE_X5Y138_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y137_SLICE_X4Y137_CO5),
.O6(CLBLL_L_X4Y137_SLICE_X4Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0eeeef0f000ee)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_BLUT (
.I0(CLBLL_L_X4Y135_SLICE_X4Y135_DQ),
.I1(CLBLL_L_X4Y137_SLICE_X4Y137_BQ),
.I2(CLBLL_L_X4Y137_SLICE_X5Y137_C5Q),
.I3(CLBLL_L_X4Y136_SLICE_X4Y136_D5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_CQ),
.O5(CLBLL_L_X4Y137_SLICE_X4Y137_BO5),
.O6(CLBLL_L_X4Y137_SLICE_X4Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfa00ccccfafa)
  ) CLBLL_L_X4Y137_SLICE_X4Y137_ALUT (
.I0(CLBLL_L_X4Y131_SLICE_X4Y131_DQ),
.I1(CLBLL_L_X4Y139_SLICE_X4Y139_DQ),
.I2(CLBLL_L_X4Y137_SLICE_X4Y137_AQ),
.I3(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X4Y135_SLICE_X5Y135_CQ),
.O5(CLBLL_L_X4Y137_SLICE_X4Y137_AO5),
.O6(CLBLL_L_X4Y137_SLICE_X4Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y137_SLICE_X5Y137_AO5),
.Q(CLBLL_L_X4Y137_SLICE_X5Y137_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y137_SLICE_X5Y137_BO5),
.Q(CLBLL_L_X4Y137_SLICE_X5Y137_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y137_SLICE_X5Y137_CO5),
.Q(CLBLL_L_X4Y137_SLICE_X5Y137_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y137_SLICE_X5Y137_DO5),
.Q(CLBLL_L_X4Y137_SLICE_X5Y137_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y137_SLICE_X5Y137_AO6),
.Q(CLBLL_L_X4Y137_SLICE_X5Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y137_SLICE_X5Y137_BO6),
.Q(CLBLL_L_X4Y137_SLICE_X5Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y137_SLICE_X5Y137_CO6),
.Q(CLBLL_L_X4Y137_SLICE_X5Y137_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y137_SLICE_X5Y137_DO6),
.Q(CLBLL_L_X4Y137_SLICE_X5Y137_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccaaf0fff000)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_DLUT (
.I0(CLBLM_R_X5Y133_SLICE_X7Y133_A5Q),
.I1(CLBLM_R_X5Y138_SLICE_X6Y138_BQ),
.I2(CLBLL_L_X4Y137_SLICE_X5Y137_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y138_SLICE_X5Y138_DQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y137_SLICE_X5Y137_DO5),
.O6(CLBLL_L_X4Y137_SLICE_X5Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa50d8d8dddd)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y137_SLICE_X10Y137_BQ),
.I2(CLBLM_R_X5Y130_SLICE_X7Y130_DQ),
.I3(CLBLM_R_X5Y136_SLICE_X6Y136_DQ),
.I4(CLBLL_L_X4Y137_SLICE_X5Y137_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y137_SLICE_X5Y137_CO5),
.O6(CLBLL_L_X4Y137_SLICE_X5Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfc0cfafa0a0a)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_BLUT (
.I0(CLBLL_L_X4Y137_SLICE_X5Y137_CQ),
.I1(RIOB33_X105Y119_IOB_X1Y119_I),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y138_SLICE_X9Y138_C5Q),
.I4(CLBLL_L_X4Y133_SLICE_X5Y133_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y137_SLICE_X5Y137_BO5),
.O6(CLBLL_L_X4Y137_SLICE_X5Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddddd88e4e4e4e4)
  ) CLBLL_L_X4Y137_SLICE_X5Y137_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y137_SLICE_X5Y137_BQ),
.I2(CLBLM_R_X3Y135_SLICE_X2Y135_BQ),
.I3(CLBLM_R_X5Y131_SLICE_X6Y131_BQ),
.I4(CLBLM_L_X10Y137_SLICE_X13Y137_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y137_SLICE_X5Y137_AO5),
.O6(CLBLL_L_X4Y137_SLICE_X5Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y138_SLICE_X4Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLL_L_X4Y137_SLICE_X4Y137_BQ),
.Q(CLBLL_L_X4Y138_SLICE_X4Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y138_SLICE_X4Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLL_L_X4Y138_SLICE_X5Y138_CQ),
.Q(CLBLL_L_X4Y138_SLICE_X4Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cccccccc)
  ) CLBLL_L_X4Y138_SLICE_X4Y138_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y138_SLICE_X9Y138_B5Q),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X5Y138_SLICE_X7Y138_CO6),
.O5(CLBLL_L_X4Y138_SLICE_X4Y138_DO5),
.O6(CLBLL_L_X4Y138_SLICE_X4Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffcfffc)
  ) CLBLL_L_X4Y138_SLICE_X4Y138_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y139_SLICE_X3Y139_AQ),
.I2(CLBLM_R_X5Y139_SLICE_X7Y139_A5Q),
.I3(CLBLL_L_X4Y137_SLICE_X4Y137_CQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y133_SLICE_X4Y133_C5Q),
.O5(CLBLL_L_X4Y138_SLICE_X4Y138_CO5),
.O6(CLBLL_L_X4Y138_SLICE_X4Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccaf0000f0f0)
  ) CLBLL_L_X4Y138_SLICE_X4Y138_BLUT (
.I0(CLBLM_R_X11Y141_SLICE_X14Y141_AQ),
.I1(CLBLM_R_X7Y131_SLICE_X9Y131_D5Q),
.I2(CLBLM_R_X3Y136_SLICE_X2Y136_CQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y135_SLICE_X4Y135_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y138_SLICE_X4Y138_BO5),
.O6(CLBLL_L_X4Y138_SLICE_X4Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa30aa3c3c3c3c3c)
  ) CLBLL_L_X4Y138_SLICE_X4Y138_ALUT (
.I0(CLBLM_R_X3Y137_SLICE_X3Y137_B5Q),
.I1(CLBLL_L_X4Y135_SLICE_X4Y135_AQ),
.I2(CLBLM_R_X3Y136_SLICE_X2Y136_CQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y138_SLICE_X5Y138_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y138_SLICE_X4Y138_AO5),
.O6(CLBLL_L_X4Y138_SLICE_X4Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y138_SLICE_X5Y138_AO5),
.Q(CLBLL_L_X4Y138_SLICE_X5Y138_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y138_SLICE_X6Y138_DO6),
.Q(CLBLL_L_X4Y138_SLICE_X5Y138_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y138_SLICE_X4Y138_AO6),
.Q(CLBLL_L_X4Y138_SLICE_X5Y138_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y140_SLICE_X4Y140_DO5),
.Q(CLBLL_L_X4Y138_SLICE_X5Y138_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y138_SLICE_X5Y138_AO6),
.Q(CLBLL_L_X4Y138_SLICE_X5Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y138_SLICE_X5Y138_BO6),
.Q(CLBLL_L_X4Y138_SLICE_X5Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y138_SLICE_X5Y138_CO6),
.Q(CLBLL_L_X4Y138_SLICE_X5Y138_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y138_SLICE_X5Y138_DO6),
.Q(CLBLL_L_X4Y138_SLICE_X5Y138_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccdecc00001200)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_DLUT (
.I0(CLBLM_R_X5Y138_SLICE_X6Y138_DO5),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y138_SLICE_X5Y138_DQ),
.I3(CLBLM_R_X5Y138_SLICE_X7Y138_AQ),
.I4(CLBLM_R_X5Y130_SLICE_X7Y130_DQ),
.I5(CLBLL_L_X4Y140_SLICE_X4Y140_AQ),
.O5(CLBLL_L_X4Y138_SLICE_X5Y138_DO5),
.O6(CLBLL_L_X4Y138_SLICE_X5Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf808fa0afb0bfa0a)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_CLUT (
.I0(CLBLL_L_X4Y138_SLICE_X5Y138_BQ),
.I1(CLBLL_L_X4Y135_SLICE_X4Y135_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y138_SLICE_X13Y138_DQ),
.I4(CLBLM_R_X3Y136_SLICE_X2Y136_CQ),
.I5(CLBLM_L_X10Y140_SLICE_X13Y140_B5Q),
.O5(CLBLL_L_X4Y138_SLICE_X5Y138_CO5),
.O6(CLBLL_L_X4Y138_SLICE_X5Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hecefeeee20232222)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_BLUT (
.I0(CLBLM_R_X5Y138_SLICE_X6Y138_CQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y135_SLICE_X4Y135_AQ),
.I3(CLBLM_L_X12Y136_SLICE_X16Y136_AQ),
.I4(CLBLM_R_X3Y136_SLICE_X2Y136_CQ),
.I5(CLBLM_L_X8Y140_SLICE_X11Y140_AQ),
.O5(CLBLL_L_X4Y138_SLICE_X5Y138_BO5),
.O6(CLBLL_L_X4Y138_SLICE_X5Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb88bb88c0c0f3f3)
  ) CLBLL_L_X4Y138_SLICE_X5Y138_ALUT (
.I0(CLBLM_R_X5Y139_SLICE_X6Y139_CQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y137_SLICE_X5Y137_CQ),
.I3(CLBLM_R_X3Y138_SLICE_X3Y138_CO6),
.I4(CLBLM_L_X12Y136_SLICE_X16Y136_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y138_SLICE_X5Y138_AO5),
.O6(CLBLL_L_X4Y138_SLICE_X5Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y139_SLICE_X4Y139_AO5),
.Q(CLBLL_L_X4Y139_SLICE_X4Y139_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y139_SLICE_X4Y139_AO6),
.Q(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y139_SLICE_X4Y139_BO6),
.Q(CLBLL_L_X4Y139_SLICE_X4Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y139_SLICE_X4Y139_CO6),
.Q(CLBLL_L_X4Y139_SLICE_X4Y139_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y139_SLICE_X4Y139_DO6),
.Q(CLBLL_L_X4Y139_SLICE_X4Y139_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc0a0aa0a0)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_DLUT (
.I0(CLBLM_R_X5Y141_SLICE_X7Y141_AO6),
.I1(CLBLM_R_X7Y136_SLICE_X8Y136_B5Q),
.I2(CLBLL_L_X4Y139_SLICE_X4Y139_DQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y140_SLICE_X4Y140_CO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y139_SLICE_X4Y139_DO5),
.O6(CLBLL_L_X4Y139_SLICE_X4Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff000e0e0e0e)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_CLUT (
.I0(CLBLL_L_X4Y137_SLICE_X4Y137_BQ),
.I1(CLBLL_L_X4Y139_SLICE_X4Y139_CQ),
.I2(CLBLM_L_X12Y132_SLICE_X16Y132_AO6),
.I3(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLL_L_X4Y139_SLICE_X4Y139_CO5),
.O6(CLBLL_L_X4Y139_SLICE_X4Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f0bbf0aa)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_BLUT (
.I0(CLBLM_L_X8Y140_SLICE_X10Y140_DQ),
.I1(CLBLL_L_X4Y139_SLICE_X5Y139_DO6),
.I2(CLBLL_L_X4Y138_SLICE_X5Y138_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y139_SLICE_X4Y139_BQ),
.I5(CLBLL_L_X4Y141_SLICE_X5Y141_BO6),
.O5(CLBLL_L_X4Y139_SLICE_X4Y139_BO5),
.O6(CLBLL_L_X4Y139_SLICE_X4Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8b8b8ddee1122)
  ) CLBLL_L_X4Y139_SLICE_X4Y139_ALUT (
.I0(CLBLM_R_X5Y137_SLICE_X7Y137_BQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y139_SLICE_X3Y139_BO6),
.I3(CLBLM_R_X7Y137_SLICE_X8Y137_BQ),
.I4(CLBLM_R_X3Y136_SLICE_X3Y136_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y139_SLICE_X4Y139_AO5),
.O6(CLBLL_L_X4Y139_SLICE_X4Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y139_SLICE_X5Y139_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y139_SLICE_X5Y139_CO5),
.Q(CLBLL_L_X4Y139_SLICE_X5Y139_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y139_SLICE_X5Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y139_SLICE_X5Y139_AO6),
.Q(CLBLL_L_X4Y139_SLICE_X5Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y139_SLICE_X5Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y139_SLICE_X5Y139_BO6),
.Q(CLBLL_L_X4Y139_SLICE_X5Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y139_SLICE_X5Y139_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y139_SLICE_X5Y139_CO6),
.Q(CLBLL_L_X4Y139_SLICE_X5Y139_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033003350505050)
  ) CLBLL_L_X4Y139_SLICE_X5Y139_DLUT (
.I0(CLBLM_R_X7Y140_SLICE_X8Y140_C5Q),
.I1(CLBLM_R_X3Y139_SLICE_X2Y139_AQ),
.I2(CLBLM_R_X5Y129_SLICE_X7Y129_B5Q),
.I3(CLBLM_R_X3Y139_SLICE_X2Y139_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y139_SLICE_X5Y139_DO5),
.O6(CLBLL_L_X4Y139_SLICE_X5Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0f0faaaaf0f0)
  ) CLBLL_L_X4Y139_SLICE_X5Y139_CLUT (
.I0(CLBLM_R_X5Y139_SLICE_X7Y139_BQ),
.I1(CLBLM_L_X8Y135_SLICE_X11Y135_AQ),
.I2(CLBLM_R_X5Y140_SLICE_X7Y140_B5Q),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y139_SLICE_X5Y139_CO5),
.O6(CLBLL_L_X4Y139_SLICE_X5Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44fa50fa50)
  ) CLBLL_L_X4Y139_SLICE_X5Y139_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y139_SLICE_X5Y139_BQ),
.I2(CLBLL_L_X4Y140_SLICE_X5Y140_AQ),
.I3(CLBLM_R_X3Y139_SLICE_X2Y139_AQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.O5(CLBLL_L_X4Y139_SLICE_X5Y139_BO5),
.O6(CLBLL_L_X4Y139_SLICE_X5Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haafcaafcaa00aafc)
  ) CLBLL_L_X4Y139_SLICE_X5Y139_ALUT (
.I0(CLBLM_R_X5Y130_SLICE_X6Y130_B5Q),
.I1(CLBLM_R_X7Y138_SLICE_X9Y138_C5Q),
.I2(CLBLL_L_X4Y139_SLICE_X5Y139_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y136_SLICE_X4Y136_D5Q),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_CQ),
.O5(CLBLL_L_X4Y139_SLICE_X5Y139_AO5),
.O6(CLBLL_L_X4Y139_SLICE_X5Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X5Y133_SLICE_X7Y133_AQ),
.Q(CLBLL_L_X4Y140_SLICE_X4Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5f5ccccf5f5)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_DLUT (
.I0(CLBLL_L_X4Y138_SLICE_X5Y138_C5Q),
.I1(CLBLL_L_X4Y139_SLICE_X4Y139_A5Q),
.I2(CLBLL_L_X4Y140_SLICE_X4Y140_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X4Y140_DO5),
.O6(CLBLL_L_X4Y140_SLICE_X4Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h300030005fffffff)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_CLUT (
.I0(CLBLL_L_X4Y139_SLICE_X4Y139_DQ),
.I1(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.I2(CLBLL_L_X4Y141_SLICE_X4Y141_DQ),
.I3(CLBLM_R_X3Y140_SLICE_X3Y140_DQ),
.I4(CLBLL_L_X4Y140_SLICE_X5Y140_DQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X4Y140_CO5),
.O6(CLBLL_L_X4Y140_SLICE_X4Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2d0f0f0f20000000)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_BLUT (
.I0(CLBLL_L_X4Y141_SLICE_X4Y141_DQ),
.I1(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.I2(CLBLL_L_X4Y140_SLICE_X5Y140_DQ),
.I3(CLBLM_R_X3Y140_SLICE_X3Y140_DQ),
.I4(CLBLL_L_X4Y139_SLICE_X4Y139_DQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X4Y140_BO5),
.O6(CLBLL_L_X4Y140_SLICE_X4Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ee22ff000000)
  ) CLBLL_L_X4Y140_SLICE_X4Y140_ALUT (
.I0(CLBLL_L_X4Y131_SLICE_X5Y131_B5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLL_L_X4Y141_SLICE_X4Y141_BQ),
.I4(CLBLL_L_X4Y141_SLICE_X4Y141_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X4Y140_AO5),
.O6(CLBLL_L_X4Y140_SLICE_X4Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y140_SLICE_X5Y140_CO5),
.Q(CLBLL_L_X4Y140_SLICE_X5Y140_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y140_SLICE_X5Y140_AO6),
.Q(CLBLL_L_X4Y140_SLICE_X5Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y140_SLICE_X5Y140_BO6),
.Q(CLBLL_L_X4Y140_SLICE_X5Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y140_SLICE_X5Y140_CO6),
.Q(CLBLL_L_X4Y140_SLICE_X5Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y140_SLICE_X5Y140_DO6),
.Q(CLBLL_L_X4Y140_SLICE_X5Y140_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0afa0a0a0afa0a0)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_DLUT (
.I0(CLBLL_L_X4Y139_SLICE_X5Y139_AQ),
.I1(1'b1),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y140_SLICE_X4Y140_BO6),
.I4(CLBLM_R_X5Y141_SLICE_X7Y141_AO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X5Y140_DO5),
.O6(CLBLL_L_X4Y140_SLICE_X5Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccaaccaacc)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_CLUT (
.I0(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.I1(CLBLL_L_X4Y138_SLICE_X5Y138_DQ),
.I2(CLBLL_L_X4Y134_SLICE_X5Y134_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y140_SLICE_X5Y140_CO5),
.O6(CLBLL_L_X4Y140_SLICE_X5Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h88bb888888888888)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_BLUT (
.I0(CLBLL_L_X4Y136_SLICE_X4Y136_DQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I4(CLBLM_R_X3Y135_SLICE_X2Y135_AQ),
.I5(CLBLL_L_X4Y141_SLICE_X5Y141_CO6),
.O5(CLBLL_L_X4Y140_SLICE_X5Y140_BO5),
.O6(CLBLL_L_X4Y140_SLICE_X5Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccaaccf0ccf0)
  ) CLBLL_L_X4Y140_SLICE_X5Y140_ALUT (
.I0(CLBLL_L_X4Y136_SLICE_X4Y136_DQ),
.I1(CLBLL_L_X4Y138_SLICE_X5Y138_B5Q),
.I2(CLBLL_L_X4Y140_SLICE_X5Y140_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y135_SLICE_X9Y135_C5Q),
.I5(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.O5(CLBLL_L_X4Y140_SLICE_X5Y140_AO5),
.O6(CLBLL_L_X4Y140_SLICE_X5Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y141_SLICE_X4Y141_AO6),
.Q(CLBLL_L_X4Y141_SLICE_X4Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y141_SLICE_X4Y141_BO6),
.Q(CLBLL_L_X4Y141_SLICE_X4Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y141_SLICE_X4Y141_CO6),
.Q(CLBLL_L_X4Y141_SLICE_X4Y141_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y141_SLICE_X4Y141_DO6),
.Q(CLBLL_L_X4Y141_SLICE_X4Y141_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff82a0000082a0)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_DLUT (
.I0(CLBLM_R_X5Y141_SLICE_X7Y141_AO6),
.I1(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.I2(CLBLL_L_X4Y141_SLICE_X4Y141_DQ),
.I3(CLBLM_R_X3Y140_SLICE_X3Y140_DQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X4Y130_SLICE_X4Y130_D5Q),
.O5(CLBLL_L_X4Y141_SLICE_X4Y141_DO5),
.O6(CLBLL_L_X4Y141_SLICE_X4Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ffb0bff0ff303)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_CLUT (
.I0(CLBLL_L_X4Y141_SLICE_X4Y141_BQ),
.I1(CLBLL_L_X4Y141_SLICE_X4Y141_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y138_SLICE_X5Y138_A5Q),
.I4(CLBLM_R_X5Y142_SLICE_X6Y142_B5Q),
.I5(CLBLL_L_X4Y141_SLICE_X4Y141_AQ),
.O5(CLBLL_L_X4Y141_SLICE_X4Y141_CO5),
.O6(CLBLL_L_X4Y141_SLICE_X4Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff101400001014)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_BLUT (
.I0(CLBLM_R_X5Y142_SLICE_X6Y142_B5Q),
.I1(CLBLL_L_X4Y141_SLICE_X4Y141_BQ),
.I2(CLBLL_L_X4Y141_SLICE_X4Y141_CQ),
.I3(CLBLL_L_X4Y141_SLICE_X4Y141_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X4Y136_SLICE_X4Y136_CQ),
.O5(CLBLL_L_X4Y141_SLICE_X4Y141_BO5),
.O6(CLBLL_L_X4Y141_SLICE_X4Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f01111f0f04400)
  ) CLBLL_L_X4Y141_SLICE_X4Y141_ALUT (
.I0(CLBLM_R_X5Y142_SLICE_X6Y142_B5Q),
.I1(CLBLL_L_X4Y141_SLICE_X4Y141_BQ),
.I2(CLBLM_R_X3Y139_SLICE_X3Y139_AQ),
.I3(CLBLL_L_X4Y141_SLICE_X4Y141_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X4Y141_SLICE_X4Y141_AQ),
.O5(CLBLL_L_X4Y141_SLICE_X4Y141_AO5),
.O6(CLBLL_L_X4Y141_SLICE_X4Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y141_SLICE_X5Y141_AO6),
.Q(CLBLL_L_X4Y141_SLICE_X5Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cccccccc)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y140_SLICE_X10Y140_C5Q),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X7Y137_SLICE_X8Y137_C5Q),
.O5(CLBLL_L_X4Y141_SLICE_X5Y141_DO5),
.O6(CLBLL_L_X4Y141_SLICE_X5Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cc00cc00)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I2(1'b1),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y140_SLICE_X10Y140_DQ),
.O5(CLBLL_L_X4Y141_SLICE_X5Y141_CO5),
.O6(CLBLL_L_X4Y141_SLICE_X5Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55df55dfdfdfdfdf)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_L_X8Y140_SLICE_X10Y140_DQ),
.I2(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.I3(CLBLM_R_X3Y135_SLICE_X2Y135_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y141_SLICE_X5Y141_BO5),
.O6(CLBLL_L_X4Y141_SLICE_X5Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'habba0110effe4554)
  ) CLBLL_L_X4Y141_SLICE_X5Y141_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y141_SLICE_X7Y141_AO5),
.I2(CLBLL_L_X4Y141_SLICE_X5Y141_AQ),
.I3(CLBLM_R_X5Y141_SLICE_X7Y141_BO6),
.I4(CLBLM_R_X5Y136_SLICE_X6Y136_AQ),
.I5(CLBLM_L_X10Y130_SLICE_X12Y130_B5Q),
.O5(CLBLL_L_X4Y141_SLICE_X5Y141_AO5),
.O6(CLBLL_L_X4Y141_SLICE_X5Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y142_SLICE_X4Y142_BO5),
.Q(CLBLL_L_X4Y142_SLICE_X4Y142_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y142_SLICE_X4Y142_AO6),
.Q(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y142_SLICE_X4Y142_DO5),
.O6(CLBLL_L_X4Y142_SLICE_X4Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y142_SLICE_X4Y142_CO5),
.O6(CLBLL_L_X4Y142_SLICE_X4Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00fffa50fa50)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLM_L_X12Y141_SLICE_X16Y141_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y142_SLICE_X4Y142_BO5),
.O6(CLBLL_L_X4Y142_SLICE_X4Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haffa0550aaaa0000)
  ) CLBLL_L_X4Y142_SLICE_X4Y142_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.I3(CLBLL_L_X4Y143_SLICE_X5Y143_BO5),
.I4(CLBLL_L_X4Y139_SLICE_X5Y139_BQ),
.I5(CLBLM_R_X5Y141_SLICE_X7Y141_AO6),
.O5(CLBLL_L_X4Y142_SLICE_X4Y142_AO5),
.O6(CLBLL_L_X4Y142_SLICE_X4Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y142_SLICE_X5Y142_CO6),
.Q(CLBLL_L_X4Y142_SLICE_X5Y142_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y142_SLICE_X5Y142_AO6),
.Q(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y142_SLICE_X5Y142_BO6),
.Q(CLBLL_L_X4Y142_SLICE_X5Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0200000000000000)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_DLUT (
.I0(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.I1(CLBLL_L_X4Y140_SLICE_X4Y140_CO5),
.I2(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.I3(CLBLL_L_X4Y142_SLICE_X5Y142_A5Q),
.I4(CLBLM_R_X5Y141_SLICE_X6Y141_DQ),
.I5(CLBLM_R_X5Y142_SLICE_X6Y142_CQ),
.O5(CLBLL_L_X4Y142_SLICE_X5Y142_DO5),
.O6(CLBLL_L_X4Y142_SLICE_X5Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0cc055555555)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_CLUT (
.I0(CLBLL_L_X4Y141_SLICE_X5Y141_AQ),
.I1(CLBLM_R_X5Y141_SLICE_X7Y141_AO6),
.I2(CLBLL_L_X4Y140_SLICE_X4Y140_BO5),
.I3(CLBLL_L_X4Y142_SLICE_X5Y142_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y142_SLICE_X5Y142_CO5),
.O6(CLBLL_L_X4Y142_SLICE_X5Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf6f00600f6f00600)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_BLUT (
.I0(CLBLL_L_X4Y142_SLICE_X5Y142_DO6),
.I1(CLBLL_L_X4Y142_SLICE_X5Y142_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y141_SLICE_X7Y141_AO6),
.I4(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y142_SLICE_X5Y142_BO5),
.O6(CLBLL_L_X4Y142_SLICE_X5Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3333deee1222)
  ) CLBLL_L_X4Y142_SLICE_X5Y142_ALUT (
.I0(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLL_L_X4Y141_SLICE_X4Y141_AQ),
.I3(CLBLL_L_X4Y141_SLICE_X4Y141_BQ),
.I4(CLBLM_R_X5Y135_SLICE_X6Y135_B5Q),
.I5(CLBLM_R_X5Y142_SLICE_X6Y142_B5Q),
.O5(CLBLL_L_X4Y142_SLICE_X5Y142_AO5),
.O6(CLBLL_L_X4Y142_SLICE_X5Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y143_SLICE_X4Y143_DO5),
.O6(CLBLL_L_X4Y143_SLICE_X4Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y143_SLICE_X4Y143_CO5),
.O6(CLBLL_L_X4Y143_SLICE_X4Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y143_SLICE_X4Y143_BO5),
.O6(CLBLL_L_X4Y143_SLICE_X4Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f5f5f5f5f)
  ) CLBLL_L_X4Y143_SLICE_X4Y143_ALUT (
.I0(CLBLM_R_X5Y141_SLICE_X6Y141_CQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y136_SLICE_X5Y136_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y143_SLICE_X4Y143_AO5),
.O6(CLBLL_L_X4Y143_SLICE_X4Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y143_SLICE_X5Y143_AO6),
.Q(CLBLL_L_X4Y143_SLICE_X5Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777ffffffffffff)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_DLUT (
.I0(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.I1(CLBLM_R_X5Y142_SLICE_X6Y142_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X4Y143_SLICE_X5Y143_AQ),
.I5(CLBLL_L_X4Y142_SLICE_X5Y142_BQ),
.O5(CLBLL_L_X4Y143_SLICE_X5Y143_DO5),
.O6(CLBLL_L_X4Y143_SLICE_X5Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0800000000000000)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_CLUT (
.I0(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.I1(CLBLM_R_X5Y142_SLICE_X6Y142_CQ),
.I2(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.I3(CLBLL_L_X4Y142_SLICE_X5Y142_BQ),
.I4(CLBLL_L_X4Y143_SLICE_X5Y143_AQ),
.I5(CLBLM_R_X5Y142_SLICE_X7Y142_BO6),
.O5(CLBLL_L_X4Y143_SLICE_X5Y143_CO5),
.O6(CLBLL_L_X4Y143_SLICE_X5Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4000000044000000)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_BLUT (
.I0(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.I1(CLBLM_R_X5Y142_SLICE_X6Y142_CQ),
.I2(CLBLL_L_X4Y142_SLICE_X4Y142_AQ),
.I3(CLBLL_L_X4Y142_SLICE_X5Y142_BQ),
.I4(CLBLM_R_X5Y142_SLICE_X7Y142_BO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y143_SLICE_X5Y143_BO5),
.O6(CLBLL_L_X4Y143_SLICE_X5Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haeeaaeea04400440)
  ) CLBLL_L_X4Y143_SLICE_X5Y143_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y141_SLICE_X7Y141_AO6),
.I2(CLBLL_L_X4Y143_SLICE_X5Y143_AQ),
.I3(CLBLL_L_X4Y143_SLICE_X5Y143_BO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y140_SLICE_X9Y140_CQ),
.O5(CLBLL_L_X4Y143_SLICE_X5Y143_AO5),
.O6(CLBLL_L_X4Y143_SLICE_X5Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y130_SLICE_X10Y130_AO6),
.Q(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000800000000000)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_DLUT (
.I0(CLBLM_L_X8Y138_SLICE_X11Y138_AQ),
.I1(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I2(CLBLM_L_X8Y131_SLICE_X11Y131_BQ),
.I3(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y130_SLICE_X8Y130_DO6),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_DO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_CLUT (
.I0(CLBLM_L_X8Y138_SLICE_X11Y138_AQ),
.I1(CLBLM_L_X8Y131_SLICE_X11Y131_BQ),
.I2(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.I3(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.I4(CLBLM_R_X7Y130_SLICE_X8Y130_CO6),
.I5(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_CO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_BLUT (
.I0(CLBLM_L_X8Y131_SLICE_X11Y131_BQ),
.I1(CLBLM_L_X8Y138_SLICE_X11Y138_AQ),
.I2(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I3(CLBLM_L_X8Y131_SLICE_X10Y131_BQ),
.I4(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.I5(CLBLM_R_X7Y130_SLICE_X8Y130_DO6),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_BO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaacc0fccaaccf0)
  ) CLBLM_L_X8Y130_SLICE_X10Y130_ALUT (
.I0(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I1(CLBLL_L_X4Y134_SLICE_X5Y134_D5Q),
.I2(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y133_SLICE_X6Y133_A5Q),
.I5(CLBLM_L_X8Y130_SLICE_X10Y130_CO6),
.O5(CLBLM_L_X8Y130_SLICE_X10Y130_AO5),
.O6(CLBLM_L_X8Y130_SLICE_X10Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_DO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a00000000000000)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_CLUT (
.I0(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y134_SLICE_X8Y134_DO6),
.I3(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.I4(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.I5(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_CO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000080000000)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_BLUT (
.I0(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I1(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I2(CLBLM_L_X8Y138_SLICE_X11Y138_AQ),
.I3(CLBLM_L_X8Y131_SLICE_X10Y131_BQ),
.I4(CLBLM_L_X8Y130_SLICE_X11Y130_AO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_BO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000800000000000)
  ) CLBLM_L_X8Y130_SLICE_X11Y130_ALUT (
.I0(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.I1(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.I2(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.I3(CLBLM_L_X8Y131_SLICE_X11Y131_BQ),
.I4(CLBLM_R_X7Y134_SLICE_X8Y134_DO6),
.I5(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.O5(CLBLM_L_X8Y130_SLICE_X11Y130_AO5),
.O6(CLBLM_L_X8Y130_SLICE_X11Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X10Y131_AO6),
.Q(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X10Y131_BO6),
.Q(CLBLM_L_X8Y131_SLICE_X10Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X10Y131_CO6),
.Q(CLBLM_L_X8Y131_SLICE_X10Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_DO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fffc00000f0c)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y131_SLICE_X10Y131_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y131_SLICE_X9Y131_BQ),
.I4(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.I5(CLBLM_L_X8Y137_SLICE_X11Y137_D5Q),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_CO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heafb4051fbea5140)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y133_SLICE_X6Y133_A5Q),
.I2(CLBLM_L_X8Y137_SLICE_X10Y137_C5Q),
.I3(CLBLM_L_X8Y130_SLICE_X10Y130_DO6),
.I4(CLBLM_L_X8Y140_SLICE_X10Y140_C5Q),
.I5(CLBLM_L_X8Y131_SLICE_X10Y131_BQ),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_BO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffcca50000cca5)
  ) CLBLM_L_X8Y131_SLICE_X10Y131_ALUT (
.I0(CLBLM_R_X7Y134_SLICE_X8Y134_DO6),
.I1(CLBLM_L_X8Y138_SLICE_X11Y138_BQ),
.I2(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.I3(CLBLM_R_X5Y133_SLICE_X6Y133_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.O5(CLBLM_L_X8Y131_SLICE_X10Y131_AO5),
.O6(CLBLM_L_X8Y131_SLICE_X10Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X11Y131_CO5),
.Q(CLBLM_L_X8Y131_SLICE_X11Y131_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X11Y131_DO5),
.Q(CLBLM_L_X8Y131_SLICE_X11Y131_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X11Y131_AO6),
.Q(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X11Y131_BO6),
.Q(CLBLM_L_X8Y131_SLICE_X11Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X11Y131_CO6),
.Q(CLBLM_L_X8Y131_SLICE_X11Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y131_SLICE_X11Y131_DO6),
.Q(CLBLM_L_X8Y131_SLICE_X11Y131_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccaaffaa00aa)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_DLUT (
.I0(CLBLM_R_X3Y135_SLICE_X3Y135_DQ),
.I1(CLBLM_L_X8Y133_SLICE_X11Y133_AQ),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_DO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000ff0fc0c0cfcf)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y131_SLICE_X10Y131_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y136_SLICE_X5Y136_DQ),
.I4(CLBLL_L_X4Y131_SLICE_X5Y131_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_CO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfabb5011faee5044)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y131_SLICE_X11Y131_BQ),
.I2(CLBLM_R_X5Y133_SLICE_X7Y133_C5Q),
.I3(CLBLM_R_X5Y133_SLICE_X6Y133_A5Q),
.I4(CLBLM_L_X10Y136_SLICE_X13Y136_BQ),
.I5(CLBLM_L_X8Y130_SLICE_X11Y130_CO6),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_BO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb8b888bbbb888b8)
  ) CLBLM_L_X8Y131_SLICE_X11Y131_ALUT (
.I0(CLBLM_R_X7Y133_SLICE_X9Y133_DQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X8Y130_SLICE_X10Y130_BO6),
.I3(CLBLM_R_X5Y133_SLICE_X6Y133_A5Q),
.I4(CLBLM_L_X10Y131_SLICE_X12Y131_C5Q),
.I5(CLBLM_L_X8Y131_SLICE_X11Y131_AQ),
.O5(CLBLM_L_X8Y131_SLICE_X11Y131_AO5),
.O6(CLBLM_L_X8Y131_SLICE_X11Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y132_SLICE_X10Y132_AO5),
.Q(CLBLM_L_X8Y132_SLICE_X10Y132_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y132_SLICE_X10Y132_BO5),
.Q(CLBLM_L_X8Y132_SLICE_X10Y132_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y132_SLICE_X10Y132_AO6),
.Q(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y132_SLICE_X10Y132_BO6),
.Q(CLBLM_L_X8Y132_SLICE_X10Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y132_SLICE_X10Y132_CO6),
.Q(CLBLM_L_X8Y132_SLICE_X10Y132_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000018081000)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_DLUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I1(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I2(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I3(CLBLM_L_X8Y131_SLICE_X10Y131_CQ),
.I4(CLBLM_R_X7Y132_SLICE_X9Y132_AQ),
.I5(CLBLM_R_X11Y132_SLICE_X15Y132_AO5),
.O5(CLBLM_L_X8Y132_SLICE_X10Y132_DO5),
.O6(CLBLM_L_X8Y132_SLICE_X10Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff55f0f0cc44)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_CLUT (
.I0(CLBLM_R_X7Y131_SLICE_X9Y131_D5Q),
.I1(CLBLM_L_X8Y132_SLICE_X10Y132_CQ),
.I2(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.I3(CLBLM_L_X10Y140_SLICE_X13Y140_D5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y135_SLICE_X9Y135_D5Q),
.O5(CLBLM_L_X8Y132_SLICE_X10Y132_CO5),
.O6(CLBLM_L_X8Y132_SLICE_X10Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf055f055cc55cc55)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_BLUT (
.I0(CLBLM_L_X10Y140_SLICE_X13Y140_B5Q),
.I1(CLBLL_L_X4Y131_SLICE_X4Y131_CQ),
.I2(CLBLM_L_X10Y134_SLICE_X12Y134_B5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y132_SLICE_X10Y132_BO5),
.O6(CLBLM_L_X8Y132_SLICE_X10Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88dd88dda0f5a0f5)
  ) CLBLM_L_X8Y132_SLICE_X10Y132_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y132_SLICE_X9Y132_CQ),
.I2(CLBLL_L_X4Y136_SLICE_X4Y136_B5Q),
.I3(CLBLM_R_X11Y142_SLICE_X14Y142_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y132_SLICE_X10Y132_AO5),
.O6(CLBLM_L_X8Y132_SLICE_X10Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y132_SLICE_X11Y132_AO6),
.Q(CLBLM_L_X8Y132_SLICE_X11Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y132_SLICE_X11Y132_BO6),
.Q(CLBLM_L_X8Y132_SLICE_X11Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6f6ff6f66f6ff6f6)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_DLUT (
.I0(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I1(CLBLL_L_X4Y132_SLICE_X4Y132_DQ),
.I2(CLBLM_R_X3Y132_SLICE_X3Y132_CQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y132_SLICE_X5Y132_DQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y132_SLICE_X11Y132_DO5),
.O6(CLBLM_L_X8Y132_SLICE_X11Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800000088000000)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_CLUT (
.I0(CLBLM_L_X8Y132_SLICE_X11Y132_BQ),
.I1(CLBLM_L_X10Y132_SLICE_X12Y132_AQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y135_SLICE_X11Y135_BO6),
.I4(CLBLM_L_X8Y132_SLICE_X11Y132_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y132_SLICE_X11Y132_CO5),
.O6(CLBLM_L_X8Y132_SLICE_X11Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hae04ea40ee44aa00)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.I2(CLBLM_L_X10Y132_SLICE_X12Y132_AQ),
.I3(CLBLM_L_X8Y135_SLICE_X10Y135_C5Q),
.I4(CLBLM_L_X8Y132_SLICE_X11Y132_BQ),
.I5(CLBLM_L_X8Y132_SLICE_X11Y132_AO5),
.O5(CLBLM_L_X8Y132_SLICE_X11Y132_BO5),
.O6(CLBLM_L_X8Y132_SLICE_X11Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdecc1200a0a0a0a0)
  ) CLBLM_L_X8Y132_SLICE_X11Y132_ALUT (
.I0(CLBLM_L_X8Y135_SLICE_X11Y135_BO6),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X8Y132_SLICE_X11Y132_AQ),
.I3(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.I4(CLBLM_L_X10Y134_SLICE_X12Y134_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y132_SLICE_X11Y132_AO5),
.O6(CLBLM_L_X8Y132_SLICE_X11Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y133_SLICE_X10Y133_CO5),
.Q(CLBLM_L_X8Y133_SLICE_X10Y133_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y133_SLICE_X10Y133_AO6),
.Q(CLBLM_L_X8Y133_SLICE_X10Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y133_SLICE_X10Y133_BO6),
.Q(CLBLM_L_X8Y133_SLICE_X10Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y133_SLICE_X10Y133_CO6),
.Q(CLBLM_L_X8Y133_SLICE_X10Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdcffffffdcffdc)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_DLUT (
.I0(CLBLM_L_X8Y136_SLICE_X11Y136_CO5),
.I1(CLBLM_L_X8Y134_SLICE_X10Y134_CO6),
.I2(CLBLM_L_X8Y132_SLICE_X10Y132_A5Q),
.I3(CLBLM_L_X8Y132_SLICE_X10Y132_DO6),
.I4(CLBLM_R_X11Y133_SLICE_X14Y133_CO5),
.I5(CLBLM_R_X5Y132_SLICE_X7Y132_BQ),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_DO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff00ff00e4e4)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_CLUT (
.I0(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.I1(CLBLM_L_X8Y132_SLICE_X10Y132_CQ),
.I2(CLBLM_L_X8Y133_SLICE_X10Y133_C5Q),
.I3(CLBLM_R_X5Y134_SLICE_X6Y134_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_CO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0aaff88cc)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_BLUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_CQ),
.I1(CLBLM_L_X8Y133_SLICE_X10Y133_BQ),
.I2(CLBLM_L_X10Y132_SLICE_X12Y132_BQ),
.I3(CLBLL_L_X4Y136_SLICE_X4Y136_D5Q),
.I4(CLBLM_R_X5Y131_SLICE_X7Y131_D5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_BO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00aaaae2e2)
  ) CLBLM_L_X8Y133_SLICE_X10Y133_ALUT (
.I0(CLBLM_L_X8Y131_SLICE_X11Y131_DQ),
.I1(CLBLL_L_X4Y136_SLICE_X4Y136_D5Q),
.I2(CLBLM_L_X8Y133_SLICE_X10Y133_AQ),
.I3(CLBLM_L_X10Y134_SLICE_X13Y134_AQ),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_CQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y133_SLICE_X10Y133_AO5),
.O6(CLBLM_L_X8Y133_SLICE_X10Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y133_SLICE_X11Y133_AO5),
.Q(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y133_SLICE_X11Y133_BO5),
.Q(CLBLM_L_X8Y133_SLICE_X11Y133_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y133_SLICE_X11Y133_AO6),
.Q(CLBLM_L_X8Y133_SLICE_X11Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y133_SLICE_X11Y133_BO6),
.Q(CLBLM_L_X8Y133_SLICE_X11Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3ff3cffc3ff3cffc)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y132_SLICE_X4Y132_DQ),
.I2(CLBLM_R_X3Y132_SLICE_X3Y132_CQ),
.I3(CLBLM_R_X5Y133_SLICE_X7Y133_B5Q),
.I4(CLBLM_R_X7Y134_SLICE_X8Y134_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_DO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h008c008c00800080)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_CLUT (
.I0(CLBLM_R_X7Y133_SLICE_X9Y133_C5Q),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I2(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I3(CLBLM_L_X10Y133_SLICE_X12Y133_CO6),
.I4(1'b1),
.I5(CLBLM_L_X8Y137_SLICE_X11Y137_D5Q),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_CO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff660066f0aaf0aa)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_BLUT (
.I0(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.I1(CLBLM_R_X5Y137_SLICE_X7Y137_AQ),
.I2(CLBLM_R_X5Y130_SLICE_X7Y130_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y136_SLICE_X12Y136_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_BO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccaaffaa00)
  ) CLBLM_L_X8Y133_SLICE_X11Y133_ALUT (
.I0(CLBLM_L_X8Y137_SLICE_X11Y137_CQ),
.I1(CLBLM_L_X10Y134_SLICE_X13Y134_AQ),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y137_SLICE_X4Y137_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y133_SLICE_X11Y133_AO5),
.O6(CLBLM_L_X8Y133_SLICE_X11Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y134_SLICE_X10Y134_AO5),
.Q(CLBLM_L_X8Y134_SLICE_X10Y134_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y134_SLICE_X10Y134_AO6),
.Q(CLBLM_L_X8Y134_SLICE_X10Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff6f6ffffff6f6)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_DLUT (
.I0(CLBLM_L_X10Y132_SLICE_X12Y132_AQ),
.I1(CLBLM_R_X7Y136_SLICE_X8Y136_BQ),
.I2(CLBLM_R_X7Y136_SLICE_X9Y136_CQ),
.I3(1'b1),
.I4(CLBLM_R_X3Y136_SLICE_X3Y136_AQ),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_A5Q),
.O5(CLBLM_L_X8Y134_SLICE_X10Y134_DO5),
.O6(CLBLM_L_X8Y134_SLICE_X10Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5404050554040000)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_CLUT (
.I0(CLBLM_R_X11Y133_SLICE_X15Y133_AO6),
.I1(CLBLM_R_X7Y132_SLICE_X9Y132_A5Q),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I3(CLBLM_R_X7Y136_SLICE_X9Y136_A5Q),
.I4(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I5(CLBLM_R_X5Y134_SLICE_X6Y134_A5Q),
.O5(CLBLM_L_X8Y134_SLICE_X10Y134_CO5),
.O6(CLBLM_L_X8Y134_SLICE_X10Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffbfffe)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_BLUT (
.I0(CLBLM_L_X8Y136_SLICE_X10Y136_DO6),
.I1(CLBLM_L_X8Y132_SLICE_X11Y132_BQ),
.I2(CLBLM_L_X8Y132_SLICE_X11Y132_DO6),
.I3(CLBLM_L_X8Y134_SLICE_X10Y134_DO6),
.I4(CLBLM_R_X7Y132_SLICE_X9Y132_DQ),
.I5(CLBLM_L_X8Y134_SLICE_X11Y134_DO6),
.O5(CLBLM_L_X8Y134_SLICE_X10Y134_BO5),
.O6(CLBLM_L_X8Y134_SLICE_X10Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaccf0ccf0cc)
  ) CLBLM_L_X8Y134_SLICE_X10Y134_ALUT (
.I0(CLBLL_L_X4Y139_SLICE_X5Y139_CQ),
.I1(CLBLM_R_X11Y141_SLICE_X14Y141_AQ),
.I2(CLBLM_L_X8Y136_SLICE_X11Y136_B5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y134_SLICE_X10Y134_AO5),
.O6(CLBLM_L_X8Y134_SLICE_X10Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y134_SLICE_X11Y134_BO5),
.Q(CLBLM_L_X8Y134_SLICE_X11Y134_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y134_SLICE_X11Y134_AO6),
.Q(CLBLM_L_X8Y134_SLICE_X11Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y134_SLICE_X11Y134_BO6),
.Q(CLBLM_L_X8Y134_SLICE_X11Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5ff55ff5affaaffa)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_DLUT (
.I0(CLBLL_L_X4Y136_SLICE_X5Y136_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y137_SLICE_X8Y137_B5Q),
.I3(CLBLM_L_X8Y132_SLICE_X11Y132_AQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y136_SLICE_X6Y136_BQ),
.O5(CLBLM_L_X8Y134_SLICE_X11Y134_DO5),
.O6(CLBLM_L_X8Y134_SLICE_X11Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff7fffffffb)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_CLUT (
.I0(CLBLM_R_X3Y133_SLICE_X3Y133_BQ),
.I1(CLBLM_L_X8Y135_SLICE_X11Y135_CO6),
.I2(CLBLM_L_X10Y134_SLICE_X12Y134_DO6),
.I3(CLBLM_L_X8Y135_SLICE_X11Y135_DO6),
.I4(CLBLM_L_X8Y133_SLICE_X11Y133_DO6),
.I5(CLBLM_L_X8Y132_SLICE_X11Y132_AQ),
.O5(CLBLM_L_X8Y134_SLICE_X11Y134_CO5),
.O6(CLBLM_L_X8Y134_SLICE_X11Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aafff000f0)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_BLUT (
.I0(CLBLM_R_X7Y140_SLICE_X9Y140_D5Q),
.I1(1'b1),
.I2(CLBLM_R_X7Y133_SLICE_X9Y133_C5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y133_SLICE_X7Y133_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y134_SLICE_X11Y134_BO5),
.O6(CLBLM_L_X8Y134_SLICE_X11Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaccc0fff0)
  ) CLBLM_L_X8Y134_SLICE_X11Y134_ALUT (
.I0(CLBLM_R_X3Y134_SLICE_X3Y134_BQ),
.I1(CLBLM_L_X10Y140_SLICE_X13Y140_D5Q),
.I2(CLBLM_L_X8Y134_SLICE_X11Y134_AQ),
.I3(CLBLM_R_X7Y136_SLICE_X9Y136_D5Q),
.I4(CLBLM_R_X7Y131_SLICE_X9Y131_D5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y134_SLICE_X11Y134_AO5),
.O6(CLBLM_L_X8Y134_SLICE_X11Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y135_SLICE_X10Y135_BO5),
.Q(CLBLM_L_X8Y135_SLICE_X10Y135_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y135_SLICE_X10Y135_CO5),
.Q(CLBLM_L_X8Y135_SLICE_X10Y135_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y135_SLICE_X10Y135_DO5),
.Q(CLBLM_L_X8Y135_SLICE_X10Y135_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y135_SLICE_X10Y135_AO6),
.Q(CLBLM_L_X8Y135_SLICE_X10Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y135_SLICE_X10Y135_BO6),
.Q(CLBLM_L_X8Y135_SLICE_X10Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y135_SLICE_X10Y135_CO6),
.Q(CLBLM_L_X8Y135_SLICE_X10Y135_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y135_SLICE_X10Y135_DO6),
.Q(CLBLM_L_X8Y135_SLICE_X10Y135_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h88dddd88f5f5a0a0)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y131_SLICE_X11Y131_DQ),
.I2(CLBLM_R_X7Y135_SLICE_X9Y135_CQ),
.I3(CLBLM_R_X3Y133_SLICE_X3Y133_B5Q),
.I4(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y135_SLICE_X10Y135_DO5),
.O6(CLBLM_L_X8Y135_SLICE_X10Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500d8d8d8d8)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y136_SLICE_X8Y136_CQ),
.I2(CLBLM_R_X5Y135_SLICE_X7Y135_CQ),
.I3(CLBLM_L_X12Y136_SLICE_X16Y136_A5Q),
.I4(CLBLM_L_X8Y136_SLICE_X11Y136_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y135_SLICE_X10Y135_CO5),
.O6(CLBLM_L_X8Y135_SLICE_X10Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaaaff00f0f0)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_BLUT (
.I0(CLBLM_L_X12Y136_SLICE_X16Y136_A5Q),
.I1(CLBLM_R_X7Y133_SLICE_X8Y133_BQ),
.I2(CLBLM_L_X8Y135_SLICE_X10Y135_AQ),
.I3(CLBLM_R_X7Y132_SLICE_X9Y132_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y135_SLICE_X10Y135_BO5),
.O6(CLBLM_L_X8Y135_SLICE_X10Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf5facccc0000)
  ) CLBLM_L_X8Y135_SLICE_X10Y135_ALUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_CQ),
.I1(CLBLM_L_X8Y132_SLICE_X10Y132_A5Q),
.I2(CLBLM_L_X8Y135_SLICE_X10Y135_AQ),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y135_SLICE_X9Y135_B5Q),
.O5(CLBLM_L_X8Y135_SLICE_X10Y135_AO5),
.O6(CLBLM_L_X8Y135_SLICE_X10Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y135_SLICE_X11Y135_AO6),
.Q(CLBLM_L_X8Y135_SLICE_X11Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6f6f6f6ff6f6f6f6)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_DLUT (
.I0(CLBLL_L_X4Y136_SLICE_X5Y136_AQ),
.I1(CLBLM_L_X8Y137_SLICE_X10Y137_BQ),
.I2(CLBLM_L_X10Y140_SLICE_X13Y140_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y139_SLICE_X11Y139_BQ),
.O5(CLBLM_L_X8Y135_SLICE_X11Y135_DO5),
.O6(CLBLM_L_X8Y135_SLICE_X11Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8040080420100201)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_CLUT (
.I0(CLBLM_L_X8Y132_SLICE_X10Y132_A5Q),
.I1(CLBLM_L_X8Y136_SLICE_X11Y136_AQ),
.I2(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.I3(CLBLM_L_X8Y137_SLICE_X11Y137_BQ),
.I4(CLBLM_R_X7Y136_SLICE_X9Y136_CQ),
.I5(CLBLM_L_X8Y137_SLICE_X11Y137_DQ),
.O5(CLBLM_L_X8Y135_SLICE_X11Y135_CO5),
.O6(CLBLM_L_X8Y135_SLICE_X11Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_BLUT (
.I0(CLBLM_R_X7Y136_SLICE_X9Y136_CQ),
.I1(CLBLM_L_X8Y136_SLICE_X11Y136_AQ),
.I2(CLBLL_L_X4Y136_SLICE_X5Y136_AQ),
.I3(CLBLM_L_X8Y139_SLICE_X11Y139_BQ),
.I4(CLBLM_R_X3Y136_SLICE_X3Y136_AQ),
.I5(CLBLM_L_X8Y137_SLICE_X11Y137_BQ),
.O5(CLBLM_L_X8Y135_SLICE_X11Y135_BO5),
.O6(CLBLM_L_X8Y135_SLICE_X11Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcfcfc0cfcfc0)
  ) CLBLM_L_X8Y135_SLICE_X11Y135_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y137_SLICE_X11Y137_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X3Y135_SLICE_X3Y135_A5Q),
.I4(CLBLM_R_X3Y136_SLICE_X3Y136_AQ),
.I5(CLBLM_L_X8Y134_SLICE_X11Y134_CO6),
.O5(CLBLM_L_X8Y135_SLICE_X11Y135_AO5),
.O6(CLBLM_L_X8Y135_SLICE_X11Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.Q(CLBLM_L_X8Y136_SLICE_X10Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X10Y132_SLICE_X12Y132_CQ),
.Q(CLBLM_L_X8Y136_SLICE_X10Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7dbe7dbe7dbe7dbe)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_DLUT (
.I0(CLBLM_L_X8Y136_SLICE_X11Y136_AQ),
.I1(CLBLM_L_X10Y136_SLICE_X12Y136_C5Q),
.I2(CLBLM_L_X8Y137_SLICE_X11Y137_BQ),
.I3(CLBLM_R_X7Y133_SLICE_X9Y133_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y136_SLICE_X10Y136_DO5),
.O6(CLBLM_L_X8Y136_SLICE_X10Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f000a0000000a)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_CLUT (
.I0(CLBLM_L_X8Y131_SLICE_X11Y131_CQ),
.I1(1'b1),
.I2(CLBLM_R_X11Y133_SLICE_X15Y133_AO6),
.I3(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I5(CLBLM_R_X7Y137_SLICE_X8Y137_BQ),
.O5(CLBLM_L_X8Y136_SLICE_X10Y136_CO5),
.O6(CLBLM_L_X8Y136_SLICE_X10Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1202100000000000)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_BLUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I1(CLBLM_R_X11Y132_SLICE_X15Y132_AO5),
.I2(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I3(CLBLM_R_X7Y136_SLICE_X8Y136_B5Q),
.I4(CLBLL_L_X4Y139_SLICE_X5Y139_BQ),
.I5(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.O5(CLBLM_L_X8Y136_SLICE_X10Y136_BO5),
.O6(CLBLM_L_X8Y136_SLICE_X10Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000a000a000)
  ) CLBLM_L_X8Y136_SLICE_X10Y136_ALUT (
.I0(CLBLM_R_X3Y136_SLICE_X3Y136_AQ),
.I1(CLBLM_L_X8Y137_SLICE_X11Y137_BQ),
.I2(CLBLL_L_X4Y136_SLICE_X5Y136_AQ),
.I3(CLBLM_L_X8Y139_SLICE_X11Y139_BQ),
.I4(CLBLM_L_X8Y136_SLICE_X11Y136_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y136_SLICE_X10Y136_AO5),
.O6(CLBLM_L_X8Y136_SLICE_X10Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y136_SLICE_X11Y136_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y136_SLICE_X11Y136_BO5),
.Q(CLBLM_L_X8Y136_SLICE_X11Y136_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y136_SLICE_X11Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y136_SLICE_X11Y136_AO6),
.Q(CLBLM_L_X8Y136_SLICE_X11Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y136_SLICE_X11Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y136_SLICE_X11Y136_BO6),
.Q(CLBLM_L_X8Y136_SLICE_X11Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000c0000a00ca00)
  ) CLBLM_L_X8Y136_SLICE_X11Y136_DLUT (
.I0(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.I1(CLBLM_L_X8Y135_SLICE_X10Y135_BQ),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I3(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I4(CLBLM_R_X11Y133_SLICE_X15Y133_AO6),
.I5(CLBLM_L_X12Y132_SLICE_X16Y132_BO6),
.O5(CLBLM_L_X8Y136_SLICE_X11Y136_DO5),
.O6(CLBLM_L_X8Y136_SLICE_X11Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h04050400fafffaff)
  ) CLBLM_L_X8Y136_SLICE_X11Y136_CLUT (
.I0(CLBLM_L_X12Y132_SLICE_X16Y132_BO6),
.I1(CLBLM_R_X3Y135_SLICE_X3Y135_A5Q),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I3(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I4(CLBLM_R_X7Y134_SLICE_X8Y134_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y136_SLICE_X11Y136_CO5),
.O6(CLBLM_L_X8Y136_SLICE_X11Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0dd88dd88)
  ) CLBLM_L_X8Y136_SLICE_X11Y136_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y140_SLICE_X12Y140_D5Q),
.I2(CLBLM_R_X5Y139_SLICE_X6Y139_C5Q),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_L_X8Y137_SLICE_X11Y137_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y136_SLICE_X11Y136_BO5),
.O6(CLBLM_L_X8Y136_SLICE_X11Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdefccccc12300000)
  ) CLBLM_L_X8Y136_SLICE_X11Y136_ALUT (
.I0(CLBLM_L_X8Y136_SLICE_X10Y136_AO5),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X8Y136_SLICE_X11Y136_AQ),
.I3(CLBLM_L_X8Y137_SLICE_X11Y137_BQ),
.I4(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.I5(CLBLM_L_X10Y140_SLICE_X12Y140_CQ),
.O5(CLBLM_L_X8Y136_SLICE_X11Y136_AO5),
.O6(CLBLM_L_X8Y136_SLICE_X11Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y137_SLICE_X10Y137_BO5),
.Q(CLBLM_L_X8Y137_SLICE_X10Y137_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y137_SLICE_X10Y137_CO5),
.Q(CLBLM_L_X8Y137_SLICE_X10Y137_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y137_SLICE_X10Y137_DO5),
.Q(CLBLM_L_X8Y137_SLICE_X10Y137_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y137_SLICE_X10Y137_AO6),
.Q(CLBLM_L_X8Y137_SLICE_X10Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y137_SLICE_X10Y137_BO6),
.Q(CLBLM_L_X8Y137_SLICE_X10Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y137_SLICE_X10Y137_CO6),
.Q(CLBLM_L_X8Y137_SLICE_X10Y137_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y137_SLICE_X10Y137_DO6),
.Q(CLBLM_L_X8Y137_SLICE_X10Y137_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ccccff00aaaa)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_DLUT (
.I0(CLBLM_L_X8Y132_SLICE_X10Y132_BQ),
.I1(CLBLL_L_X4Y139_SLICE_X5Y139_CQ),
.I2(CLBLM_R_X5Y126_SLICE_X6Y126_A5Q),
.I3(CLBLM_L_X10Y137_SLICE_X12Y137_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y137_SLICE_X10Y137_DO5),
.O6(CLBLM_L_X8Y137_SLICE_X10Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf055f055ccffcc00)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_CLUT (
.I0(CLBLM_R_X3Y135_SLICE_X2Y135_AQ),
.I1(CLBLM_R_X7Y137_SLICE_X8Y137_BQ),
.I2(CLBLM_R_X11Y140_SLICE_X15Y140_B5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y137_SLICE_X11Y137_D5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y137_SLICE_X10Y137_CO5),
.O6(CLBLM_L_X8Y137_SLICE_X10Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccf055f0aa)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_BLUT (
.I0(CLBLM_R_X3Y135_SLICE_X3Y135_DQ),
.I1(CLBLM_L_X10Y140_SLICE_X13Y140_BQ),
.I2(CLBLM_R_X7Y140_SLICE_X8Y140_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y132_SLICE_X9Y132_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y137_SLICE_X10Y137_BO5),
.O6(CLBLM_L_X8Y137_SLICE_X10Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeaafefe54005454)
  ) CLBLM_L_X8Y137_SLICE_X10Y137_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y135_SLICE_X10Y135_D5Q),
.I2(CLBLM_L_X8Y137_SLICE_X10Y137_AQ),
.I3(CLBLM_L_X10Y140_SLICE_X13Y140_D5Q),
.I4(CLBLM_R_X7Y131_SLICE_X9Y131_D5Q),
.I5(CLBLM_R_X5Y139_SLICE_X7Y139_CQ),
.O5(CLBLM_L_X8Y137_SLICE_X10Y137_AO5),
.O6(CLBLM_L_X8Y137_SLICE_X10Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y137_SLICE_X11Y137_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y137_SLICE_X11Y137_DO5),
.Q(CLBLM_L_X8Y137_SLICE_X11Y137_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y137_SLICE_X11Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y137_SLICE_X11Y137_AO6),
.Q(CLBLM_L_X8Y137_SLICE_X11Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y137_SLICE_X11Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y137_SLICE_X11Y137_BO6),
.Q(CLBLM_L_X8Y137_SLICE_X11Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y137_SLICE_X11Y137_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y137_SLICE_X11Y137_CO6),
.Q(CLBLM_L_X8Y137_SLICE_X11Y137_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y137_SLICE_X11Y137_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y137_SLICE_X11Y137_DO6),
.Q(CLBLM_L_X8Y137_SLICE_X11Y137_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccff0033e2e2e2e2)
  ) CLBLM_L_X8Y137_SLICE_X11Y137_DLUT (
.I0(CLBLM_R_X5Y134_SLICE_X7Y134_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y142_SLICE_X9Y142_AQ),
.I3(CLBLL_L_X4Y131_SLICE_X5Y131_B5Q),
.I4(CLBLM_R_X5Y131_SLICE_X6Y131_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y137_SLICE_X11Y137_DO5),
.O6(CLBLM_L_X8Y137_SLICE_X11Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000fc00fc)
  ) CLBLM_L_X8Y137_SLICE_X11Y137_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y137_SLICE_X11Y137_CQ),
.I2(CLBLM_R_X7Y140_SLICE_X9Y140_AQ),
.I3(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.I4(CLBLM_R_X3Y136_SLICE_X2Y136_DQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y137_SLICE_X11Y137_CO5),
.O6(CLBLM_L_X8Y137_SLICE_X11Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa3c003c00)
  ) CLBLM_L_X8Y137_SLICE_X11Y137_BLUT (
.I0(CLBLM_R_X7Y138_SLICE_X8Y138_DQ),
.I1(CLBLM_L_X8Y137_SLICE_X11Y137_BQ),
.I2(CLBLM_L_X8Y136_SLICE_X10Y136_AO5),
.I3(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y137_SLICE_X11Y137_BO5),
.O6(CLBLM_L_X8Y137_SLICE_X11Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f6f60000)
  ) CLBLM_L_X8Y137_SLICE_X11Y137_ALUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_C5Q),
.I2(CLBLM_L_X8Y137_SLICE_X11Y137_AQ),
.I3(CLBLM_L_X8Y138_SLICE_X11Y138_CQ),
.I4(CLBLM_R_X7Y135_SLICE_X9Y135_B5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y137_SLICE_X11Y137_AO5),
.O6(CLBLM_L_X8Y137_SLICE_X11Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y138_SLICE_X10Y138_AO5),
.Q(CLBLM_L_X8Y138_SLICE_X10Y138_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y138_SLICE_X10Y138_BO5),
.Q(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y138_SLICE_X10Y138_CO5),
.Q(CLBLM_L_X8Y138_SLICE_X10Y138_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y138_SLICE_X10Y138_DO5),
.Q(CLBLM_L_X8Y138_SLICE_X10Y138_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y138_SLICE_X10Y138_AO6),
.Q(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y138_SLICE_X10Y138_BO6),
.Q(CLBLM_L_X8Y138_SLICE_X10Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y138_SLICE_X10Y138_CO6),
.Q(CLBLM_L_X8Y138_SLICE_X10Y138_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y138_SLICE_X10Y138_DO6),
.Q(CLBLM_L_X8Y138_SLICE_X10Y138_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0afa0afa0)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_DLUT (
.I0(CLBLM_L_X10Y140_SLICE_X12Y140_DQ),
.I1(CLBLL_L_X4Y135_SLICE_X5Y135_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y137_SLICE_X10Y137_D5Q),
.I4(CLBLM_R_X7Y130_SLICE_X9Y130_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y138_SLICE_X10Y138_DO5),
.O6(CLBLM_L_X8Y138_SLICE_X10Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ff000afafa0a0)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_CLUT (
.I0(CLBLL_L_X4Y138_SLICE_X5Y138_C5Q),
.I1(1'b1),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y140_SLICE_X13Y140_BQ),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y138_SLICE_X10Y138_CO5),
.O6(CLBLM_L_X8Y138_SLICE_X10Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaf05058d8d8d8d)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y138_SLICE_X5Y138_D5Q),
.I2(CLBLM_L_X12Y136_SLICE_X16Y136_AQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y138_SLICE_X10Y138_BO5),
.O6(CLBLM_L_X8Y138_SLICE_X10Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888ddddaa00ff55)
  ) CLBLM_L_X8Y138_SLICE_X10Y138_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y137_SLICE_X10Y137_D5Q),
.I2(1'b1),
.I3(CLBLM_R_X7Y137_SLICE_X9Y137_BQ),
.I4(CLBLM_R_X11Y142_SLICE_X14Y142_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y138_SLICE_X10Y138_AO5),
.O6(CLBLM_L_X8Y138_SLICE_X10Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y138_SLICE_X11Y138_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y138_SLICE_X11Y138_BO5),
.Q(CLBLM_L_X8Y138_SLICE_X11Y138_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y138_SLICE_X11Y138_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y138_SLICE_X11Y138_CO5),
.Q(CLBLM_L_X8Y138_SLICE_X11Y138_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y138_SLICE_X11Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y138_SLICE_X11Y138_AO6),
.Q(CLBLM_L_X8Y138_SLICE_X11Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y138_SLICE_X11Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y138_SLICE_X11Y138_BO6),
.Q(CLBLM_L_X8Y138_SLICE_X11Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y138_SLICE_X11Y138_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y138_SLICE_X11Y138_CO6),
.Q(CLBLM_L_X8Y138_SLICE_X11Y138_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000bc8cb080)
  ) CLBLM_L_X8Y138_SLICE_X11Y138_DLUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I1(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I3(CLBLM_R_X3Y137_SLICE_X3Y137_B5Q),
.I4(CLBLM_L_X8Y138_SLICE_X11Y138_B5Q),
.I5(CLBLM_L_X10Y133_SLICE_X12Y133_CO6),
.O5(CLBLM_L_X8Y138_SLICE_X11Y138_DO5),
.O6(CLBLM_L_X8Y138_SLICE_X11Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf0aaffaa00)
  ) CLBLM_L_X8Y138_SLICE_X11Y138_CLUT (
.I0(CLBLM_L_X8Y137_SLICE_X11Y137_AQ),
.I1(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I2(CLBLM_R_X5Y137_SLICE_X7Y137_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y138_SLICE_X11Y138_CO5),
.O6(CLBLM_L_X8Y138_SLICE_X11Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888fa50fa50)
  ) CLBLM_L_X8Y138_SLICE_X11Y138_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_D5Q),
.I2(CLBLM_R_X7Y132_SLICE_X8Y132_BQ),
.I3(CLBLM_L_X8Y138_SLICE_X11Y138_BQ),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y138_SLICE_X11Y138_BO5),
.O6(CLBLM_L_X8Y138_SLICE_X11Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44af05fa50)
  ) CLBLM_L_X8Y138_SLICE_X11Y138_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_D5Q),
.I2(CLBLM_L_X8Y138_SLICE_X11Y138_AQ),
.I3(CLBLM_L_X8Y141_SLICE_X11Y141_BQ),
.I4(CLBLM_L_X8Y130_SLICE_X11Y130_AO6),
.I5(CLBLM_R_X5Y133_SLICE_X6Y133_A5Q),
.O5(CLBLM_L_X8Y138_SLICE_X11Y138_AO5),
.O6(CLBLM_L_X8Y138_SLICE_X11Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X7Y133_SLICE_X9Y133_BQ),
.Q(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1044104410001000)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_DLUT (
.I0(CLBLM_L_X10Y133_SLICE_X12Y133_CO6),
.I1(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I2(CLBLM_L_X8Y137_SLICE_X10Y137_D5Q),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I4(1'b1),
.I5(CLBLL_L_X4Y134_SLICE_X4Y134_D5Q),
.O5(CLBLM_L_X8Y139_SLICE_X10Y139_DO5),
.O6(CLBLM_L_X8Y139_SLICE_X10Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_CLUT (
.I0(CLBLM_L_X12Y134_SLICE_X17Y134_AO5),
.I1(CLBLL_L_X4Y130_SLICE_X5Y130_DO5),
.I2(CLBLM_L_X8Y139_SLICE_X11Y139_DO6),
.I3(CLBLM_R_X7Y139_SLICE_X8Y139_DO6),
.I4(CLBLM_R_X7Y139_SLICE_X9Y139_CO6),
.I5(CLBLM_L_X8Y144_SLICE_X10Y144_BO6),
.O5(CLBLM_L_X8Y139_SLICE_X10Y139_CO5),
.O6(CLBLM_L_X8Y139_SLICE_X10Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_BLUT (
.I0(CLBLM_R_X3Y133_SLICE_X3Y133_DO6),
.I1(CLBLM_L_X8Y144_SLICE_X10Y144_BO6),
.I2(CLBLM_R_X7Y134_SLICE_X8Y134_DO6),
.I3(CLBLM_R_X7Y139_SLICE_X8Y139_DO6),
.I4(CLBLM_R_X7Y139_SLICE_X8Y139_AO5),
.I5(CLBLM_L_X8Y139_SLICE_X11Y139_DO6),
.O5(CLBLM_L_X8Y139_SLICE_X10Y139_BO5),
.O6(CLBLM_L_X8Y139_SLICE_X10Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00df0020ffff0000)
  ) CLBLM_L_X8Y139_SLICE_X10Y139_ALUT (
.I0(CLBLM_L_X8Y140_SLICE_X11Y140_B5Q),
.I1(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.I2(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I3(CLBLM_L_X8Y141_SLICE_X11Y141_BQ),
.I4(CLBLM_R_X5Y137_SLICE_X7Y137_B5Q),
.I5(CLBLM_R_X7Y133_SLICE_X8Y133_A5Q),
.O5(CLBLM_L_X8Y139_SLICE_X10Y139_AO5),
.O6(CLBLM_L_X8Y139_SLICE_X10Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y139_SLICE_X11Y139_CO5),
.Q(CLBLM_L_X8Y139_SLICE_X11Y139_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y139_SLICE_X11Y139_AO6),
.Q(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y139_SLICE_X11Y139_BO6),
.Q(CLBLM_L_X8Y139_SLICE_X11Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y139_SLICE_X11Y139_CO6),
.Q(CLBLM_L_X8Y139_SLICE_X11Y139_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffefff)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_DLUT (
.I0(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.I1(CLBLM_R_X11Y141_SLICE_X14Y141_AQ),
.I2(CLBLM_L_X10Y140_SLICE_X13Y140_C5Q),
.I3(CLBLM_L_X10Y140_SLICE_X13Y140_B5Q),
.I4(CLBLL_L_X4Y133_SLICE_X4Y133_AQ),
.I5(CLBLM_L_X10Y139_SLICE_X12Y139_AO5),
.O5(CLBLM_L_X8Y139_SLICE_X11Y139_DO5),
.O6(CLBLM_L_X8Y139_SLICE_X11Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaff00ccccf0f0)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_CLUT (
.I0(CLBLM_L_X8Y138_SLICE_X11Y138_C5Q),
.I1(CLBLM_L_X8Y139_SLICE_X11Y139_CQ),
.I2(CLBLM_L_X10Y140_SLICE_X13Y140_BQ),
.I3(CLBLM_R_X5Y137_SLICE_X7Y137_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y139_SLICE_X11Y139_CO5),
.O6(CLBLM_L_X8Y139_SLICE_X11Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa33330000)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_BLUT (
.I0(CLBLM_L_X8Y140_SLICE_X11Y140_B5Q),
.I1(CLBLM_L_X8Y139_SLICE_X11Y139_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X8Y139_SLICE_X11Y139_BO5),
.O6(CLBLM_L_X8Y139_SLICE_X11Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefebaba54541010)
  ) CLBLM_L_X8Y139_SLICE_X11Y139_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X11Y131_SLICE_X14Y131_BO6),
.I2(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y140_SLICE_X6Y140_AQ),
.I5(CLBLM_L_X10Y140_SLICE_X13Y140_B5Q),
.O5(CLBLM_L_X8Y139_SLICE_X11Y139_AO5),
.O6(CLBLM_L_X8Y139_SLICE_X11Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X10Y140_CO5),
.Q(CLBLM_L_X8Y140_SLICE_X10Y140_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X10Y140_DO5),
.Q(CLBLM_L_X8Y140_SLICE_X10Y140_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X10Y140_AO6),
.Q(CLBLM_L_X8Y140_SLICE_X10Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X10Y140_BO6),
.Q(CLBLM_L_X8Y140_SLICE_X10Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X10Y140_CO6),
.Q(CLBLM_L_X8Y140_SLICE_X10Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X10Y140_DO6),
.Q(CLBLM_L_X8Y140_SLICE_X10Y140_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaaaccaacc)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_DLUT (
.I0(CLBLM_L_X10Y139_SLICE_X12Y139_AQ),
.I1(CLBLM_R_X5Y140_SLICE_X6Y140_CQ),
.I2(CLBLM_R_X5Y140_SLICE_X6Y140_A5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y140_SLICE_X10Y140_DO5),
.O6(CLBLM_L_X8Y140_SLICE_X10Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaccf0fff000)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_CLUT (
.I0(CLBLM_R_X7Y140_SLICE_X8Y140_BQ),
.I1(CLBLM_L_X8Y142_SLICE_X10Y142_A5Q),
.I2(CLBLM_L_X10Y141_SLICE_X13Y141_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(RIOB33_X105Y123_IOB_X1Y124_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y140_SLICE_X10Y140_CO5),
.O6(CLBLM_L_X8Y140_SLICE_X10Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffccf0f05544)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_BLUT (
.I0(CLBLL_L_X4Y136_SLICE_X4Y136_D5Q),
.I1(CLBLM_L_X8Y140_SLICE_X10Y140_BQ),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_AQ),
.I3(CLBLM_L_X8Y140_SLICE_X10Y140_D5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_CQ),
.O5(CLBLM_L_X8Y140_SLICE_X10Y140_BO5),
.O6(CLBLM_L_X8Y140_SLICE_X10Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbbb8b888bb88b8)
  ) CLBLM_L_X8Y140_SLICE_X10Y140_ALUT (
.I0(CLBLM_R_X5Y140_SLICE_X6Y140_CQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X8Y140_SLICE_X10Y140_AQ),
.I3(CLBLL_L_X4Y136_SLICE_X4Y136_D5Q),
.I4(CLBLM_R_X7Y140_SLICE_X8Y140_BQ),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_CQ),
.O5(CLBLM_L_X8Y140_SLICE_X10Y140_AO5),
.O6(CLBLM_L_X8Y140_SLICE_X10Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X11Y140_BO5),
.Q(CLBLM_L_X8Y140_SLICE_X11Y140_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X11Y140_AO6),
.Q(CLBLM_L_X8Y140_SLICE_X11Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X11Y140_BO6),
.Q(CLBLM_L_X8Y140_SLICE_X11Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y140_SLICE_X11Y140_CO6),
.Q(CLBLM_L_X8Y140_SLICE_X11Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffefffee)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_DLUT (
.I0(CLBLM_L_X10Y141_SLICE_X12Y141_BQ),
.I1(CLBLM_R_X7Y140_SLICE_X9Y140_D5Q),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_DO6),
.I3(CLBLM_L_X8Y134_SLICE_X11Y134_BQ),
.I4(CLBLM_L_X10Y140_SLICE_X12Y140_CQ),
.I5(CLBLM_R_X7Y136_SLICE_X8Y136_D5Q),
.O5(CLBLM_L_X8Y140_SLICE_X11Y140_DO5),
.O6(CLBLM_L_X8Y140_SLICE_X11Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe54fe54ae04ae04)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y140_SLICE_X11Y140_CQ),
.I2(CLBLM_R_X13Y134_SLICE_X18Y134_AO6),
.I3(CLBLM_L_X8Y134_SLICE_X11Y134_BQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y140_SLICE_X9Y140_CQ),
.O5(CLBLM_L_X8Y140_SLICE_X11Y140_CO5),
.O6(CLBLM_L_X8Y140_SLICE_X11Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaccffcc00)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_BLUT (
.I0(CLBLM_R_X3Y134_SLICE_X2Y134_CO6),
.I1(CLBLM_L_X10Y140_SLICE_X12Y140_BQ),
.I2(CLBLM_R_X7Y137_SLICE_X8Y137_CQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y141_SLICE_X11Y141_CO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y140_SLICE_X11Y140_BO5),
.O6(CLBLM_L_X8Y140_SLICE_X11Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haafcaaffaa30aa00)
  ) CLBLM_L_X8Y140_SLICE_X11Y140_ALUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_BQ),
.I1(CLBLM_R_X5Y133_SLICE_X7Y133_AQ),
.I2(CLBLM_L_X8Y140_SLICE_X11Y140_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y135_SLICE_X4Y135_D5Q),
.I5(CLBLM_L_X8Y139_SLICE_X11Y139_CQ),
.O5(CLBLM_L_X8Y140_SLICE_X11Y140_AO5),
.O6(CLBLM_L_X8Y140_SLICE_X11Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y141_SLICE_X10Y141_AO6),
.Q(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y141_SLICE_X10Y141_BO6),
.Q(CLBLM_L_X8Y141_SLICE_X10Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff77ffffffffffff)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_DLUT (
.I0(CLBLM_L_X10Y141_SLICE_X13Y141_CQ),
.I1(CLBLM_R_X7Y142_SLICE_X9Y142_AQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y142_SLICE_X10Y142_DO6),
.I4(CLBLM_L_X10Y141_SLICE_X13Y141_DQ),
.I5(CLBLM_L_X10Y141_SLICE_X12Y141_AQ),
.O5(CLBLM_L_X8Y141_SLICE_X10Y141_DO5),
.O6(CLBLM_L_X8Y141_SLICE_X10Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffcfcf3f3f2f3f)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_CLUT (
.I0(CLBLM_L_X8Y144_SLICE_X10Y144_AO6),
.I1(CLBLM_L_X8Y141_SLICE_X11Y141_BQ),
.I2(CLBLM_R_X7Y133_SLICE_X8Y133_A5Q),
.I3(CLBLM_L_X8Y141_SLICE_X10Y141_BQ),
.I4(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y141_SLICE_X10Y141_CO5),
.O6(CLBLM_L_X8Y141_SLICE_X10Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44aa00ef45ab01)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_BQ),
.I2(CLBLM_L_X8Y144_SLICE_X10Y144_AO6),
.I3(CLBLM_R_X5Y137_SLICE_X7Y137_A5Q),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_CO5),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_CO6),
.O5(CLBLM_L_X8Y141_SLICE_X10Y141_BO5),
.O6(CLBLM_L_X8Y141_SLICE_X10Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30cc00fd31cd01)
  ) CLBLM_L_X8Y141_SLICE_X10Y141_ALUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_BO5),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I3(CLBLM_R_X5Y134_SLICE_X7Y134_AQ),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_CO5),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_CO6),
.O5(CLBLM_L_X8Y141_SLICE_X10Y141_AO5),
.O6(CLBLM_L_X8Y141_SLICE_X10Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y141_SLICE_X11Y141_AO6),
.Q(CLBLM_L_X8Y141_SLICE_X11Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y141_SLICE_X11Y141_BO6),
.Q(CLBLM_L_X8Y141_SLICE_X11Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000022000000)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_DLUT (
.I0(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_CO6),
.I2(1'b1),
.I3(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.I4(CLBLM_L_X8Y143_SLICE_X11Y143_AQ),
.I5(CLBLM_L_X8Y143_SLICE_X10Y143_BO6),
.O5(CLBLM_L_X8Y141_SLICE_X11Y141_DO5),
.O6(CLBLM_L_X8Y141_SLICE_X11Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h30f0307833ff3333)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_CLUT (
.I0(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I1(CLBLM_R_X7Y133_SLICE_X8Y133_A5Q),
.I2(CLBLM_L_X8Y140_SLICE_X11Y140_B5Q),
.I3(CLBLM_L_X8Y141_SLICE_X11Y141_BQ),
.I4(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y141_SLICE_X11Y141_CO5),
.O6(CLBLM_L_X8Y141_SLICE_X11Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0eef0aaf0ccf000)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_BLUT (
.I0(CLBLM_L_X8Y141_SLICE_X11Y141_DO6),
.I1(CLBLM_L_X8Y141_SLICE_X11Y141_BQ),
.I2(CLBLM_R_X5Y132_SLICE_X6Y132_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y141_SLICE_X11Y141_CO5),
.I5(CLBLM_L_X10Y141_SLICE_X12Y141_CQ),
.O5(CLBLM_L_X8Y141_SLICE_X11Y141_BO5),
.O6(CLBLM_L_X8Y141_SLICE_X11Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff06000688888888)
  ) CLBLM_L_X8Y141_SLICE_X11Y141_ALUT (
.I0(CLBLM_L_X8Y141_SLICE_X11Y141_AQ),
.I1(CLBLM_L_X10Y134_SLICE_X12Y134_AQ),
.I2(CLBLM_R_X5Y140_SLICE_X7Y140_A5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X11Y140_SLICE_X14Y140_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y141_SLICE_X11Y141_AO5),
.O6(CLBLM_L_X8Y141_SLICE_X11Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X10Y142_BO6),
.Q(CLBLM_L_X8Y142_SLICE_X10Y142_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X10Y142_AO6),
.Q(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff7fffffffffff)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_DLUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I1(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.I2(CLBLM_R_X7Y142_SLICE_X9Y142_CQ),
.I3(CLBLM_R_X7Y142_SLICE_X9Y142_BQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y141_SLICE_X11Y141_AQ),
.O5(CLBLM_L_X8Y142_SLICE_X10Y142_DO5),
.O6(CLBLM_L_X8Y142_SLICE_X10Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h80000000c0000000)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_CLUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I1(CLBLM_L_X10Y134_SLICE_X12Y134_AQ),
.I2(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.I3(CLBLM_L_X8Y141_SLICE_X11Y141_AQ),
.I4(CLBLM_R_X7Y142_SLICE_X9Y142_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y142_SLICE_X10Y142_CO5),
.O6(CLBLM_L_X8Y142_SLICE_X10Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00ffcc00cc00)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_BLUT (
.I0(CLBLM_L_X8Y134_SLICE_X10Y134_A5Q),
.I1(CLBLM_L_X8Y141_SLICE_X11Y141_BQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y133_SLICE_X8Y133_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y142_SLICE_X10Y142_BO5),
.O6(CLBLM_L_X8Y142_SLICE_X10Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff007800000078)
  ) CLBLM_L_X8Y142_SLICE_X10Y142_ALUT (
.I0(CLBLM_R_X7Y142_SLICE_X9Y142_CQ),
.I1(CLBLM_L_X8Y141_SLICE_X11Y141_AO5),
.I2(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.I3(CLBLM_R_X5Y140_SLICE_X7Y140_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X10Y141_SLICE_X12Y141_C5Q),
.O5(CLBLM_L_X8Y142_SLICE_X10Y142_AO5),
.O6(CLBLM_L_X8Y142_SLICE_X10Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X11Y142_AO6),
.Q(CLBLM_L_X8Y142_SLICE_X11Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y142_SLICE_X11Y142_BO6),
.Q(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0080000000000000)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_DLUT (
.I0(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.I1(CLBLM_L_X8Y143_SLICE_X11Y143_AQ),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_BO5),
.I4(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I5(CLBLM_R_X7Y143_SLICE_X8Y143_A5Q),
.O5(CLBLM_L_X8Y142_SLICE_X11Y142_DO5),
.O6(CLBLM_L_X8Y142_SLICE_X11Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5fffff7f7fffff)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_CLUT (
.I0(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I1(CLBLM_L_X8Y142_SLICE_X11Y142_AQ),
.I2(CLBLM_L_X8Y140_SLICE_X11Y140_B5Q),
.I3(1'b1),
.I4(CLBLM_R_X5Y137_SLICE_X7Y137_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y142_SLICE_X11Y142_CO5),
.O6(CLBLM_L_X8Y142_SLICE_X11Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff008888ff00b8b8)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_BLUT (
.I0(CLBLM_L_X8Y143_SLICE_X11Y143_BO6),
.I1(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.I2(CLBLM_L_X8Y143_SLICE_X11Y143_AQ),
.I3(CLBLM_L_X10Y135_SLICE_X12Y135_B5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X8Y143_SLICE_X11Y143_CO6),
.O5(CLBLM_L_X8Y142_SLICE_X11Y142_BO5),
.O6(CLBLM_L_X8Y142_SLICE_X11Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb888b888b888b8bb)
  ) CLBLM_L_X8Y142_SLICE_X11Y142_ALUT (
.I0(CLBLM_L_X8Y138_SLICE_X11Y138_B5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_DO6),
.I3(CLBLM_L_X8Y142_SLICE_X11Y142_AQ),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_CO6),
.I5(CLBLM_L_X8Y142_SLICE_X11Y142_CO6),
.O5(CLBLM_L_X8Y142_SLICE_X11Y142_AO5),
.O6(CLBLM_L_X8Y142_SLICE_X11Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X10Y143_AO6),
.Q(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff007f00ff)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_DLUT (
.I0(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I1(CLBLM_R_X5Y137_SLICE_X7Y137_B5Q),
.I2(CLBLM_L_X8Y140_SLICE_X11Y140_B5Q),
.I3(CLBLM_L_X8Y142_SLICE_X10Y142_BO5),
.I4(CLBLM_L_X8Y142_SLICE_X11Y142_AQ),
.I5(CLBLM_R_X7Y143_SLICE_X9Y143_BO5),
.O5(CLBLM_L_X8Y143_SLICE_X10Y143_DO5),
.O6(CLBLM_L_X8Y143_SLICE_X10Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffff7ffff)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_CLUT (
.I0(CLBLM_R_X7Y133_SLICE_X8Y133_A5Q),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I2(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.I3(CLBLM_L_X8Y144_SLICE_X10Y144_AO6),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_BQ),
.I5(CLBLM_L_X8Y141_SLICE_X11Y141_BQ),
.O5(CLBLM_L_X8Y143_SLICE_X10Y143_CO5),
.O6(CLBLM_L_X8Y143_SLICE_X10Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff7fffffff33ff33)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_BLUT (
.I0(CLBLM_R_X7Y143_SLICE_X8Y143_A5Q),
.I1(CLBLM_L_X8Y141_SLICE_X10Y141_BQ),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I3(CLBLM_L_X8Y144_SLICE_X10Y144_AO6),
.I4(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y143_SLICE_X10Y143_BO5),
.O6(CLBLM_L_X8Y143_SLICE_X10Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaffaa3caa3c)
  ) CLBLM_L_X8Y143_SLICE_X10Y143_ALUT (
.I0(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I1(CLBLM_L_X8Y142_SLICE_X10Y142_CO5),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(CLBLM_R_X5Y140_SLICE_X7Y140_A5Q),
.O5(CLBLM_L_X8Y143_SLICE_X10Y143_AO5),
.O6(CLBLM_L_X8Y143_SLICE_X10Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y143_SLICE_X11Y143_AO6),
.Q(CLBLM_L_X8Y143_SLICE_X11Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y143_SLICE_X11Y143_DO5),
.O6(CLBLM_L_X8Y143_SLICE_X11Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff7ffffffffffff)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_CLUT (
.I0(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.I1(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I2(CLBLM_L_X8Y143_SLICE_X10Y143_BO5),
.I3(CLBLM_L_X8Y141_SLICE_X10Y141_CO6),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I5(CLBLM_R_X7Y143_SLICE_X8Y143_A5Q),
.O5(CLBLM_L_X8Y143_SLICE_X11Y143_CO5),
.O6(CLBLM_L_X8Y143_SLICE_X11Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ef00ffffffffff)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_BLUT (
.I0(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.I1(CLBLM_L_X8Y143_SLICE_X10Y143_BO6),
.I2(CLBLM_L_X8Y143_SLICE_X11Y143_AQ),
.I3(CLBLM_L_X8Y141_SLICE_X11Y141_BQ),
.I4(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.I5(CLBLM_R_X7Y133_SLICE_X8Y133_A5Q),
.O5(CLBLM_L_X8Y143_SLICE_X11Y143_BO5),
.O6(CLBLM_L_X8Y143_SLICE_X11Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfccc3000ffcf3303)
  ) CLBLM_L_X8Y143_SLICE_X11Y143_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X8Y143_SLICE_X11Y143_AQ),
.I3(CLBLM_L_X8Y143_SLICE_X11Y143_BO6),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_AQ),
.I5(CLBLM_L_X8Y143_SLICE_X11Y143_CO6),
.O5(CLBLM_L_X8Y143_SLICE_X11Y143_AO5),
.O6(CLBLM_L_X8Y143_SLICE_X11Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y144_SLICE_X10Y144_DO5),
.O6(CLBLM_L_X8Y144_SLICE_X10Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y144_SLICE_X10Y144_CO5),
.O6(CLBLM_L_X8Y144_SLICE_X10Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffff7fff)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_BLUT (
.I0(CLBLM_R_X5Y137_SLICE_X7Y137_B5Q),
.I1(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I2(CLBLM_L_X8Y142_SLICE_X11Y142_AQ),
.I3(CLBLM_L_X8Y140_SLICE_X11Y140_B5Q),
.I4(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_CO6),
.O5(CLBLM_L_X8Y144_SLICE_X10Y144_BO5),
.O6(CLBLM_L_X8Y144_SLICE_X10Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffffffffffff)
  ) CLBLM_L_X8Y144_SLICE_X10Y144_ALUT (
.I0(CLBLM_R_X5Y137_SLICE_X7Y137_B5Q),
.I1(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I2(CLBLM_L_X8Y142_SLICE_X11Y142_AQ),
.I3(CLBLM_L_X8Y140_SLICE_X11Y140_B5Q),
.I4(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I5(CLBLM_L_X10Y141_SLICE_X12Y141_C5Q),
.O5(CLBLM_L_X8Y144_SLICE_X10Y144_AO5),
.O6(CLBLM_L_X8Y144_SLICE_X10Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y144_SLICE_X11Y144_DO5),
.O6(CLBLM_L_X8Y144_SLICE_X11Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y144_SLICE_X11Y144_CO5),
.O6(CLBLM_L_X8Y144_SLICE_X11Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y144_SLICE_X11Y144_BO5),
.O6(CLBLM_L_X8Y144_SLICE_X11Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y144_SLICE_X11Y144_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y144_SLICE_X11Y144_AO5),
.O6(CLBLM_L_X8Y144_SLICE_X11Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y130_SLICE_X12Y130_BO5),
.Q(CLBLM_L_X10Y130_SLICE_X12Y130_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y130_SLICE_X12Y130_CO5),
.Q(CLBLM_L_X10Y130_SLICE_X12Y130_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y130_SLICE_X12Y130_AO6),
.Q(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y130_SLICE_X12Y130_BO6),
.Q(CLBLM_L_X10Y130_SLICE_X12Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y130_SLICE_X12Y130_CO6),
.Q(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_DO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfc0cacacacac)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_CLUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_AQ),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_CO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0f0ccccff00)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_BLUT (
.I0(CLBLM_L_X10Y135_SLICE_X12Y135_A5Q),
.I1(CLBLM_L_X10Y130_SLICE_X12Y130_BQ),
.I2(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.I3(RIOB33_X105Y127_IOB_X1Y128_I),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_BO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccca0aaaaa0)
  ) CLBLM_L_X10Y130_SLICE_X12Y130_ALUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_B5Q),
.I1(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I2(CLBLM_L_X10Y130_SLICE_X12Y130_AQ),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(CLBLM_L_X10Y130_SLICE_X12Y130_C5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X10Y130_SLICE_X12Y130_AO5),
.O6(CLBLM_L_X10Y130_SLICE_X12Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_DO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_CO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_BO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y130_SLICE_X13Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y130_SLICE_X13Y130_AO5),
.O6(CLBLM_L_X10Y130_SLICE_X13Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X12Y131_CO5),
.Q(CLBLM_L_X10Y131_SLICE_X12Y131_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X12Y131_DO5),
.Q(CLBLM_L_X10Y131_SLICE_X12Y131_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X12Y131_AO6),
.Q(CLBLM_L_X10Y131_SLICE_X12Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X12Y131_BO6),
.Q(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X12Y131_CO6),
.Q(CLBLM_L_X10Y131_SLICE_X12Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X12Y131_DO6),
.Q(CLBLM_L_X10Y131_SLICE_X12Y131_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ff000acacacac)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_DLUT (
.I0(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y131_SLICE_X11Y131_D5Q),
.I4(CLBLL_L_X4Y136_SLICE_X4Y136_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_DO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0f0ccccff00)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_CLUT (
.I0(CLBLM_L_X10Y132_SLICE_X12Y132_C5Q),
.I1(CLBLM_L_X10Y131_SLICE_X12Y131_CQ),
.I2(CLBLM_R_X3Y135_SLICE_X3Y135_DQ),
.I3(CLBLM_R_X3Y137_SLICE_X3Y137_B5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_CO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000fffc00fc)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.I2(CLBLL_L_X4Y131_SLICE_X5Y131_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y131_SLICE_X12Y131_C5Q),
.I5(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_BO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88d8d8dd88)
  ) CLBLM_L_X10Y131_SLICE_X12Y131_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y131_SLICE_X11Y131_BQ),
.I2(CLBLM_L_X10Y131_SLICE_X12Y131_AQ),
.I3(CLBLM_L_X10Y131_SLICE_X12Y131_CQ),
.I4(CLBLM_R_X7Y131_SLICE_X9Y131_D5Q),
.I5(CLBLM_L_X10Y140_SLICE_X13Y140_D5Q),
.O5(CLBLM_L_X10Y131_SLICE_X12Y131_AO5),
.O6(CLBLM_L_X10Y131_SLICE_X12Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X13Y131_AO6),
.Q(CLBLM_L_X10Y131_SLICE_X13Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y131_SLICE_X13Y131_BO6),
.Q(CLBLM_L_X10Y131_SLICE_X13Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5d0c5d0cffff5d0c)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_DLUT (
.I0(CLBLM_R_X11Y131_SLICE_X14Y131_AO6),
.I1(CLBLM_R_X5Y126_SLICE_X6Y126_A5Q),
.I2(CLBLM_R_X11Y132_SLICE_X15Y132_BO6),
.I3(CLBLM_L_X8Y139_SLICE_X11Y139_C5Q),
.I4(CLBLM_R_X7Y131_SLICE_X8Y131_CQ),
.I5(CLBLM_R_X11Y131_SLICE_X14Y131_AO5),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_DO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f773f335f550f00)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_CLUT (
.I0(CLBLM_R_X11Y131_SLICE_X14Y131_AO6),
.I1(CLBLM_R_X11Y131_SLICE_X14Y131_AO5),
.I2(CLBLM_R_X11Y132_SLICE_X15Y132_BO6),
.I3(CLBLL_L_X4Y130_SLICE_X5Y130_B5Q),
.I4(CLBLM_R_X7Y134_SLICE_X8Y134_AQ),
.I5(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_CO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd8ddd8ddd8d8888)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y132_SLICE_X13Y132_AQ),
.I2(CLBLL_L_X4Y135_SLICE_X5Y135_CQ),
.I3(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I4(CLBLM_L_X10Y131_SLICE_X13Y131_BQ),
.I5(CLBLM_R_X7Y131_SLICE_X9Y131_DQ),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_BO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88d8d8dd88dd88)
  ) CLBLM_L_X10Y131_SLICE_X13Y131_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y131_SLICE_X13Y131_BQ),
.I2(CLBLM_L_X10Y131_SLICE_X13Y131_AQ),
.I3(CLBLM_L_X8Y131_SLICE_X11Y131_D5Q),
.I4(CLBLM_R_X5Y133_SLICE_X7Y133_AQ),
.I5(CLBLL_L_X4Y135_SLICE_X4Y135_D5Q),
.O5(CLBLM_L_X10Y131_SLICE_X13Y131_AO5),
.O6(CLBLM_L_X10Y131_SLICE_X13Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y132_SLICE_X12Y132_CO5),
.Q(CLBLM_L_X10Y132_SLICE_X12Y132_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y132_SLICE_X12Y132_AO6),
.Q(CLBLM_L_X10Y132_SLICE_X12Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y132_SLICE_X12Y132_BO6),
.Q(CLBLM_L_X10Y132_SLICE_X12Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y132_SLICE_X12Y132_CO6),
.Q(CLBLM_L_X10Y132_SLICE_X12Y132_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0010000000000000)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_DLUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I1(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I2(CLBLM_R_X7Y132_SLICE_X9Y132_CQ),
.I3(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I4(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I5(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_DO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ff000cfc0cfc0)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y135_SLICE_X2Y135_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y131_SLICE_X12Y131_DQ),
.I4(CLBLM_L_X8Y131_SLICE_X11Y131_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_CO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hefeaefea45404540)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y132_SLICE_X12Y132_BQ),
.I2(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.I3(CLBLM_R_X5Y130_SLICE_X7Y130_AQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_BO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbeaa1400eeaa4400)
  ) CLBLM_L_X10Y132_SLICE_X12Y132_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y132_SLICE_X12Y132_AQ),
.I2(CLBLM_L_X8Y132_SLICE_X11Y132_AQ),
.I3(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.I4(CLBLM_L_X10Y131_SLICE_X12Y131_AQ),
.I5(CLBLM_L_X8Y135_SLICE_X11Y135_BO6),
.O5(CLBLM_L_X10Y132_SLICE_X12Y132_AO5),
.O6(CLBLM_L_X10Y132_SLICE_X12Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y132_SLICE_X13Y132_AO6),
.Q(CLBLM_L_X10Y132_SLICE_X13Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5040504000400040)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_DLUT (
.I0(CLBLM_R_X11Y131_SLICE_X15Y131_AO6),
.I1(CLBLM_L_X8Y139_SLICE_X11Y139_C5Q),
.I2(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I4(1'b1),
.I5(CLBLM_R_X7Y131_SLICE_X8Y131_CQ),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_DO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4000400070304000)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_CLUT (
.I0(CLBLM_L_X12Y132_SLICE_X16Y132_BO6),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I2(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I3(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.I4(CLBLM_L_X8Y134_SLICE_X10Y134_AQ),
.I5(CLBLM_R_X11Y131_SLICE_X15Y131_AO6),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_CO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a0a0a0a0ace0a)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_BLUT (
.I0(CLBLM_L_X8Y132_SLICE_X10Y132_B5Q),
.I1(CLBLL_L_X4Y132_SLICE_X5Y132_DQ),
.I2(CLBLM_R_X11Y131_SLICE_X14Y131_AO6),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I4(CLBLM_L_X12Y132_SLICE_X16Y132_BO6),
.I5(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_BO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0ffcc00f000cc)
  ) CLBLM_L_X10Y132_SLICE_X13Y132_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y134_SLICE_X5Y134_BQ),
.I2(CLBLM_L_X10Y132_SLICE_X13Y132_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X12Y132_SLICE_X16Y132_AO6),
.I5(CLBLL_L_X4Y134_SLICE_X4Y134_C5Q),
.O5(CLBLM_L_X10Y132_SLICE_X13Y132_AO5),
.O6(CLBLM_L_X10Y132_SLICE_X13Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y133_SLICE_X12Y133_AO5),
.Q(CLBLM_L_X10Y133_SLICE_X12Y133_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y133_SLICE_X12Y133_AO6),
.Q(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y133_SLICE_X12Y133_BO6),
.Q(CLBLM_L_X10Y133_SLICE_X12Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000e000e00040004)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_DLUT (
.I0(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I1(CLBLM_R_X7Y135_SLICE_X8Y135_AQ),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I3(CLBLM_L_X10Y133_SLICE_X12Y133_CO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y130_SLICE_X12Y130_BQ),
.O5(CLBLM_L_X10Y133_SLICE_X12Y133_DO5),
.O6(CLBLM_L_X10Y133_SLICE_X12Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_CLUT (
.I0(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.I1(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I2(CLBLM_R_X7Y137_SLICE_X8Y137_CQ),
.I3(CLBLL_L_X4Y136_SLICE_X5Y136_D5Q),
.I4(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I5(CLBLM_L_X8Y134_SLICE_X10Y134_A5Q),
.O5(CLBLM_L_X10Y133_SLICE_X12Y133_CO5),
.O6(CLBLM_L_X10Y133_SLICE_X12Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffe4ffe400e400e4)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_BLUT (
.I0(CLBLM_R_X13Y134_SLICE_X18Y134_AO6),
.I1(CLBLM_L_X10Y133_SLICE_X12Y133_BQ),
.I2(CLBLM_L_X10Y131_SLICE_X13Y131_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y134_SLICE_X11Y134_B5Q),
.O5(CLBLM_L_X10Y133_SLICE_X12Y133_BO5),
.O6(CLBLM_L_X10Y133_SLICE_X12Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000ccaaccaa)
  ) CLBLM_L_X10Y133_SLICE_X12Y133_ALUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(CLBLM_L_X8Y133_SLICE_X10Y133_CQ),
.I2(CLBLM_R_X3Y131_SLICE_X2Y131_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X11Y141_SLICE_X14Y141_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y133_SLICE_X12Y133_AO5),
.O6(CLBLM_L_X10Y133_SLICE_X12Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y133_SLICE_X13Y133_AO6),
.Q(CLBLM_L_X10Y133_SLICE_X13Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff50ff50ffdcffdc)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_DLUT (
.I0(CLBLM_R_X11Y131_SLICE_X14Y131_AO6),
.I1(CLBLM_R_X7Y137_SLICE_X8Y137_B5Q),
.I2(CLBLL_L_X4Y134_SLICE_X4Y134_A5Q),
.I3(CLBLM_L_X10Y133_SLICE_X13Y133_CO6),
.I4(1'b1),
.I5(CLBLM_R_X11Y134_SLICE_X14Y134_AO6),
.O5(CLBLM_L_X10Y133_SLICE_X13Y133_DO5),
.O6(CLBLM_L_X10Y133_SLICE_X13Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0022f0f20022f0f2)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_CLUT (
.I0(CLBLL_L_X4Y131_SLICE_X5Y131_B5Q),
.I1(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I2(CLBLM_R_X5Y134_SLICE_X6Y134_B5Q),
.I3(CLBLM_L_X12Y136_SLICE_X17Y136_BO6),
.I4(CLBLM_R_X11Y132_SLICE_X15Y132_BO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y133_SLICE_X13Y133_CO5),
.O6(CLBLM_L_X10Y133_SLICE_X13Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0cff0cff5dff0c)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_BLUT (
.I0(CLBLM_L_X12Y136_SLICE_X17Y136_BO6),
.I1(CLBLM_R_X7Y133_SLICE_X9Y133_DQ),
.I2(CLBLM_R_X11Y132_SLICE_X15Y132_BO6),
.I3(CLBLM_L_X10Y132_SLICE_X13Y132_CO6),
.I4(CLBLM_R_X11Y141_SLICE_X14Y141_AQ),
.I5(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.O5(CLBLM_L_X10Y133_SLICE_X13Y133_BO5),
.O6(CLBLM_L_X10Y133_SLICE_X13Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccffcca0ccf0)
  ) CLBLM_L_X10Y133_SLICE_X13Y133_ALUT (
.I0(CLBLM_R_X5Y133_SLICE_X7Y133_AQ),
.I1(CLBLM_R_X7Y133_SLICE_X8Y133_A5Q),
.I2(CLBLM_L_X10Y133_SLICE_X13Y133_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y135_SLICE_X4Y135_D5Q),
.I5(CLBLM_L_X8Y133_SLICE_X11Y133_B5Q),
.O5(CLBLM_L_X10Y133_SLICE_X13Y133_AO5),
.O6(CLBLM_L_X10Y133_SLICE_X13Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y134_SLICE_X12Y134_AO5),
.Q(CLBLM_L_X10Y134_SLICE_X12Y134_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y134_SLICE_X12Y134_BO5),
.Q(CLBLM_L_X10Y134_SLICE_X12Y134_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y134_SLICE_X12Y134_AO6),
.Q(CLBLM_L_X10Y134_SLICE_X12Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y134_SLICE_X12Y134_BO6),
.Q(CLBLM_L_X10Y134_SLICE_X12Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7b7b7b7bdededede)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_DLUT (
.I0(CLBLM_L_X10Y132_SLICE_X12Y132_AQ),
.I1(CLBLM_L_X10Y134_SLICE_X13Y134_A5Q),
.I2(CLBLM_L_X10Y134_SLICE_X12Y134_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y132_SLICE_X11Y132_BQ),
.O5(CLBLM_L_X10Y134_SLICE_X12Y134_DO5),
.O6(CLBLM_L_X10Y134_SLICE_X12Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000551100004400)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_CLUT (
.I0(CLBLM_R_X11Y133_SLICE_X15Y133_AO6),
.I1(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I2(1'b1),
.I3(CLBLM_L_X10Y135_SLICE_X13Y135_AQ),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I5(CLBLM_R_X7Y133_SLICE_X9Y133_AQ),
.O5(CLBLM_L_X10Y134_SLICE_X12Y134_CO5),
.O6(CLBLM_L_X10Y134_SLICE_X12Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccffaa00aa)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_BLUT (
.I0(CLBLL_L_X4Y137_SLICE_X5Y137_A5Q),
.I1(CLBLM_R_X11Y141_SLICE_X14Y141_AQ),
.I2(CLBLM_L_X8Y134_SLICE_X11Y134_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y139_SLICE_X13Y139_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y134_SLICE_X12Y134_BO5),
.O6(CLBLM_L_X10Y134_SLICE_X12Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaf0ccffcc00)
  ) CLBLM_L_X10Y134_SLICE_X12Y134_ALUT (
.I0(CLBLM_R_X7Y139_SLICE_X9Y139_AQ),
.I1(CLBLM_L_X8Y132_SLICE_X11Y132_AQ),
.I2(CLBLM_L_X10Y132_SLICE_X12Y132_C5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y135_SLICE_X10Y135_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y134_SLICE_X12Y134_AO5),
.O6(CLBLM_L_X10Y134_SLICE_X12Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y134_SLICE_X13Y134_AO5),
.Q(CLBLM_L_X10Y134_SLICE_X13Y134_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y134_SLICE_X13Y134_AO6),
.Q(CLBLM_L_X10Y134_SLICE_X13Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff0faf0faf0fa)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_DLUT (
.I0(CLBLM_L_X10Y139_SLICE_X13Y139_AQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y133_SLICE_X12Y133_DO6),
.I3(CLBLM_R_X11Y136_SLICE_X15Y136_AO5),
.I4(CLBLM_R_X7Y134_SLICE_X9Y134_CQ),
.I5(CLBLM_L_X12Y132_SLICE_X16Y132_AO6),
.O5(CLBLM_L_X10Y134_SLICE_X13Y134_DO5),
.O6(CLBLM_L_X10Y134_SLICE_X13Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h30baffff30ba30ba)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_CLUT (
.I0(CLBLM_R_X5Y131_SLICE_X6Y131_AQ),
.I1(CLBLM_L_X12Y134_SLICE_X16Y134_AO6),
.I2(CLBLL_L_X4Y136_SLICE_X5Y136_DQ),
.I3(CLBLM_R_X11Y136_SLICE_X15Y136_AO5),
.I4(CLBLM_L_X12Y134_SLICE_X16Y134_AO5),
.I5(CLBLM_L_X8Y136_SLICE_X11Y136_BQ),
.O5(CLBLM_L_X10Y134_SLICE_X13Y134_CO5),
.O6(CLBLM_L_X10Y134_SLICE_X13Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2200000022000030)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_BLUT (
.I0(CLBLM_R_X7Y139_SLICE_X9Y139_AQ),
.I1(CLBLM_R_X11Y136_SLICE_X14Y136_CO6),
.I2(CLBLM_L_X8Y133_SLICE_X10Y133_AQ),
.I3(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I5(CLBLM_R_X11Y140_SLICE_X14Y140_BO6),
.O5(CLBLM_L_X10Y134_SLICE_X13Y134_BO5),
.O6(CLBLM_L_X10Y134_SLICE_X13Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aaffcc00ccff)
  ) CLBLM_L_X10Y134_SLICE_X13Y134_ALUT (
.I0(CLBLM_L_X10Y136_SLICE_X13Y136_AQ),
.I1(CLBLM_L_X8Y136_SLICE_X11Y136_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y140_SLICE_X13Y140_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y134_SLICE_X13Y134_AO5),
.O6(CLBLM_L_X10Y134_SLICE_X13Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y135_SLICE_X12Y135_AO5),
.Q(CLBLM_L_X10Y135_SLICE_X12Y135_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y135_SLICE_X12Y135_BO5),
.Q(CLBLM_L_X10Y135_SLICE_X12Y135_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y135_SLICE_X12Y135_AO6),
.Q(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y135_SLICE_X12Y135_BO6),
.Q(CLBLM_L_X10Y135_SLICE_X12Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0202000002020f00)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_DLUT (
.I0(CLBLM_R_X7Y139_SLICE_X9Y139_BQ),
.I1(CLBLM_R_X11Y136_SLICE_X14Y136_CO6),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I3(CLBLM_L_X10Y137_SLICE_X12Y137_AQ),
.I4(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I5(CLBLM_L_X10Y133_SLICE_X12Y133_CO6),
.O5(CLBLM_L_X10Y135_SLICE_X12Y135_DO5),
.O6(CLBLM_L_X10Y135_SLICE_X12Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8f888f88ffff8f88)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_CLUT (
.I0(CLBLM_L_X12Y132_SLICE_X16Y132_AO6),
.I1(CLBLM_R_X3Y135_SLICE_X2Y135_CQ),
.I2(CLBLM_L_X12Y135_SLICE_X16Y135_AO5),
.I3(CLBLM_L_X10Y132_SLICE_X12Y132_CQ),
.I4(CLBLM_L_X10Y135_SLICE_X12Y135_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y135_SLICE_X12Y135_CO5),
.O6(CLBLM_L_X10Y135_SLICE_X12Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacacacfc0cfc0c)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_BLUT (
.I0(CLBLM_R_X7Y135_SLICE_X8Y135_AQ),
.I1(CLBLM_L_X12Y136_SLICE_X16Y136_A5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y140_SLICE_X8Y140_D5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y135_SLICE_X12Y135_BO5),
.O6(CLBLM_L_X10Y135_SLICE_X12Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f0f0ccccaaaa)
  ) CLBLM_L_X10Y135_SLICE_X12Y135_ALUT (
.I0(CLBLM_L_X10Y135_SLICE_X12Y135_B5Q),
.I1(CLBLM_L_X10Y138_SLICE_X13Y138_CQ),
.I2(CLBLL_L_X4Y134_SLICE_X4Y134_C5Q),
.I3(CLBLM_L_X8Y135_SLICE_X10Y135_D5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y135_SLICE_X12Y135_AO5),
.O6(CLBLM_L_X10Y135_SLICE_X12Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y136_SLICE_X13Y136_CO5),
.Q(CLBLM_L_X10Y135_SLICE_X13Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff0a0acece)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_DLUT (
.I0(CLBLM_L_X8Y140_SLICE_X11Y140_AQ),
.I1(CLBLM_R_X5Y135_SLICE_X7Y135_B5Q),
.I2(CLBLM_R_X11Y131_SLICE_X14Y131_BO6),
.I3(1'b1),
.I4(CLBLM_L_X12Y134_SLICE_X17Y134_AO5),
.I5(CLBLM_R_X11Y140_SLICE_X14Y140_BO6),
.O5(CLBLM_L_X10Y135_SLICE_X13Y135_DO5),
.O6(CLBLM_L_X10Y135_SLICE_X13Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55f500f0ddfdccfc)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_CLUT (
.I0(CLBLM_L_X12Y134_SLICE_X16Y134_AO6),
.I1(CLBLM_R_X5Y135_SLICE_X7Y135_AQ),
.I2(CLBLM_R_X5Y136_SLICE_X6Y136_CQ),
.I3(CLBLM_L_X12Y136_SLICE_X17Y136_AO6),
.I4(CLBLM_R_X3Y134_SLICE_X3Y134_A5Q),
.I5(CLBLM_R_X11Y136_SLICE_X15Y136_AO5),
.O5(CLBLM_L_X10Y135_SLICE_X13Y135_CO5),
.O6(CLBLM_L_X10Y135_SLICE_X13Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaffeefffafffe)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_BLUT (
.I0(CLBLM_L_X10Y135_SLICE_X13Y135_DO6),
.I1(CLBLM_L_X10Y137_SLICE_X12Y137_AQ),
.I2(CLBLM_R_X7Y139_SLICE_X9Y139_BQ),
.I3(CLBLM_L_X10Y135_SLICE_X12Y135_CO6),
.I4(CLBLM_R_X11Y136_SLICE_X15Y136_AO6),
.I5(CLBLM_L_X12Y136_SLICE_X17Y136_AO6),
.O5(CLBLM_L_X10Y135_SLICE_X13Y135_BO5),
.O6(CLBLM_L_X10Y135_SLICE_X13Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcfcfcfffefefe)
  ) CLBLM_L_X10Y135_SLICE_X13Y135_ALUT (
.I0(CLBLM_R_X7Y137_SLICE_X9Y137_BQ),
.I1(CLBLM_R_X11Y140_SLICE_X14Y140_BO6),
.I2(CLBLM_L_X8Y133_SLICE_X11Y133_CO6),
.I3(CLBLM_L_X10Y138_SLICE_X13Y138_CQ),
.I4(CLBLM_R_X11Y133_SLICE_X14Y133_CO6),
.I5(CLBLM_L_X12Y136_SLICE_X17Y136_AO6),
.O5(CLBLM_L_X10Y135_SLICE_X13Y135_AO5),
.O6(CLBLM_L_X10Y135_SLICE_X13Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y136_SLICE_X12Y136_CO5),
.Q(CLBLM_L_X10Y136_SLICE_X12Y136_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y136_SLICE_X12Y136_AO6),
.Q(CLBLM_L_X10Y136_SLICE_X12Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y136_SLICE_X12Y136_BO6),
.Q(CLBLM_L_X10Y136_SLICE_X12Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y136_SLICE_X12Y136_CO6),
.Q(CLBLM_L_X10Y136_SLICE_X12Y136_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_DLUT (
.I0(CLBLM_L_X10Y139_SLICE_X12Y139_CO6),
.I1(CLBLM_L_X10Y132_SLICE_X12Y132_DO6),
.I2(CLBLM_L_X8Y136_SLICE_X11Y136_DO6),
.I3(CLBLM_L_X10Y137_SLICE_X12Y137_AO5),
.I4(CLBLM_L_X10Y139_SLICE_X12Y139_DO6),
.I5(CLBLM_L_X8Y136_SLICE_X10Y136_BO6),
.O5(CLBLM_L_X10Y136_SLICE_X12Y136_DO5),
.O6(CLBLM_L_X10Y136_SLICE_X12Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500f5a0f5a0)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(CLBLM_L_X10Y131_SLICE_X13Y131_AQ),
.I3(CLBLM_L_X12Y136_SLICE_X16Y136_AQ),
.I4(CLBLM_R_X5Y132_SLICE_X7Y132_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y136_SLICE_X12Y136_CO5),
.O6(CLBLM_L_X10Y136_SLICE_X12Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aafff0f088cc)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_BLUT (
.I0(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I1(CLBLM_L_X10Y136_SLICE_X12Y136_BQ),
.I2(CLBLM_L_X10Y136_SLICE_X12Y136_AQ),
.I3(CLBLL_L_X4Y135_SLICE_X5Y135_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y136_SLICE_X9Y136_DQ),
.O5(CLBLM_L_X10Y136_SLICE_X12Y136_BO5),
.O6(CLBLM_L_X10Y136_SLICE_X12Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafff0aaaa3330)
  ) CLBLM_L_X10Y136_SLICE_X12Y136_ALUT (
.I0(CLBLM_L_X10Y140_SLICE_X13Y140_CQ),
.I1(CLBLL_L_X4Y135_SLICE_X5Y135_CQ),
.I2(CLBLM_L_X10Y136_SLICE_X12Y136_AQ),
.I3(CLBLM_L_X8Y133_SLICE_X10Y133_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.O5(CLBLM_L_X10Y136_SLICE_X12Y136_AO5),
.O6(CLBLM_L_X10Y136_SLICE_X12Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y136_SLICE_X13Y136_AO6),
.Q(CLBLM_L_X10Y136_SLICE_X13Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y136_SLICE_X13Y136_BO6),
.Q(CLBLM_L_X10Y136_SLICE_X13Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffafaabfbb)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_DLUT (
.I0(CLBLM_R_X11Y136_SLICE_X14Y136_BO6),
.I1(CLBLM_L_X10Y140_SLICE_X13Y140_B5Q),
.I2(CLBLM_R_X11Y134_SLICE_X14Y134_AO6),
.I3(CLBLM_R_X5Y136_SLICE_X6Y136_BQ),
.I4(CLBLM_L_X12Y135_SLICE_X17Y135_DO6),
.I5(CLBLM_L_X10Y132_SLICE_X13Y132_BO6),
.O5(CLBLM_L_X10Y136_SLICE_X13Y136_DO5),
.O6(CLBLM_L_X10Y136_SLICE_X13Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69966996f0f03333)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_CLUT (
.I0(CLBLM_L_X12Y136_SLICE_X16Y136_AQ),
.I1(CLBLM_L_X10Y140_SLICE_X13Y140_B5Q),
.I2(CLBLM_R_X11Y142_SLICE_X14Y142_AQ),
.I3(CLBLL_L_X4Y131_SLICE_X5Y131_B5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y136_SLICE_X13Y136_CO5),
.O6(CLBLM_L_X10Y136_SLICE_X13Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5e4f5e4a0a0f5e4)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y136_SLICE_X13Y136_BQ),
.I2(CLBLM_R_X11Y133_SLICE_X14Y133_AQ),
.I3(CLBLM_L_X8Y138_SLICE_X11Y138_CQ),
.I4(CLBLL_L_X4Y135_SLICE_X5Y135_CQ),
.I5(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.O5(CLBLM_L_X10Y136_SLICE_X13Y136_BO5),
.O6(CLBLM_L_X10Y136_SLICE_X13Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50ee44fa50ee44)
  ) CLBLM_L_X10Y136_SLICE_X13Y136_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y140_SLICE_X8Y140_AQ),
.I2(CLBLM_L_X10Y136_SLICE_X13Y136_AQ),
.I3(CLBLM_L_X10Y137_SLICE_X13Y137_AQ),
.I4(CLBLM_L_X12Y132_SLICE_X16Y132_AO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y136_SLICE_X13Y136_AO5),
.O6(CLBLM_L_X10Y136_SLICE_X13Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X3Y137_SLICE_X3Y137_C5Q),
.Q(CLBLM_L_X10Y137_SLICE_X12Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.Q(CLBLM_L_X10Y137_SLICE_X12Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfbbbfbbafaaafaa)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_DLUT (
.I0(CLBLM_L_X8Y136_SLICE_X11Y136_CO6),
.I1(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.I2(CLBLM_L_X10Y137_SLICE_X13Y137_BO5),
.I3(CLBLM_L_X10Y136_SLICE_X12Y136_CQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y137_SLICE_X8Y137_AQ),
.O5(CLBLM_L_X10Y137_SLICE_X12Y137_DO5),
.O6(CLBLM_L_X10Y137_SLICE_X12Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000f0aa00)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_CLUT (
.I0(CLBLM_L_X8Y135_SLICE_X10Y135_B5Q),
.I1(1'b1),
.I2(CLBLL_L_X4Y137_SLICE_X4Y137_C5Q),
.I3(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I5(CLBLM_L_X10Y133_SLICE_X12Y133_CO6),
.O5(CLBLM_L_X10Y137_SLICE_X12Y137_CO5),
.O6(CLBLM_L_X10Y137_SLICE_X12Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbaffffffbaba)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_BLUT (
.I0(CLBLM_R_X7Y135_SLICE_X8Y135_CO6),
.I1(CLBLM_L_X10Y137_SLICE_X13Y137_BO5),
.I2(CLBLM_L_X10Y136_SLICE_X12Y136_CQ),
.I3(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.I4(CLBLM_L_X8Y136_SLICE_X11Y136_CO6),
.I5(CLBLM_R_X7Y137_SLICE_X8Y137_AQ),
.O5(CLBLM_L_X10Y137_SLICE_X12Y137_BO5),
.O6(CLBLM_L_X10Y137_SLICE_X12Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f3f3ff01ff00)
  ) CLBLM_L_X10Y137_SLICE_X12Y137_ALUT (
.I0(CLBLM_L_X10Y133_SLICE_X12Y133_CO6),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I2(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I3(CLBLM_R_X11Y140_SLICE_X14Y140_BO6),
.I4(CLBLM_L_X8Y136_SLICE_X10Y136_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X12Y137_AO5),
.O6(CLBLM_L_X10Y137_SLICE_X12Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y137_SLICE_X13Y137_AO5),
.Q(CLBLM_L_X10Y137_SLICE_X13Y137_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y137_SLICE_X13Y137_AO6),
.Q(CLBLM_L_X10Y137_SLICE_X13Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4444f4f4ff44fff4)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_DLUT (
.I0(CLBLM_R_X11Y133_SLICE_X14Y133_CO5),
.I1(CLBLM_L_X8Y137_SLICE_X11Y137_CQ),
.I2(CLBLM_R_X3Y137_SLICE_X3Y137_DQ),
.I3(CLBLM_L_X10Y140_SLICE_X12Y140_DQ),
.I4(CLBLM_L_X10Y137_SLICE_X13Y137_BO5),
.I5(CLBLM_L_X10Y137_SLICE_X13Y137_BO6),
.O5(CLBLM_L_X10Y137_SLICE_X13Y137_DO5),
.O6(CLBLM_L_X10Y137_SLICE_X13Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffdcffdcdc)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_CLUT (
.I0(CLBLM_R_X11Y133_SLICE_X14Y133_CO6),
.I1(CLBLM_L_X10Y137_SLICE_X12Y137_CO6),
.I2(CLBLM_L_X10Y138_SLICE_X13Y138_DQ),
.I3(CLBLM_R_X11Y136_SLICE_X15Y136_AO5),
.I4(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.I5(CLBLM_R_X11Y140_SLICE_X14Y140_BO6),
.O5(CLBLM_L_X10Y137_SLICE_X13Y137_CO5),
.O6(CLBLM_L_X10Y137_SLICE_X13Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff7fffffffffdf)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_BLUT (
.I0(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I1(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I2(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I4(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X13Y137_BO5),
.O6(CLBLM_L_X10Y137_SLICE_X13Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbb8888ffcc3300)
  ) CLBLM_L_X10Y137_SLICE_X13Y137_ALUT (
.I0(CLBLM_R_X7Y133_SLICE_X8Y133_D5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLM_L_X10Y132_SLICE_X12Y132_CQ),
.I4(CLBLM_R_X7Y137_SLICE_X8Y137_DQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y137_SLICE_X13Y137_AO5),
.O6(CLBLM_L_X10Y137_SLICE_X13Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y138_SLICE_X12Y138_AO6),
.Q(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y138_SLICE_X12Y138_BO6),
.Q(CLBLM_L_X10Y138_SLICE_X12Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff5fff55ff0fff00)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_DLUT (
.I0(CLBLM_L_X12Y132_SLICE_X16Y132_AO6),
.I1(1'b1),
.I2(CLBLM_R_X11Y136_SLICE_X15Y136_AO6),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_CO6),
.I4(CLBLL_L_X4Y138_SLICE_X4Y138_BQ),
.I5(CLBLM_L_X8Y140_SLICE_X10Y140_BQ),
.O5(CLBLM_L_X10Y138_SLICE_X12Y138_DO5),
.O6(CLBLM_L_X10Y138_SLICE_X12Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4400000074003000)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_CLUT (
.I0(CLBLM_L_X10Y133_SLICE_X12Y133_CO6),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I3(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I4(CLBLM_R_X7Y133_SLICE_X8Y133_D5Q),
.I5(CLBLM_R_X11Y136_SLICE_X14Y136_CO6),
.O5(CLBLM_L_X10Y138_SLICE_X12Y138_CO5),
.O6(CLBLM_L_X10Y138_SLICE_X12Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe0ef404fe0ef404)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_BLUT (
.I0(CLBLM_R_X13Y134_SLICE_X18Y134_AO6),
.I1(CLBLM_L_X10Y138_SLICE_X12Y138_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.I4(CLBLM_R_X3Y137_SLICE_X2Y137_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y138_SLICE_X12Y138_BO5),
.O6(CLBLM_L_X10Y138_SLICE_X12Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd31ec20fd31ec20)
  ) CLBLM_L_X10Y138_SLICE_X12Y138_ALUT (
.I0(CLBLM_L_X12Y132_SLICE_X16Y132_AO6),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I3(CLBLM_L_X8Y140_SLICE_X10Y140_BQ),
.I4(CLBLM_L_X8Y133_SLICE_X10Y133_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y138_SLICE_X12Y138_AO5),
.O6(CLBLM_L_X10Y138_SLICE_X12Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y138_SLICE_X13Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y138_SLICE_X13Y138_AO6),
.Q(CLBLM_L_X10Y138_SLICE_X13Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y138_SLICE_X13Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y138_SLICE_X13Y138_BO6),
.Q(CLBLM_L_X10Y138_SLICE_X13Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y138_SLICE_X13Y138_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y138_SLICE_X13Y138_CO6),
.Q(CLBLM_L_X10Y138_SLICE_X13Y138_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y138_SLICE_X13Y138_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y138_SLICE_X13Y138_DO6),
.Q(CLBLM_L_X10Y138_SLICE_X13Y138_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfacc00ccfaccfa)
  ) CLBLM_L_X10Y138_SLICE_X13Y138_DLUT (
.I0(CLBLM_L_X10Y140_SLICE_X13Y140_C5Q),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_BQ),
.I2(CLBLM_L_X10Y138_SLICE_X13Y138_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y133_SLICE_X7Y133_AQ),
.I5(CLBLL_L_X4Y135_SLICE_X4Y135_D5Q),
.O5(CLBLM_L_X10Y138_SLICE_X13Y138_DO5),
.O6(CLBLM_L_X10Y138_SLICE_X13Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffd080000fd08)
  ) CLBLM_L_X10Y138_SLICE_X13Y138_CLUT (
.I0(CLBLL_L_X4Y135_SLICE_X4Y135_D5Q),
.I1(CLBLM_L_X10Y138_SLICE_X13Y138_CQ),
.I2(CLBLM_R_X5Y133_SLICE_X7Y133_AQ),
.I3(CLBLM_R_X7Y138_SLICE_X9Y138_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X8Y133_SLICE_X10Y133_BQ),
.O5(CLBLM_L_X10Y138_SLICE_X13Y138_CO5),
.O6(CLBLM_L_X10Y138_SLICE_X13Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd88d8d8dd88dd88d)
  ) CLBLM_L_X10Y138_SLICE_X13Y138_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X12Y136_SLICE_X16Y136_A5Q),
.I2(CLBLM_R_X11Y137_SLICE_X14Y137_DO6),
.I3(CLBLM_R_X11Y140_SLICE_X15Y140_B5Q),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_L_X10Y138_SLICE_X13Y138_BO5),
.O6(CLBLM_L_X10Y138_SLICE_X13Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccffccf0cc00)
  ) CLBLM_L_X10Y138_SLICE_X13Y138_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y134_SLICE_X12Y134_BQ),
.I2(CLBLM_L_X10Y138_SLICE_X13Y138_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.I5(CLBLL_L_X4Y133_SLICE_X5Y133_AQ),
.O5(CLBLM_L_X10Y138_SLICE_X13Y138_AO5),
.O6(CLBLM_L_X10Y138_SLICE_X13Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y139_SLICE_X12Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X10Y140_SLICE_X13Y140_AQ),
.Q(CLBLM_L_X10Y139_SLICE_X12Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2220222002000200)
  ) CLBLM_L_X10Y139_SLICE_X12Y139_DLUT (
.I0(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I1(CLBLM_R_X11Y136_SLICE_X14Y136_CO6),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I3(CLBLM_R_X5Y139_SLICE_X6Y139_AQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y136_SLICE_X9Y136_BQ),
.O5(CLBLM_L_X10Y139_SLICE_X12Y139_DO5),
.O6(CLBLM_L_X10Y139_SLICE_X12Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4044404440004000)
  ) CLBLM_L_X10Y139_SLICE_X12Y139_CLUT (
.I0(CLBLM_L_X10Y133_SLICE_X12Y133_CO6),
.I1(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I2(CLBLM_L_X10Y135_SLICE_X12Y135_B5Q),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I4(1'b1),
.I5(CLBLM_L_X10Y133_SLICE_X12Y133_A5Q),
.O5(CLBLM_L_X10Y139_SLICE_X12Y139_CO5),
.O6(CLBLM_L_X10Y139_SLICE_X12Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haafaeefeaafaeefe)
  ) CLBLM_L_X10Y139_SLICE_X12Y139_BLUT (
.I0(CLBLM_L_X8Y139_SLICE_X10Y139_DO6),
.I1(CLBLL_L_X4Y136_SLICE_X4Y136_BQ),
.I2(CLBLM_L_X10Y139_SLICE_X12Y139_AQ),
.I3(CLBLM_R_X11Y136_SLICE_X15Y136_AO6),
.I4(CLBLM_L_X12Y132_SLICE_X16Y132_AO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y139_SLICE_X12Y139_BO5),
.O6(CLBLM_L_X10Y139_SLICE_X12Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00ff44444444)
  ) CLBLM_L_X10Y139_SLICE_X12Y139_ALUT (
.I0(CLBLM_R_X5Y133_SLICE_X7Y133_AQ),
.I1(CLBLL_L_X4Y135_SLICE_X4Y135_D5Q),
.I2(1'b1),
.I3(CLBLM_R_X11Y140_SLICE_X14Y140_BO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y139_SLICE_X12Y139_AO5),
.O6(CLBLM_L_X10Y139_SLICE_X12Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y139_SLICE_X12Y139_AO6),
.Q(CLBLM_L_X10Y139_SLICE_X13Y139_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y139_SLICE_X13Y139_AO6),
.Q(CLBLM_L_X10Y139_SLICE_X13Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y139_SLICE_X13Y139_BO6),
.Q(CLBLM_L_X10Y139_SLICE_X13Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y139_SLICE_X13Y139_CO6),
.Q(CLBLM_L_X10Y139_SLICE_X13Y139_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff7f5fffff3f0)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_DLUT (
.I0(CLBLM_L_X12Y134_SLICE_X17Y134_AO5),
.I1(CLBLM_R_X11Y136_SLICE_X15Y136_AO6),
.I2(CLBLM_L_X10Y135_SLICE_X13Y135_CO6),
.I3(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.I4(CLBLM_R_X11Y140_SLICE_X14Y140_BO6),
.I5(CLBLM_R_X7Y140_SLICE_X8Y140_D5Q),
.O5(CLBLM_L_X10Y139_SLICE_X13Y139_DO5),
.O6(CLBLM_L_X10Y139_SLICE_X13Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfc0cfa0afa0a)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_CLUT (
.I0(CLBLM_L_X10Y139_SLICE_X13Y139_BQ),
.I1(CLBLM_L_X10Y139_SLICE_X13Y139_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y141_SLICE_X12Y141_CQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.O5(CLBLM_L_X10Y139_SLICE_X13Y139_CO5),
.O6(CLBLM_L_X10Y139_SLICE_X13Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5f5e4a0e4e4)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y139_SLICE_X13Y139_BQ),
.I2(CLBLM_R_X11Y138_SLICE_X14Y138_AQ),
.I3(CLBLM_L_X10Y140_SLICE_X13Y140_D5Q),
.I4(CLBLM_R_X7Y131_SLICE_X9Y131_D5Q),
.I5(CLBLM_R_X7Y136_SLICE_X8Y136_A5Q),
.O5(CLBLM_L_X10Y139_SLICE_X13Y139_BO5),
.O6(CLBLM_L_X10Y139_SLICE_X13Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0cacacaca)
  ) CLBLM_L_X10Y139_SLICE_X13Y139_ALUT (
.I0(CLBLM_L_X10Y139_SLICE_X13Y139_AQ),
.I1(CLBLM_L_X10Y139_SLICE_X13Y139_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(1'b1),
.I4(CLBLM_L_X10Y140_SLICE_X13Y140_AQ),
.I5(CLBLM_R_X11Y131_SLICE_X14Y131_BO6),
.O5(CLBLM_L_X10Y139_SLICE_X13Y139_AO5),
.O6(CLBLM_L_X10Y139_SLICE_X13Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y140_SLICE_X12Y140_DO5),
.Q(CLBLM_L_X10Y140_SLICE_X12Y140_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y140_SLICE_X12Y140_AO6),
.Q(CLBLM_L_X10Y140_SLICE_X12Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y140_SLICE_X12Y140_BO6),
.Q(CLBLM_L_X10Y140_SLICE_X12Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y140_SLICE_X12Y140_CO6),
.Q(CLBLM_L_X10Y140_SLICE_X12Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y140_SLICE_X12Y140_DO6),
.Q(CLBLM_L_X10Y140_SLICE_X12Y140_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f0ffcc00ccff)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y140_SLICE_X12Y140_AQ),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y140_SLICE_X13Y140_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y140_SLICE_X12Y140_DO5),
.O6(CLBLM_L_X10Y140_SLICE_X12Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aaccaa3c)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_CLUT (
.I0(CLBLM_R_X11Y139_SLICE_X14Y139_AQ),
.I1(CLBLM_L_X10Y140_SLICE_X12Y140_CQ),
.I2(CLBLM_L_X10Y134_SLICE_X12Y134_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_DO6),
.I5(CLBLM_R_X5Y140_SLICE_X7Y140_A5Q),
.O5(CLBLM_L_X10Y140_SLICE_X12Y140_CO5),
.O6(CLBLM_L_X10Y140_SLICE_X12Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0ccf055f0aa)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_BLUT (
.I0(CLBLM_L_X8Y130_SLICE_X11Y130_BO6),
.I1(CLBLM_L_X10Y137_SLICE_X13Y137_A5Q),
.I2(CLBLM_R_X7Y136_SLICE_X8Y136_C5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y140_SLICE_X12Y140_BQ),
.I5(CLBLM_R_X5Y133_SLICE_X6Y133_A5Q),
.O5(CLBLM_L_X10Y140_SLICE_X12Y140_BO5),
.O6(CLBLM_L_X10Y140_SLICE_X12Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000ff0ff808)
  ) CLBLM_L_X10Y140_SLICE_X12Y140_ALUT (
.I0(CLBLM_L_X8Y130_SLICE_X11Y130_BO6),
.I1(CLBLM_L_X10Y140_SLICE_X12Y140_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X11Y140_SLICE_X15Y140_AQ),
.I4(CLBLM_L_X10Y140_SLICE_X12Y140_AQ),
.I5(CLBLM_R_X5Y133_SLICE_X6Y133_A5Q),
.O5(CLBLM_L_X10Y140_SLICE_X12Y140_AO5),
.O6(CLBLM_L_X10Y140_SLICE_X12Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y140_SLICE_X13Y140_BO5),
.Q(CLBLM_L_X10Y140_SLICE_X13Y140_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y140_SLICE_X13Y140_CO5),
.Q(CLBLM_L_X10Y140_SLICE_X13Y140_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y140_SLICE_X13Y140_DO5),
.Q(CLBLM_L_X10Y140_SLICE_X13Y140_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y140_SLICE_X13Y140_AO6),
.Q(CLBLM_L_X10Y140_SLICE_X13Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y140_SLICE_X13Y140_BO6),
.Q(CLBLM_L_X10Y140_SLICE_X13Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y140_SLICE_X13Y140_CO6),
.Q(CLBLM_L_X10Y140_SLICE_X13Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y140_SLICE_X13Y140_DO6),
.Q(CLBLM_L_X10Y140_SLICE_X13Y140_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0ee44ee44)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(CLBLM_R_X3Y140_SLICE_X3Y140_AQ),
.I3(CLBLM_L_X8Y140_SLICE_X10Y140_AQ),
.I4(CLBLM_L_X10Y140_SLICE_X13Y140_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y140_SLICE_X13Y140_DO5),
.O6(CLBLM_L_X10Y140_SLICE_X13Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8b8b8fc30fc30)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_CLUT (
.I0(CLBLL_L_X4Y140_SLICE_X5Y140_C5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y140_SLICE_X6Y140_CQ),
.I3(CLBLM_L_X12Y140_SLICE_X16Y140_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y140_SLICE_X13Y140_CO5),
.O6(CLBLM_L_X10Y140_SLICE_X13Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33cc008b8b8b8b)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_BLUT (
.I0(CLBLM_L_X10Y134_SLICE_X13Y134_A5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X11Y136_SLICE_X15Y136_BO6),
.I3(CLBLM_L_X10Y137_SLICE_X13Y137_A5Q),
.I4(CLBLM_R_X11Y135_SLICE_X15Y135_BO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y140_SLICE_X13Y140_BO5),
.O6(CLBLM_L_X10Y140_SLICE_X13Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeffecfc22332030)
  ) CLBLM_L_X10Y140_SLICE_X13Y140_ALUT (
.I0(CLBLM_R_X5Y133_SLICE_X7Y133_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y140_SLICE_X13Y140_AQ),
.I3(CLBLL_L_X4Y135_SLICE_X4Y135_D5Q),
.I4(CLBLL_L_X4Y140_SLICE_X5Y140_C5Q),
.I5(CLBLM_L_X8Y133_SLICE_X11Y133_B5Q),
.O5(CLBLM_L_X10Y140_SLICE_X13Y140_AO5),
.O6(CLBLM_L_X10Y140_SLICE_X13Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y141_SLICE_X12Y141_CO5),
.Q(CLBLM_L_X10Y141_SLICE_X12Y141_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y141_SLICE_X12Y141_AO6),
.Q(CLBLM_L_X10Y141_SLICE_X12Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y141_SLICE_X12Y141_BO6),
.Q(CLBLM_L_X10Y141_SLICE_X12Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y141_SLICE_X12Y141_CO6),
.Q(CLBLM_L_X10Y141_SLICE_X12Y141_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f0f077ffffff)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_DLUT (
.I0(CLBLM_R_X7Y142_SLICE_X9Y142_DO5),
.I1(CLBLM_L_X10Y141_SLICE_X12Y141_AQ),
.I2(CLBLM_L_X10Y134_SLICE_X12Y134_AQ),
.I3(CLBLM_L_X10Y141_SLICE_X13Y141_CQ),
.I4(CLBLM_L_X8Y141_SLICE_X10Y141_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y141_SLICE_X12Y141_DO5),
.O6(CLBLM_L_X10Y141_SLICE_X12Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaccfff000f0)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_CLUT (
.I0(CLBLM_L_X8Y138_SLICE_X11Y138_AQ),
.I1(CLBLM_L_X10Y142_SLICE_X12Y142_CO6),
.I2(CLBLM_L_X10Y142_SLICE_X12Y142_BO6),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y140_SLICE_X13Y140_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y141_SLICE_X12Y141_CO5),
.O6(CLBLM_L_X10Y141_SLICE_X12Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd1d1d1d1c0c0c0c0)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_BLUT (
.I0(CLBLM_L_X8Y141_SLICE_X10Y141_DO6),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y140_SLICE_X12Y140_CQ),
.O5(CLBLM_L_X10Y141_SLICE_X12Y141_BO5),
.O6(CLBLM_L_X10Y141_SLICE_X12Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55be14ff55fa50)
  ) CLBLM_L_X10Y141_SLICE_X12Y141_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y142_SLICE_X9Y142_DO5),
.I2(CLBLM_L_X10Y141_SLICE_X12Y141_AQ),
.I3(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.I4(CLBLM_R_X5Y140_SLICE_X7Y140_A5Q),
.I5(CLBLM_L_X10Y141_SLICE_X13Y141_CQ),
.O5(CLBLM_L_X10Y141_SLICE_X12Y141_AO5),
.O6(CLBLM_L_X10Y141_SLICE_X12Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y141_SLICE_X13Y141_AO6),
.Q(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y141_SLICE_X13Y141_BO6),
.Q(CLBLM_L_X10Y141_SLICE_X13Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y141_SLICE_X13Y141_CO6),
.Q(CLBLM_L_X10Y141_SLICE_X13Y141_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y141_SLICE_X13Y141_DO6),
.Q(CLBLM_L_X10Y141_SLICE_X13Y141_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hefff2333eeff2233)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_DLUT (
.I0(CLBLM_R_X5Y140_SLICE_X7Y140_A5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_L_X10Y141_SLICE_X12Y141_DO6),
.I3(CLBLM_L_X10Y141_SLICE_X12Y141_DO5),
.I4(CLBLM_L_X8Y140_SLICE_X10Y140_CQ),
.I5(CLBLM_L_X10Y141_SLICE_X13Y141_DQ),
.O5(CLBLM_L_X10Y141_SLICE_X13Y141_DO5),
.O6(CLBLM_L_X10Y141_SLICE_X13Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0bbf0bbf0eef0ee)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_CLUT (
.I0(CLBLM_R_X5Y140_SLICE_X7Y140_A5Q),
.I1(CLBLM_L_X10Y141_SLICE_X13Y141_CQ),
.I2(CLBLM_L_X10Y136_SLICE_X12Y136_C5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y142_SLICE_X9Y142_DO5),
.O5(CLBLM_L_X10Y141_SLICE_X13Y141_CO5),
.O6(CLBLM_L_X10Y141_SLICE_X13Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaf8c0000af8c)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_BLUT (
.I0(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I1(CLBLM_L_X10Y141_SLICE_X13Y141_BQ),
.I2(CLBLL_L_X4Y135_SLICE_X5Y135_CQ),
.I3(CLBLM_L_X10Y140_SLICE_X13Y140_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X10Y139_SLICE_X13Y139_A5Q),
.O5(CLBLM_L_X10Y141_SLICE_X13Y141_BO5),
.O6(CLBLM_L_X10Y141_SLICE_X13Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff70ff5200700052)
  ) CLBLM_L_X10Y141_SLICE_X13Y141_ALUT (
.I0(CLBLM_R_X7Y133_SLICE_X8Y133_A5Q),
.I1(CLBLM_L_X8Y141_SLICE_X11Y141_BQ),
.I2(CLBLM_L_X10Y141_SLICE_X13Y141_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.I5(CLBLM_R_X7Y138_SLICE_X9Y138_CQ),
.O5(CLBLM_L_X10Y141_SLICE_X13Y141_AO5),
.O6(CLBLM_L_X10Y141_SLICE_X13Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y142_SLICE_X12Y142_AO6),
.Q(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y142_SLICE_X12Y142_DO5),
.O6(CLBLM_L_X10Y142_SLICE_X12Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h44cc14cc44cc44cc)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_CLUT (
.I0(CLBLM_L_X8Y141_SLICE_X11Y141_BQ),
.I1(CLBLM_L_X10Y141_SLICE_X12Y141_CQ),
.I2(CLBLM_L_X8Y142_SLICE_X11Y142_DO6),
.I3(CLBLM_R_X7Y133_SLICE_X8Y133_A5Q),
.I4(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.I5(CLBLM_L_X8Y142_SLICE_X11Y142_BQ),
.O5(CLBLM_L_X10Y142_SLICE_X12Y142_CO5),
.O6(CLBLM_L_X10Y142_SLICE_X12Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h30f030f030f012f0)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_BLUT (
.I0(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I1(CLBLM_L_X8Y141_SLICE_X11Y141_BQ),
.I2(CLBLM_L_X10Y141_SLICE_X12Y141_C5Q),
.I3(CLBLM_R_X7Y133_SLICE_X8Y133_A5Q),
.I4(CLBLM_L_X8Y142_SLICE_X11Y142_CO5),
.I5(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.O5(CLBLM_L_X10Y142_SLICE_X12Y142_BO5),
.O6(CLBLM_L_X10Y142_SLICE_X12Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcac0cac0cac0cfc5)
  ) CLBLM_L_X10Y142_SLICE_X12Y142_ALUT (
.I0(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I1(CLBLM_L_X10Y133_SLICE_X12Y133_A5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_DO6),
.I4(CLBLM_L_X8Y142_SLICE_X11Y142_CO5),
.I5(CLBLM_L_X8Y141_SLICE_X10Y141_CO6),
.O5(CLBLM_L_X10Y142_SLICE_X12Y142_AO5),
.O6(CLBLM_L_X10Y142_SLICE_X12Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y142_SLICE_X13Y142_DO5),
.O6(CLBLM_L_X10Y142_SLICE_X13Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y142_SLICE_X13Y142_CO5),
.O6(CLBLM_L_X10Y142_SLICE_X13Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y142_SLICE_X13Y142_BO5),
.O6(CLBLM_L_X10Y142_SLICE_X13Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y142_SLICE_X13Y142_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y142_SLICE_X13Y142_AO5),
.O6(CLBLM_L_X10Y142_SLICE_X13Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y131_SLICE_X16Y131_DO5),
.O6(CLBLM_L_X12Y131_SLICE_X16Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y131_SLICE_X16Y131_CO5),
.O6(CLBLM_L_X12Y131_SLICE_X16Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffcfc)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y136_SLICE_X5Y136_D5Q),
.I2(CLBLM_L_X8Y134_SLICE_X10Y134_A5Q),
.I3(1'b1),
.I4(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.I5(CLBLM_R_X7Y137_SLICE_X8Y137_CQ),
.O5(CLBLM_L_X12Y131_SLICE_X16Y131_BO5),
.O6(CLBLM_L_X12Y131_SLICE_X16Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffff0ff)
  ) CLBLM_L_X12Y131_SLICE_X16Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X8Y134_SLICE_X10Y134_A5Q),
.I3(CLBLL_L_X4Y136_SLICE_X5Y136_D5Q),
.I4(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.I5(CLBLM_R_X7Y137_SLICE_X8Y137_CQ),
.O5(CLBLM_L_X12Y131_SLICE_X16Y131_AO5),
.O6(CLBLM_L_X12Y131_SLICE_X16Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y131_SLICE_X17Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y131_SLICE_X17Y131_DO5),
.O6(CLBLM_L_X12Y131_SLICE_X17Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y131_SLICE_X17Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y131_SLICE_X17Y131_CO5),
.O6(CLBLM_L_X12Y131_SLICE_X17Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y131_SLICE_X17Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y131_SLICE_X17Y131_BO5),
.O6(CLBLM_L_X12Y131_SLICE_X17Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y131_SLICE_X17Y131_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y131_SLICE_X17Y131_AO5),
.O6(CLBLM_L_X12Y131_SLICE_X17Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y132_SLICE_X16Y132_DO5),
.O6(CLBLM_L_X12Y132_SLICE_X16Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y132_SLICE_X16Y132_CO5),
.O6(CLBLM_L_X12Y132_SLICE_X16Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffb)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_BLUT (
.I0(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.I1(CLBLL_L_X4Y136_SLICE_X5Y136_D5Q),
.I2(CLBLM_L_X8Y134_SLICE_X10Y134_A5Q),
.I3(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I4(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I5(CLBLM_R_X7Y137_SLICE_X8Y137_CQ),
.O5(CLBLM_L_X12Y132_SLICE_X16Y132_BO5),
.O6(CLBLM_L_X12Y132_SLICE_X16Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000100000000)
  ) CLBLM_L_X12Y132_SLICE_X16Y132_ALUT (
.I0(CLBLM_R_X11Y140_SLICE_X14Y140_BO6),
.I1(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I3(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I4(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I5(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.O5(CLBLM_L_X12Y132_SLICE_X16Y132_AO5),
.O6(CLBLM_L_X12Y132_SLICE_X16Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y132_SLICE_X17Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y132_SLICE_X17Y132_DO5),
.O6(CLBLM_L_X12Y132_SLICE_X17Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y132_SLICE_X17Y132_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y132_SLICE_X17Y132_CO5),
.O6(CLBLM_L_X12Y132_SLICE_X17Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y132_SLICE_X17Y132_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y132_SLICE_X17Y132_BO5),
.O6(CLBLM_L_X12Y132_SLICE_X17Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y132_SLICE_X17Y132_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y132_SLICE_X17Y132_AO5),
.O6(CLBLM_L_X12Y132_SLICE_X17Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0505030301010)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_DLUT (
.I0(CLBLM_R_X3Y133_SLICE_X3Y133_BQ),
.I1(CLBLM_R_X3Y133_SLICE_X3Y133_B5Q),
.I2(CLBLM_L_X12Y133_SLICE_X17Y133_DO6),
.I3(1'b1),
.I4(CLBLM_L_X8Y136_SLICE_X11Y136_CO5),
.I5(CLBLM_L_X12Y134_SLICE_X17Y134_AO5),
.O5(CLBLM_L_X12Y133_SLICE_X16Y133_DO5),
.O6(CLBLM_L_X12Y133_SLICE_X16Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4000000000000000)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_CLUT (
.I0(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I1(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I3(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I4(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I5(CLBLM_R_X5Y137_SLICE_X7Y137_AQ),
.O5(CLBLM_L_X12Y133_SLICE_X16Y133_CO5),
.O6(CLBLM_L_X12Y133_SLICE_X16Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hefef0000eeef0000)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_BLUT (
.I0(CLBLM_R_X11Y133_SLICE_X15Y133_CO6),
.I1(CLBLM_R_X5Y133_SLICE_X6Y133_CO5),
.I2(CLBLM_L_X12Y133_SLICE_X17Y133_AO6),
.I3(CLBLM_L_X12Y135_SLICE_X17Y135_BO6),
.I4(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I5(CLBLM_R_X13Y134_SLICE_X18Y134_DO6),
.O5(CLBLM_L_X12Y133_SLICE_X16Y133_BO5),
.O6(CLBLM_L_X12Y133_SLICE_X16Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffbfffbb)
  ) CLBLM_L_X12Y133_SLICE_X16Y133_ALUT (
.I0(CLBLM_L_X12Y134_SLICE_X16Y134_CO6),
.I1(CLBLM_L_X12Y133_SLICE_X17Y133_DO6),
.I2(CLBLM_L_X8Y136_SLICE_X11Y136_CO5),
.I3(CLBLM_L_X12Y133_SLICE_X16Y133_BO6),
.I4(CLBLM_R_X3Y133_SLICE_X3Y133_BQ),
.I5(CLBLM_L_X12Y133_SLICE_X16Y133_CO6),
.O5(CLBLM_L_X12Y133_SLICE_X16Y133_AO5),
.O6(CLBLM_L_X12Y133_SLICE_X16Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff5533ffff)
  ) CLBLM_L_X12Y133_SLICE_X17Y133_DLUT (
.I0(CLBLM_L_X10Y132_SLICE_X12Y132_BQ),
.I1(CLBLM_R_X11Y133_SLICE_X14Y133_BQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I4(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I5(CLBLM_L_X12Y133_SLICE_X17Y133_BO6),
.O5(CLBLM_L_X12Y133_SLICE_X17Y133_DO5),
.O6(CLBLM_L_X12Y133_SLICE_X17Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000200000)
  ) CLBLM_L_X12Y133_SLICE_X17Y133_CLUT (
.I0(CLBLM_R_X7Y132_SLICE_X9Y132_D5Q),
.I1(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I3(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I4(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I5(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.O5(CLBLM_L_X12Y133_SLICE_X17Y133_CO5),
.O6(CLBLM_L_X12Y133_SLICE_X17Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffd)
  ) CLBLM_L_X12Y133_SLICE_X17Y133_BLUT (
.I0(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I1(CLBLM_L_X8Y134_SLICE_X10Y134_A5Q),
.I2(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I3(CLBLL_L_X4Y136_SLICE_X5Y136_D5Q),
.I4(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.I5(CLBLM_R_X7Y137_SLICE_X8Y137_CQ),
.O5(CLBLM_L_X12Y133_SLICE_X17Y133_BO5),
.O6(CLBLM_L_X12Y133_SLICE_X17Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000000004c)
  ) CLBLM_L_X12Y133_SLICE_X17Y133_ALUT (
.I0(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I1(CLBLL_L_X4Y136_SLICE_X5Y136_D5Q),
.I2(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I3(CLBLM_L_X8Y134_SLICE_X10Y134_A5Q),
.I4(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.I5(CLBLM_R_X7Y137_SLICE_X8Y137_CQ),
.O5(CLBLM_L_X12Y133_SLICE_X17Y133_AO5),
.O6(CLBLM_L_X12Y133_SLICE_X17Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0022002000000020)
  ) CLBLM_L_X12Y134_SLICE_X16Y134_DLUT (
.I0(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I1(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I2(CLBLM_R_X11Y133_SLICE_X14Y133_AQ),
.I3(CLBLM_L_X12Y140_SLICE_X16Y140_AO5),
.I4(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I5(CLBLM_R_X5Y137_SLICE_X7Y137_AQ),
.O5(CLBLM_L_X12Y134_SLICE_X16Y134_DO5),
.O6(CLBLM_L_X12Y134_SLICE_X16Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffff7350)
  ) CLBLM_L_X12Y134_SLICE_X16Y134_CLUT (
.I0(CLBLM_R_X11Y136_SLICE_X15Y136_AO6),
.I1(CLBLM_L_X12Y134_SLICE_X17Y134_AO5),
.I2(CLBLM_R_X3Y134_SLICE_X2Y134_AQ),
.I3(CLBLM_R_X3Y133_SLICE_X3Y133_B5Q),
.I4(CLBLM_R_X11Y140_SLICE_X14Y140_BO6),
.I5(CLBLM_L_X12Y134_SLICE_X16Y134_BO6),
.O5(CLBLM_L_X12Y134_SLICE_X16Y134_CO5),
.O6(CLBLM_L_X12Y134_SLICE_X16Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeeffeefefefffe)
  ) CLBLM_L_X12Y134_SLICE_X16Y134_BLUT (
.I0(CLBLM_R_X11Y131_SLICE_X14Y131_DO6),
.I1(CLBLM_L_X12Y135_SLICE_X16Y135_DO6),
.I2(CLBLM_R_X11Y133_SLICE_X14Y133_AQ),
.I3(CLBLM_R_X7Y132_SLICE_X9Y132_D5Q),
.I4(CLBLM_L_X12Y134_SLICE_X16Y134_AO6),
.I5(CLBLM_R_X11Y136_SLICE_X15Y136_AO5),
.O5(CLBLM_L_X12Y134_SLICE_X16Y134_BO5),
.O6(CLBLM_L_X12Y134_SLICE_X16Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffdfffffffffd)
  ) CLBLM_L_X12Y134_SLICE_X16Y134_ALUT (
.I0(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I1(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I2(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I4(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y134_SLICE_X16Y134_AO5),
.O6(CLBLM_L_X12Y134_SLICE_X16Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000005040f0f0)
  ) CLBLM_L_X12Y134_SLICE_X17Y134_DLUT (
.I0(CLBLM_R_X11Y132_SLICE_X15Y132_CO6),
.I1(CLBLM_R_X13Y134_SLICE_X18Y134_BO6),
.I2(CLBLM_L_X12Y133_SLICE_X16Y133_DO6),
.I3(CLBLM_L_X12Y133_SLICE_X17Y133_AO6),
.I4(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I5(CLBLM_L_X12Y134_SLICE_X17Y134_BO6),
.O5(CLBLM_L_X12Y134_SLICE_X17Y134_DO5),
.O6(CLBLM_L_X12Y134_SLICE_X17Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000004)
  ) CLBLM_L_X12Y134_SLICE_X17Y134_CLUT (
.I0(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I1(CLBLM_R_X3Y134_SLICE_X2Y134_AQ),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I3(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I4(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I5(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.O5(CLBLM_L_X12Y134_SLICE_X17Y134_CO5),
.O6(CLBLM_L_X12Y134_SLICE_X17Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X12Y134_SLICE_X17Y134_BLUT (
.I0(CLBLM_R_X11Y131_SLICE_X14Y131_DO6),
.I1(CLBLM_L_X12Y134_SLICE_X16Y134_DO6),
.I2(CLBLM_R_X11Y140_SLICE_X14Y140_BO6),
.I3(CLBLM_L_X12Y135_SLICE_X16Y135_DO6),
.I4(CLBLM_L_X12Y134_SLICE_X17Y134_CO6),
.I5(CLBLM_L_X12Y133_SLICE_X17Y133_CO6),
.O5(CLBLM_L_X12Y134_SLICE_X17Y134_BO5),
.O6(CLBLM_L_X12Y134_SLICE_X17Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff7fff7ffff)
  ) CLBLM_L_X12Y134_SLICE_X17Y134_ALUT (
.I0(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I1(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I2(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I4(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y134_SLICE_X17Y134_AO5),
.O6(CLBLM_L_X12Y134_SLICE_X17Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000100000)
  ) CLBLM_L_X12Y135_SLICE_X16Y135_DLUT (
.I0(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I2(CLBLL_L_X4Y142_SLICE_X4Y142_A5Q),
.I3(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I4(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I5(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.O5(CLBLM_L_X12Y135_SLICE_X16Y135_DO5),
.O6(CLBLM_L_X12Y135_SLICE_X16Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55000c0c00000000)
  ) CLBLM_L_X12Y135_SLICE_X16Y135_CLUT (
.I0(CLBLM_R_X11Y132_SLICE_X15Y132_AO6),
.I1(CLBLM_L_X8Y135_SLICE_X10Y135_CQ),
.I2(CLBLM_R_X11Y131_SLICE_X15Y131_AO6),
.I3(CLBLM_R_X5Y132_SLICE_X7Y132_CQ),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I5(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.O5(CLBLM_L_X12Y135_SLICE_X16Y135_CO5),
.O6(CLBLM_L_X12Y135_SLICE_X16Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff5fffdfff0fffc)
  ) CLBLM_L_X12Y135_SLICE_X16Y135_BLUT (
.I0(CLBLM_L_X8Y136_SLICE_X11Y136_CO5),
.I1(CLBLM_R_X3Y140_SLICE_X3Y140_C5Q),
.I2(CLBLM_L_X10Y135_SLICE_X13Y135_AO6),
.I3(CLBLM_L_X10Y134_SLICE_X13Y134_DO6),
.I4(CLBLM_L_X12Y135_SLICE_X16Y135_AO6),
.I5(CLBLM_L_X8Y137_SLICE_X10Y137_BQ),
.O5(CLBLM_L_X12Y135_SLICE_X16Y135_BO5),
.O6(CLBLM_L_X12Y135_SLICE_X16Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfffffffffeffff)
  ) CLBLM_L_X12Y135_SLICE_X16Y135_ALUT (
.I0(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I1(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I2(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I3(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X12Y135_SLICE_X16Y135_AO5),
.O6(CLBLM_L_X12Y135_SLICE_X16Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffefefffffffff)
  ) CLBLM_L_X12Y135_SLICE_X17Y135_DLUT (
.I0(CLBLM_L_X12Y131_SLICE_X16Y131_AO6),
.I1(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I2(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I3(1'b1),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I5(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.O5(CLBLM_L_X12Y135_SLICE_X17Y135_DO5),
.O6(CLBLM_L_X12Y135_SLICE_X17Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdffffffffffffff)
  ) CLBLM_L_X12Y135_SLICE_X17Y135_CLUT (
.I0(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.I1(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I2(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I3(CLBLM_R_X7Y137_SLICE_X8Y137_CQ),
.I4(CLBLL_L_X4Y136_SLICE_X5Y136_D5Q),
.I5(CLBLM_L_X8Y134_SLICE_X10Y134_A5Q),
.O5(CLBLM_L_X12Y135_SLICE_X17Y135_CO5),
.O6(CLBLM_L_X12Y135_SLICE_X17Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7fff7fff7ffffff)
  ) CLBLM_L_X12Y135_SLICE_X17Y135_BLUT (
.I0(CLBLM_R_X13Y138_SLICE_X18Y138_BO6),
.I1(CLBLM_L_X12Y135_SLICE_X17Y135_CO6),
.I2(CLBLM_R_X13Y134_SLICE_X18Y134_AO6),
.I3(CLBLM_L_X12Y136_SLICE_X17Y136_BO6),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I5(CLBLM_L_X12Y135_SLICE_X17Y135_AO5),
.O5(CLBLM_L_X12Y135_SLICE_X17Y135_BO5),
.O6(CLBLM_L_X12Y135_SLICE_X17Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fffffffdfffffff)
  ) CLBLM_L_X12Y135_SLICE_X17Y135_ALUT (
.I0(CLBLL_L_X4Y136_SLICE_X5Y136_D5Q),
.I1(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I2(CLBLM_R_X7Y137_SLICE_X8Y137_CQ),
.I3(CLBLM_L_X8Y134_SLICE_X10Y134_A5Q),
.I4(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y135_SLICE_X17Y135_AO5),
.O6(CLBLM_L_X12Y135_SLICE_X17Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y136_SLICE_X16Y136_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y136_SLICE_X16Y136_AO5),
.Q(CLBLM_L_X12Y136_SLICE_X16Y136_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y136_SLICE_X16Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y136_SLICE_X16Y136_AO6),
.Q(CLBLM_L_X12Y136_SLICE_X16Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00aa00aa0cae0cae)
  ) CLBLM_L_X12Y136_SLICE_X16Y136_DLUT (
.I0(CLBLM_L_X10Y136_SLICE_X12Y136_C5Q),
.I1(CLBLM_L_X12Y136_SLICE_X16Y136_AQ),
.I2(CLBLM_L_X12Y136_SLICE_X17Y136_BO6),
.I3(CLBLM_R_X11Y134_SLICE_X14Y134_AO6),
.I4(1'b1),
.I5(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.O5(CLBLM_L_X12Y136_SLICE_X16Y136_DO5),
.O6(CLBLM_L_X12Y136_SLICE_X16Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcdcccdccffffcdcc)
  ) CLBLM_L_X12Y136_SLICE_X16Y136_CLUT (
.I0(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I1(CLBLM_L_X12Y135_SLICE_X16Y135_CO6),
.I2(CLBLM_L_X12Y136_SLICE_X17Y136_BO6),
.I3(CLBLM_L_X12Y136_SLICE_X16Y136_A5Q),
.I4(CLBLM_R_X7Y136_SLICE_X8Y136_BQ),
.I5(CLBLM_R_X11Y134_SLICE_X14Y134_AO6),
.O5(CLBLM_L_X12Y136_SLICE_X16Y136_CO5),
.O6(CLBLM_L_X12Y136_SLICE_X16Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haabaaabaffffaaba)
  ) CLBLM_L_X12Y136_SLICE_X16Y136_BLUT (
.I0(CLBLM_L_X10Y131_SLICE_X13Y131_CO6),
.I1(CLBLM_L_X12Y136_SLICE_X17Y136_BO6),
.I2(CLBLM_L_X12Y136_SLICE_X16Y136_AQ),
.I3(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I4(CLBLM_L_X10Y136_SLICE_X12Y136_C5Q),
.I5(CLBLM_R_X11Y134_SLICE_X14Y134_AO6),
.O5(CLBLM_L_X12Y136_SLICE_X16Y136_BO5),
.O6(CLBLM_L_X12Y136_SLICE_X16Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa55008d8d8d8d)
  ) CLBLM_L_X12Y136_SLICE_X16Y136_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y134_SLICE_X8Y134_CQ),
.I2(CLBLM_L_X12Y136_SLICE_X17Y136_CO6),
.I3(CLBLM_L_X12Y138_SLICE_X16Y138_BO6),
.I4(CLBLM_R_X11Y133_SLICE_X14Y133_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y136_SLICE_X16Y136_AO5),
.O6(CLBLM_L_X12Y136_SLICE_X16Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccccfcfffcfc)
  ) CLBLM_L_X12Y136_SLICE_X17Y136_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y137_SLICE_X18Y137_AO5),
.I2(CLBLM_R_X11Y136_SLICE_X14Y136_AQ),
.I3(CLBLM_R_X13Y138_SLICE_X18Y138_BO6),
.I4(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.I5(CLBLM_L_X12Y136_SLICE_X17Y136_BO6),
.O5(CLBLM_L_X12Y136_SLICE_X17Y136_DO5),
.O6(CLBLM_L_X12Y136_SLICE_X17Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0707070705050705)
  ) CLBLM_L_X12Y136_SLICE_X17Y136_CLUT (
.I0(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I1(CLBLM_L_X12Y136_SLICE_X16Y136_CO6),
.I2(CLBLM_L_X10Y136_SLICE_X12Y136_DO6),
.I3(CLBLM_L_X12Y135_SLICE_X17Y135_BO6),
.I4(CLBLM_L_X12Y136_SLICE_X17Y136_DO6),
.I5(CLBLM_L_X12Y133_SLICE_X17Y133_AO6),
.O5(CLBLM_L_X12Y136_SLICE_X17Y136_CO5),
.O6(CLBLM_L_X12Y136_SLICE_X17Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffdff)
  ) CLBLM_L_X12Y136_SLICE_X17Y136_BLUT (
.I0(CLBLL_L_X4Y136_SLICE_X5Y136_D5Q),
.I1(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.I2(CLBLM_L_X8Y134_SLICE_X10Y134_A5Q),
.I3(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I4(CLBLM_L_X12Y139_SLICE_X16Y139_AO6),
.I5(CLBLM_R_X7Y137_SLICE_X8Y137_CQ),
.O5(CLBLM_L_X12Y136_SLICE_X17Y136_BO5),
.O6(CLBLM_L_X12Y136_SLICE_X17Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffdfff77ff77)
  ) CLBLM_L_X12Y136_SLICE_X17Y136_ALUT (
.I0(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I1(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I2(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I4(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y136_SLICE_X17Y136_AO5),
.O6(CLBLM_L_X12Y136_SLICE_X17Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff000000ff0010)
  ) CLBLM_L_X12Y137_SLICE_X16Y137_DLUT (
.I0(CLBLM_L_X12Y137_SLICE_X16Y137_AO6),
.I1(CLBLM_R_X13Y137_SLICE_X18Y137_DO6),
.I2(CLBLM_L_X12Y135_SLICE_X17Y135_BO6),
.I3(CLBLM_R_X11Y132_SLICE_X14Y132_CO6),
.I4(CLBLM_L_X12Y133_SLICE_X17Y133_AO6),
.I5(CLBLM_R_X11Y137_SLICE_X15Y137_AO6),
.O5(CLBLM_L_X12Y137_SLICE_X16Y137_DO5),
.O6(CLBLM_L_X12Y137_SLICE_X16Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc00cc50dc00cc)
  ) CLBLM_L_X12Y137_SLICE_X16Y137_CLUT (
.I0(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I1(CLBLM_R_X3Y136_SLICE_X2Y136_DQ),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I3(CLBLM_L_X12Y136_SLICE_X17Y136_BO6),
.I4(CLBLM_L_X12Y140_SLICE_X16Y140_AQ),
.I5(CLBLM_L_X12Y135_SLICE_X17Y135_CO6),
.O5(CLBLM_L_X12Y137_SLICE_X16Y137_CO5),
.O6(CLBLM_L_X12Y137_SLICE_X16Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0fcf0f0f0f4)
  ) CLBLM_L_X12Y137_SLICE_X16Y137_BLUT (
.I0(RIOB33_X105Y143_IOB_X1Y144_I),
.I1(CLBLM_L_X12Y135_SLICE_X17Y135_BO6),
.I2(CLBLM_L_X12Y133_SLICE_X17Y133_AO6),
.I3(CLBLM_R_X11Y137_SLICE_X15Y137_AO6),
.I4(CLBLM_L_X12Y137_SLICE_X16Y137_AO6),
.I5(CLBLM_L_X12Y140_SLICE_X16Y140_BO6),
.O5(CLBLM_L_X12Y137_SLICE_X16Y137_BO5),
.O6(CLBLM_L_X12Y137_SLICE_X16Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc00cc00cca0ec)
  ) CLBLM_L_X12Y137_SLICE_X16Y137_ALUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I1(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.I2(CLBLM_R_X7Y139_SLICE_X8Y139_AQ),
.I3(CLBLM_L_X12Y136_SLICE_X17Y136_BO6),
.I4(CLBLM_L_X12Y135_SLICE_X17Y135_CO6),
.I5(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.O5(CLBLM_L_X12Y137_SLICE_X16Y137_AO5),
.O6(CLBLM_L_X12Y137_SLICE_X16Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffefffafffeeffaa)
  ) CLBLM_L_X12Y137_SLICE_X17Y137_DLUT (
.I0(CLBLM_L_X12Y137_SLICE_X17Y137_AO6),
.I1(CLBLM_L_X10Y136_SLICE_X13Y136_BQ),
.I2(CLBLM_R_X13Y137_SLICE_X18Y137_AO6),
.I3(CLBLM_L_X12Y139_SLICE_X17Y139_AO6),
.I4(CLBLM_R_X13Y134_SLICE_X18Y134_AO6),
.I5(CLBLM_L_X10Y137_SLICE_X12Y137_BQ),
.O5(CLBLM_L_X12Y137_SLICE_X17Y137_DO5),
.O6(CLBLM_L_X12Y137_SLICE_X17Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaababaaaaaaaba)
  ) CLBLM_L_X12Y137_SLICE_X17Y137_CLUT (
.I0(CLBLM_L_X12Y133_SLICE_X17Y133_AO6),
.I1(CLBLM_L_X12Y137_SLICE_X16Y137_CO6),
.I2(CLBLM_L_X12Y135_SLICE_X17Y135_BO6),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X12Y137_SLICE_X17Y137_DO6),
.I5(CLBLM_L_X12Y140_SLICE_X16Y140_BO6),
.O5(CLBLM_L_X12Y137_SLICE_X17Y137_CO5),
.O6(CLBLM_L_X12Y137_SLICE_X17Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffeffffff)
  ) CLBLM_L_X12Y137_SLICE_X17Y137_BLUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I1(CLBLM_R_X11Y140_SLICE_X14Y140_BO6),
.I2(CLBLM_L_X12Y131_SLICE_X16Y131_AO6),
.I3(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I4(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I5(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.O5(CLBLM_L_X12Y137_SLICE_X17Y137_BO5),
.O6(CLBLM_L_X12Y137_SLICE_X17Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0300000002000200)
  ) CLBLM_L_X12Y137_SLICE_X17Y137_ALUT (
.I0(CLBLM_L_X8Y140_SLICE_X10Y140_CQ),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I2(CLBLM_L_X12Y135_SLICE_X17Y135_CO6),
.I3(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y137_SLICE_X17Y137_AO5),
.O6(CLBLM_L_X12Y137_SLICE_X17Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7755f7f53300f3f0)
  ) CLBLM_L_X12Y138_SLICE_X16Y138_DLUT (
.I0(CLBLM_R_X13Y137_SLICE_X18Y137_AO6),
.I1(CLBLM_R_X13Y138_SLICE_X18Y138_BO6),
.I2(CLBLM_R_X11Y140_SLICE_X15Y140_AQ),
.I3(LIOB33_X0Y53_IOB_X0Y53_I),
.I4(CLBLM_R_X13Y138_SLICE_X18Y138_AO6),
.I5(CLBLM_R_X11Y138_SLICE_X14Y138_AQ),
.O5(CLBLM_L_X12Y138_SLICE_X16Y138_DO5),
.O6(CLBLM_L_X12Y138_SLICE_X16Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000002200000002)
  ) CLBLM_L_X12Y138_SLICE_X16Y138_CLUT (
.I0(CLBLM_L_X12Y135_SLICE_X17Y135_BO6),
.I1(CLBLM_L_X12Y140_SLICE_X16Y140_DO6),
.I2(CLBLM_L_X10Y141_SLICE_X13Y141_BQ),
.I3(CLBLM_L_X12Y139_SLICE_X16Y139_AO5),
.I4(CLBLM_L_X12Y138_SLICE_X16Y138_DO6),
.I5(CLBLM_L_X12Y137_SLICE_X17Y137_BO6),
.O5(CLBLM_L_X12Y138_SLICE_X16Y138_CO5),
.O6(CLBLM_L_X12Y138_SLICE_X16Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff88ffffff8a)
  ) CLBLM_L_X12Y138_SLICE_X16Y138_BLUT (
.I0(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I1(CLBLM_L_X12Y136_SLICE_X16Y136_BO6),
.I2(CLBLM_L_X12Y133_SLICE_X17Y133_AO6),
.I3(CLBLM_R_X11Y138_SLICE_X14Y138_AO6),
.I4(CLBLM_L_X10Y137_SLICE_X12Y137_BO6),
.I5(CLBLM_L_X12Y138_SLICE_X16Y138_CO6),
.O5(CLBLM_L_X12Y138_SLICE_X16Y138_BO5),
.O6(CLBLM_L_X12Y138_SLICE_X16Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaaaa31200000)
  ) CLBLM_L_X12Y138_SLICE_X16Y138_ALUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I1(CLBLM_L_X12Y135_SLICE_X17Y135_CO6),
.I2(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.I3(RIOB33_X105Y137_IOB_X1Y138_I),
.I4(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X12Y138_SLICE_X16Y138_AO5),
.O6(CLBLM_L_X12Y138_SLICE_X16Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafafaffaafffa)
  ) CLBLM_L_X12Y138_SLICE_X17Y138_DLUT (
.I0(CLBLM_L_X12Y138_SLICE_X17Y138_CO6),
.I1(1'b1),
.I2(CLBLM_R_X11Y138_SLICE_X14Y138_AQ),
.I3(CLBLM_L_X10Y141_SLICE_X13Y141_BQ),
.I4(CLBLM_R_X13Y137_SLICE_X18Y137_AO6),
.I5(CLBLM_L_X12Y137_SLICE_X17Y137_BO6),
.O5(CLBLM_L_X12Y138_SLICE_X17Y138_DO5),
.O6(CLBLM_L_X12Y138_SLICE_X17Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000500000ccdc)
  ) CLBLM_L_X12Y138_SLICE_X17Y138_CLUT (
.I0(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I1(LIOB33_X0Y53_IOB_X0Y53_I),
.I2(CLBLM_R_X11Y140_SLICE_X15Y140_AQ),
.I3(CLBLM_L_X12Y136_SLICE_X17Y136_AO5),
.I4(CLBLM_L_X12Y135_SLICE_X17Y135_AO6),
.I5(CLBLM_R_X13Y138_SLICE_X18Y138_BO5),
.O5(CLBLM_L_X12Y138_SLICE_X17Y138_CO5),
.O6(CLBLM_L_X12Y138_SLICE_X17Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000444400004454)
  ) CLBLM_L_X12Y138_SLICE_X17Y138_BLUT (
.I0(CLBLM_L_X12Y136_SLICE_X16Y136_DO6),
.I1(CLBLM_L_X12Y133_SLICE_X17Y133_AO6),
.I2(CLBLM_L_X12Y135_SLICE_X17Y135_BO6),
.I3(CLBLM_L_X12Y138_SLICE_X17Y138_DO6),
.I4(CLBLM_L_X10Y131_SLICE_X13Y131_CO6),
.I5(CLBLM_L_X12Y139_SLICE_X17Y139_CO6),
.O5(CLBLM_L_X12Y138_SLICE_X17Y138_BO5),
.O6(CLBLM_L_X12Y138_SLICE_X17Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h01110f1101510151)
  ) CLBLM_L_X12Y138_SLICE_X17Y138_ALUT (
.I0(CLBLM_L_X12Y135_SLICE_X17Y135_AO6),
.I1(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I3(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I4(CLBLM_L_X12Y131_SLICE_X16Y131_AO6),
.I5(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.O5(CLBLM_L_X12Y138_SLICE_X17Y138_AO5),
.O6(CLBLM_L_X12Y138_SLICE_X17Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0a0affffff0a)
  ) CLBLM_L_X12Y139_SLICE_X16Y139_DLUT (
.I0(RIOB33_X105Y147_IOB_X1Y147_I),
.I1(1'b1),
.I2(CLBLM_R_X13Y138_SLICE_X18Y138_BO6),
.I3(CLBLM_R_X3Y138_SLICE_X2Y138_CQ),
.I4(CLBLM_L_X12Y140_SLICE_X16Y140_BO5),
.I5(CLBLM_L_X12Y136_SLICE_X17Y136_BO6),
.O5(CLBLM_L_X12Y139_SLICE_X16Y139_DO5),
.O6(CLBLM_L_X12Y139_SLICE_X16Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f0a00000303)
  ) CLBLM_L_X12Y139_SLICE_X16Y139_CLUT (
.I0(CLBLM_R_X13Y134_SLICE_X18Y134_AO6),
.I1(CLBLM_R_X3Y138_SLICE_X2Y138_CQ),
.I2(CLBLM_L_X12Y139_SLICE_X17Y139_BO6),
.I3(CLBLM_R_X13Y138_SLICE_X18Y138_AO5),
.I4(CLBLM_L_X12Y140_SLICE_X16Y140_BO5),
.I5(CLBLM_L_X12Y136_SLICE_X17Y136_BO6),
.O5(CLBLM_L_X12Y139_SLICE_X16Y139_CO5),
.O6(CLBLM_L_X12Y139_SLICE_X16Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h22fff2ff2222f2f2)
  ) CLBLM_L_X12Y139_SLICE_X16Y139_BLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(CLBLM_R_X13Y138_SLICE_X18Y138_BO6),
.I2(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.I3(CLBLM_R_X13Y137_SLICE_X18Y137_BO6),
.I4(CLBLM_R_X13Y138_SLICE_X18Y138_AO6),
.I5(RIOB33_X105Y139_IOB_X1Y140_I),
.O5(CLBLM_L_X12Y139_SLICE_X16Y139_BO5),
.O6(CLBLM_L_X12Y139_SLICE_X16Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddddddd00006420)
  ) CLBLM_L_X12Y139_SLICE_X16Y139_ALUT (
.I0(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I2(RIOB33_X105Y139_IOB_X1Y139_I),
.I3(CLBLM_R_X11Y140_SLICE_X14Y140_CQ),
.I4(CLBLM_L_X12Y135_SLICE_X17Y135_CO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y139_SLICE_X16Y139_AO5),
.O6(CLBLM_L_X12Y139_SLICE_X16Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y139_SLICE_X17Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y139_SLICE_X17Y139_DO5),
.O6(CLBLM_L_X12Y139_SLICE_X17Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcceecceefcfefcfe)
  ) CLBLM_L_X12Y139_SLICE_X17Y139_CLUT (
.I0(CLBLM_L_X8Y140_SLICE_X11Y140_CQ),
.I1(CLBLM_L_X12Y139_SLICE_X16Y139_AO5),
.I2(RIOB33_X105Y143_IOB_X1Y143_I),
.I3(CLBLM_L_X12Y136_SLICE_X17Y136_BO6),
.I4(1'b1),
.I5(CLBLM_L_X12Y140_SLICE_X16Y140_BO6),
.O5(CLBLM_L_X12Y139_SLICE_X17Y139_CO5),
.O6(CLBLM_L_X12Y139_SLICE_X17Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000010000000)
  ) CLBLM_L_X12Y139_SLICE_X17Y139_BLUT (
.I0(CLBLM_L_X12Y135_SLICE_X17Y135_AO6),
.I1(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I2(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I4(RIOB33_X105Y147_IOB_X1Y147_I),
.I5(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.O5(CLBLM_L_X12Y139_SLICE_X17Y139_BO5),
.O6(CLBLM_L_X12Y139_SLICE_X17Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0010000000000000)
  ) CLBLM_L_X12Y139_SLICE_X17Y139_ALUT (
.I0(CLBLM_L_X12Y135_SLICE_X17Y135_AO6),
.I1(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I2(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I3(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I4(RIOB33_X105Y147_IOB_X1Y148_I),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.O5(CLBLM_L_X12Y139_SLICE_X17Y139_AO5),
.O6(CLBLM_L_X12Y139_SLICE_X17Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y140_SLICE_X16Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X11Y140_SLICE_X14Y140_DQ),
.Q(CLBLM_L_X12Y140_SLICE_X16Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3300330033007350)
  ) CLBLM_L_X12Y140_SLICE_X16Y140_DLUT (
.I0(CLBLM_L_X12Y135_SLICE_X17Y135_CO6),
.I1(CLBLM_L_X12Y136_SLICE_X17Y136_BO6),
.I2(RIOB33_X105Y143_IOB_X1Y143_I),
.I3(CLBLM_L_X8Y140_SLICE_X11Y140_CQ),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I5(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.O5(CLBLM_L_X12Y140_SLICE_X16Y140_DO5),
.O6(CLBLM_L_X12Y140_SLICE_X16Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff8f8f8ff888888)
  ) CLBLM_L_X12Y140_SLICE_X16Y140_CLUT (
.I0(CLBLM_R_X7Y139_SLICE_X8Y139_AQ),
.I1(RIOB33_X105Y143_IOB_X1Y144_I),
.I2(RIOB33_X105Y143_IOB_X1Y143_I),
.I3(CLBLM_R_X11Y140_SLICE_X14Y140_DQ),
.I4(RIOB33_X105Y141_IOB_X1Y142_I),
.I5(CLBLM_R_X11Y140_SLICE_X14Y140_CQ),
.O5(CLBLM_L_X12Y140_SLICE_X16Y140_CO5),
.O6(CLBLM_L_X12Y140_SLICE_X16Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeeee0000a280)
  ) CLBLM_L_X12Y140_SLICE_X16Y140_BLUT (
.I0(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I2(CLBLM_R_X11Y140_SLICE_X14Y140_BQ),
.I3(RIOB33_X105Y141_IOB_X1Y141_I),
.I4(CLBLM_L_X12Y135_SLICE_X17Y135_CO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y140_SLICE_X16Y140_BO5),
.O6(CLBLM_L_X12Y140_SLICE_X16Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000e023333ffff)
  ) CLBLM_L_X12Y140_SLICE_X16Y140_ALUT (
.I0(RIOB33_X105Y141_IOB_X1Y142_I),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I2(CLBLM_L_X12Y135_SLICE_X17Y135_CO6),
.I3(CLBLM_R_X11Y140_SLICE_X14Y140_DQ),
.I4(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X12Y140_SLICE_X16Y140_AO5),
.O6(CLBLM_L_X12Y140_SLICE_X16Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y140_SLICE_X17Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y140_SLICE_X17Y140_DO5),
.O6(CLBLM_L_X12Y140_SLICE_X17Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y140_SLICE_X17Y140_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y140_SLICE_X17Y140_CO5),
.O6(CLBLM_L_X12Y140_SLICE_X17Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y140_SLICE_X17Y140_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y140_SLICE_X17Y140_BO5),
.O6(CLBLM_L_X12Y140_SLICE_X17Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffefefe)
  ) CLBLM_L_X12Y140_SLICE_X17Y140_ALUT (
.I0(CLBLM_R_X13Y138_SLICE_X18Y138_CO6),
.I1(CLBLM_R_X11Y140_SLICE_X15Y140_CO5),
.I2(CLBLM_L_X12Y140_SLICE_X16Y140_CO6),
.I3(RIOB33_X105Y145_IOB_X1Y146_I),
.I4(CLBLM_L_X12Y140_SLICE_X16Y140_AQ),
.I5(CLBLM_R_X13Y137_SLICE_X18Y137_CO6),
.O5(CLBLM_L_X12Y140_SLICE_X17Y140_AO5),
.O6(CLBLM_L_X12Y140_SLICE_X17Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y141_SLICE_X16Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y141_SLICE_X16Y141_AO6),
.Q(CLBLM_L_X12Y141_SLICE_X16Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y141_SLICE_X16Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y141_SLICE_X16Y141_DO5),
.O6(CLBLM_L_X12Y141_SLICE_X16Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y141_SLICE_X16Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y141_SLICE_X16Y141_CO5),
.O6(CLBLM_L_X12Y141_SLICE_X16Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffc0c0c0c0c0c0)
  ) CLBLM_L_X12Y141_SLICE_X16Y141_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y141_IOB_X1Y141_I),
.I2(CLBLM_R_X11Y140_SLICE_X14Y140_BQ),
.I3(1'b1),
.I4(CLBLM_R_X11Y140_SLICE_X14Y140_AQ),
.I5(RIOB33_X105Y139_IOB_X1Y140_I),
.O5(CLBLM_L_X12Y141_SLICE_X16Y141_BO5),
.O6(CLBLM_L_X12Y141_SLICE_X16Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccfffffaaa)
  ) CLBLM_L_X12Y141_SLICE_X16Y141_ALUT (
.I0(CLBLM_L_X12Y141_SLICE_X16Y141_BO6),
.I1(CLBLM_R_X7Y135_SLICE_X9Y135_DQ),
.I2(CLBLM_R_X11Y138_SLICE_X14Y138_AQ),
.I3(RIOB33_X105Y139_IOB_X1Y139_I),
.I4(CLBLM_L_X12Y140_SLICE_X17Y140_AO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_L_X12Y141_SLICE_X16Y141_AO5),
.O6(CLBLM_L_X12Y141_SLICE_X16Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y141_SLICE_X17Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y141_SLICE_X17Y141_DO5),
.O6(CLBLM_L_X12Y141_SLICE_X17Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y141_SLICE_X17Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y141_SLICE_X17Y141_CO5),
.O6(CLBLM_L_X12Y141_SLICE_X17Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y141_SLICE_X17Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y141_SLICE_X17Y141_BO5),
.O6(CLBLM_L_X12Y141_SLICE_X17Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y141_SLICE_X17Y141_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y141_SLICE_X17Y141_AO5),
.O6(CLBLM_L_X12Y141_SLICE_X17Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y142_SLICE_X16Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y142_SLICE_X16Y142_DO5),
.O6(CLBLM_L_X12Y142_SLICE_X16Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y142_SLICE_X16Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y142_SLICE_X16Y142_CO5),
.O6(CLBLM_L_X12Y142_SLICE_X16Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffffccccffff)
  ) CLBLM_L_X12Y142_SLICE_X16Y142_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y138_SLICE_X16Y138_BO6),
.I2(CLBLM_R_X11Y135_SLICE_X14Y135_AO6),
.I3(1'b1),
.I4(CLBLM_L_X10Y139_SLICE_X13Y139_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X12Y142_SLICE_X16Y142_BO5),
.O6(CLBLM_L_X12Y142_SLICE_X16Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fff0fafafafaf)
  ) CLBLM_L_X12Y142_SLICE_X16Y142_ALUT (
.I0(CLBLM_L_X12Y133_SLICE_X16Y133_AO6),
.I1(1'b1),
.I2(CLBLM_L_X10Y139_SLICE_X13Y139_A5Q),
.I3(CLBLM_R_X11Y135_SLICE_X15Y135_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y142_SLICE_X16Y142_AO5),
.O6(CLBLM_L_X12Y142_SLICE_X16Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y142_SLICE_X17Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y142_SLICE_X17Y142_DO5),
.O6(CLBLM_L_X12Y142_SLICE_X17Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y142_SLICE_X17Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y142_SLICE_X17Y142_CO5),
.O6(CLBLM_L_X12Y142_SLICE_X17Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y142_SLICE_X17Y142_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y142_SLICE_X17Y142_BO5),
.O6(CLBLM_L_X12Y142_SLICE_X17Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y142_SLICE_X17Y142_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y142_SLICE_X17Y142_AO5),
.O6(CLBLM_L_X12Y142_SLICE_X17Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y143_SLICE_X16Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y143_SLICE_X16Y143_DO5),
.O6(CLBLM_L_X12Y143_SLICE_X16Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y143_SLICE_X16Y143_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y143_SLICE_X16Y143_CO5),
.O6(CLBLM_L_X12Y143_SLICE_X16Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y143_SLICE_X16Y143_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y143_SLICE_X16Y143_BO5),
.O6(CLBLM_L_X12Y143_SLICE_X16Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffffff33ff33)
  ) CLBLM_L_X12Y143_SLICE_X16Y143_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y139_SLICE_X13Y139_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X11Y139_SLICE_X15Y139_BO6),
.I4(CLBLM_L_X12Y136_SLICE_X17Y136_CO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y143_SLICE_X16Y143_AO5),
.O6(CLBLM_L_X12Y143_SLICE_X16Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y143_SLICE_X17Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y143_SLICE_X17Y143_DO5),
.O6(CLBLM_L_X12Y143_SLICE_X17Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y143_SLICE_X17Y143_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y143_SLICE_X17Y143_CO5),
.O6(CLBLM_L_X12Y143_SLICE_X17Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y143_SLICE_X17Y143_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y143_SLICE_X17Y143_BO5),
.O6(CLBLM_L_X12Y143_SLICE_X17Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y143_SLICE_X17Y143_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y143_SLICE_X17Y143_AO5),
.O6(CLBLM_L_X12Y143_SLICE_X17Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y130_SLICE_X2Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y130_SLICE_X2Y130_DO5),
.O6(CLBLM_R_X3Y130_SLICE_X2Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y130_SLICE_X2Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y130_SLICE_X2Y130_CO5),
.O6(CLBLM_R_X3Y130_SLICE_X2Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y130_SLICE_X2Y130_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y130_SLICE_X2Y130_BO5),
.O6(CLBLM_R_X3Y130_SLICE_X2Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y130_SLICE_X2Y130_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y130_SLICE_X2Y130_AO5),
.O6(CLBLM_R_X3Y130_SLICE_X2Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y130_SLICE_X3Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y130_SLICE_X3Y130_DO5),
.O6(CLBLM_R_X3Y130_SLICE_X3Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y130_SLICE_X3Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y130_SLICE_X3Y130_CO5),
.O6(CLBLM_R_X3Y130_SLICE_X3Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffafa)
  ) CLBLM_R_X3Y130_SLICE_X3Y130_BLUT (
.I0(CLBLL_L_X4Y130_SLICE_X4Y130_DQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y133_SLICE_X7Y133_BQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I5(CLBLL_L_X4Y132_SLICE_X5Y132_A5Q),
.O5(CLBLM_R_X3Y130_SLICE_X3Y130_BO5),
.O6(CLBLM_R_X3Y130_SLICE_X3Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000003)
  ) CLBLM_R_X3Y130_SLICE_X3Y130_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.I2(CLBLL_L_X4Y131_SLICE_X4Y131_D5Q),
.I3(CLBLM_R_X3Y130_SLICE_X3Y130_BO6),
.I4(CLBLM_R_X5Y133_SLICE_X7Y133_CQ),
.I5(CLBLL_L_X4Y130_SLICE_X4Y130_BQ),
.O5(CLBLM_R_X3Y130_SLICE_X3Y130_AO5),
.O6(CLBLM_R_X3Y130_SLICE_X3Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y131_SLICE_X2Y131_AO5),
.Q(CLBLM_R_X3Y131_SLICE_X2Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y132_SLICE_X2Y132_CO5),
.Q(CLBLM_R_X3Y131_SLICE_X2Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X2Y131_DO5),
.O6(CLBLM_R_X3Y131_SLICE_X2Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X2Y131_CO5),
.O6(CLBLM_R_X3Y131_SLICE_X2Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X2Y131_BO5),
.O6(CLBLM_R_X3Y131_SLICE_X2Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555f0f08800)
  ) CLBLM_R_X3Y131_SLICE_X2Y131_ALUT (
.I0(LIOB33_X0Y57_IOB_X0Y58_I),
.I1(CLBLM_R_X3Y131_SLICE_X2Y131_BQ),
.I2(CLBLM_R_X3Y132_SLICE_X2Y132_AQ),
.I3(CLBLM_R_X3Y131_SLICE_X3Y131_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X2Y131_AO5),
.O6(CLBLM_R_X3Y131_SLICE_X2Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y131_SLICE_X3Y131_BO5),
.Q(CLBLM_R_X3Y131_SLICE_X3Y131_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y131_SLICE_X3Y131_AO6),
.Q(CLBLM_R_X3Y131_SLICE_X3Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y131_SLICE_X3Y131_BO6),
.Q(CLBLM_R_X3Y131_SLICE_X3Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X3Y131_DO5),
.O6(CLBLM_R_X3Y131_SLICE_X3Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X3Y131_CO5),
.O6(CLBLM_R_X3Y131_SLICE_X3Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff006666ccccf0f0)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_BLUT (
.I0(LIOB33_X0Y57_IOB_X0Y58_I),
.I1(CLBLM_R_X3Y131_SLICE_X3Y131_BQ),
.I2(CLBLM_R_X7Y138_SLICE_X9Y138_B5Q),
.I3(CLBLM_R_X5Y135_SLICE_X7Y135_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y131_SLICE_X3Y131_BO5),
.O6(CLBLM_R_X3Y131_SLICE_X3Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0000f00f)
  ) CLBLM_R_X3Y131_SLICE_X3Y131_ALUT (
.I0(CLBLM_R_X5Y134_SLICE_X6Y134_AQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y130_SLICE_X5Y130_CO5),
.I3(CLBLM_R_X3Y131_SLICE_X3Y131_AQ),
.I4(CLBLM_R_X5Y130_SLICE_X6Y130_B5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y131_SLICE_X3Y131_AO5),
.O6(CLBLM_R_X3Y131_SLICE_X3Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y132_SLICE_X2Y132_AO6),
.Q(CLBLM_R_X3Y132_SLICE_X2Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y132_SLICE_X2Y132_BO6),
.Q(CLBLM_R_X3Y132_SLICE_X2Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y132_SLICE_X2Y132_DO5),
.O6(CLBLM_R_X3Y132_SLICE_X2Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ffffffb1e4f5a0)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y131_SLICE_X3Y131_BQ),
.I2(CLBLM_R_X3Y132_SLICE_X2Y132_BQ),
.I3(CLBLM_R_X3Y131_SLICE_X2Y131_BQ),
.I4(LIOB33_X0Y57_IOB_X0Y58_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y132_SLICE_X2Y132_CO5),
.O6(CLBLM_R_X3Y132_SLICE_X2Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeff0e00ee000e)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_BLUT (
.I0(CLBLM_R_X3Y132_SLICE_X3Y132_DQ),
.I1(CLBLM_R_X3Y132_SLICE_X2Y132_BQ),
.I2(CLBLM_R_X7Y131_SLICE_X9Y131_D5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y140_SLICE_X13Y140_D5Q),
.I5(CLBLM_R_X5Y133_SLICE_X6Y133_A5Q),
.O5(CLBLM_R_X3Y132_SLICE_X2Y132_BO5),
.O6(CLBLM_R_X3Y132_SLICE_X2Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbbb00000bbb0)
  ) CLBLM_R_X3Y132_SLICE_X2Y132_ALUT (
.I0(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I1(CLBLL_L_X4Y135_SLICE_X5Y135_CQ),
.I2(CLBLM_R_X3Y132_SLICE_X2Y132_AQ),
.I3(CLBLL_L_X4Y135_SLICE_X4Y135_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X8Y132_SLICE_X11Y132_BQ),
.O5(CLBLM_R_X3Y132_SLICE_X2Y132_AO5),
.O6(CLBLM_R_X3Y132_SLICE_X2Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y132_SLICE_X3Y132_DO5),
.Q(CLBLM_R_X3Y132_SLICE_X3Y132_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y132_SLICE_X3Y132_AO6),
.Q(CLBLM_R_X3Y132_SLICE_X3Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y132_SLICE_X3Y132_BO6),
.Q(CLBLM_R_X3Y132_SLICE_X3Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y132_SLICE_X3Y132_CO6),
.Q(CLBLM_R_X3Y132_SLICE_X3Y132_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y132_SLICE_X3Y132_DO6),
.Q(CLBLM_R_X3Y132_SLICE_X3Y132_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa5050d8d8d8d8)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y130_SLICE_X4Y130_B5Q),
.I2(CLBLM_R_X3Y135_SLICE_X3Y135_BQ),
.I3(1'b1),
.I4(CLBLM_R_X3Y133_SLICE_X2Y133_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y132_SLICE_X3Y132_DO5),
.O6(CLBLM_R_X3Y132_SLICE_X3Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbeaa1400eeaa4400)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y132_SLICE_X3Y132_CQ),
.I2(CLBLL_L_X4Y132_SLICE_X4Y132_DQ),
.I3(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.I4(CLBLM_R_X3Y139_SLICE_X3Y139_A5Q),
.I5(CLBLM_L_X8Y132_SLICE_X11Y132_CO6),
.O5(CLBLM_R_X3Y132_SLICE_X3Y132_CO5),
.O6(CLBLM_R_X3Y132_SLICE_X3Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0000000aa)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_BLUT (
.I0(CLBLL_L_X4Y132_SLICE_X4Y132_CQ),
.I1(1'b1),
.I2(CLBLM_R_X3Y138_SLICE_X3Y138_A5Q),
.I3(CLBLL_L_X4Y132_SLICE_X4Y132_AQ),
.I4(CLBLL_L_X4Y132_SLICE_X4Y132_BQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y132_SLICE_X3Y132_BO5),
.O6(CLBLM_R_X3Y132_SLICE_X3Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000044004400)
  ) CLBLM_R_X3Y132_SLICE_X3Y132_ALUT (
.I0(CLBLL_L_X4Y132_SLICE_X4Y132_CQ),
.I1(CLBLL_L_X4Y132_SLICE_X4Y132_AQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y132_SLICE_X4Y132_BQ),
.I4(CLBLM_R_X7Y137_SLICE_X8Y137_B5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y132_SLICE_X3Y132_AO5),
.O6(CLBLM_R_X3Y132_SLICE_X3Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y133_SLICE_X2Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y133_SLICE_X2Y133_AO6),
.Q(CLBLM_R_X3Y133_SLICE_X2Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y133_SLICE_X2Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y133_SLICE_X2Y133_BO6),
.Q(CLBLM_R_X3Y133_SLICE_X2Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff3fffffff)
  ) CLBLM_R_X3Y133_SLICE_X2Y133_DLUT (
.I0(1'b1),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLM_R_X7Y134_SLICE_X8Y134_CQ),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(CLBLL_L_X4Y138_SLICE_X4Y138_BQ),
.O5(CLBLM_R_X3Y133_SLICE_X2Y133_DO5),
.O6(CLBLM_R_X3Y133_SLICE_X2Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h80aa00aa00aa00aa)
  ) CLBLM_R_X3Y133_SLICE_X2Y133_CLUT (
.I0(CLBLM_L_X8Y140_SLICE_X11Y140_BQ),
.I1(CLBLM_R_X3Y131_SLICE_X2Y131_BQ),
.I2(LIOB33_X0Y57_IOB_X0Y58_I),
.I3(CLBLM_R_X3Y134_SLICE_X3Y134_AQ),
.I4(CLBLM_R_X3Y131_SLICE_X3Y131_BQ),
.I5(CLBLM_R_X3Y134_SLICE_X3Y134_BQ),
.O5(CLBLM_R_X3Y133_SLICE_X2Y133_CO5),
.O6(CLBLM_R_X3Y133_SLICE_X2Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0eeeef0f000ee)
  ) CLBLM_R_X3Y133_SLICE_X2Y133_BLUT (
.I0(CLBLL_L_X4Y133_SLICE_X5Y133_CQ),
.I1(CLBLM_R_X3Y133_SLICE_X2Y133_BQ),
.I2(CLBLL_L_X4Y132_SLICE_X5Y132_DQ),
.I3(CLBLL_L_X4Y135_SLICE_X5Y135_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.O5(CLBLM_R_X3Y133_SLICE_X2Y133_BO5),
.O6(CLBLM_R_X3Y133_SLICE_X2Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00aacccc00aa)
  ) CLBLM_R_X3Y133_SLICE_X2Y133_ALUT (
.I0(CLBLM_R_X3Y141_SLICE_X2Y141_CO6),
.I1(CLBLL_L_X4Y133_SLICE_X5Y133_DQ),
.I2(1'b1),
.I3(CLBLM_R_X3Y133_SLICE_X2Y133_DO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y133_SLICE_X2Y133_AO5),
.O6(CLBLM_R_X3Y133_SLICE_X2Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y133_SLICE_X3Y133_BO5),
.Q(CLBLM_R_X3Y133_SLICE_X3Y133_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y133_SLICE_X3Y133_AO6),
.Q(CLBLM_R_X3Y133_SLICE_X3Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y133_SLICE_X3Y133_BO6),
.Q(CLBLM_R_X3Y133_SLICE_X3Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000077ff0000)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_DLUT (
.I0(CLBLM_R_X3Y131_SLICE_X2Y131_BQ),
.I1(CLBLM_R_X3Y131_SLICE_X3Y131_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y57_IOB_X0Y58_I),
.I4(CLBLM_R_X5Y135_SLICE_X6Y135_A5Q),
.I5(CLBLM_R_X3Y134_SLICE_X3Y134_BQ),
.O5(CLBLM_R_X3Y133_SLICE_X3Y133_DO5),
.O6(CLBLM_R_X3Y133_SLICE_X3Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000001100)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_CLUT (
.I0(CLBLM_L_X8Y140_SLICE_X11Y140_BQ),
.I1(CLBLL_L_X4Y132_SLICE_X5Y132_CQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y132_SLICE_X6Y132_CO6),
.I4(CLBLM_R_X3Y134_SLICE_X3Y134_AQ),
.I5(CLBLM_R_X3Y134_SLICE_X3Y134_BQ),
.O5(CLBLM_R_X3Y133_SLICE_X3Y133_CO5),
.O6(CLBLM_R_X3Y133_SLICE_X3Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ff000cfcfc0c0)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y136_SLICE_X9Y136_A5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y132_SLICE_X5Y132_BQ),
.I4(CLBLL_L_X4Y134_SLICE_X4Y134_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y133_SLICE_X3Y133_BO5),
.O6(CLBLM_R_X3Y133_SLICE_X3Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaccccf0cc)
  ) CLBLM_R_X3Y133_SLICE_X3Y133_ALUT (
.I0(CLBLL_L_X4Y130_SLICE_X4Y130_AQ),
.I1(CLBLL_L_X4Y133_SLICE_X4Y133_CQ),
.I2(CLBLM_R_X3Y133_SLICE_X3Y133_AQ),
.I3(CLBLM_R_X7Y131_SLICE_X9Y131_D5Q),
.I4(CLBLM_L_X10Y140_SLICE_X13Y140_D5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y133_SLICE_X3Y133_AO5),
.O6(CLBLM_R_X3Y133_SLICE_X3Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y134_SLICE_X2Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X3Y134_SLICE_X3Y134_AQ),
.Q(CLBLM_R_X3Y134_SLICE_X2Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000004048c8c)
  ) CLBLM_R_X3Y134_SLICE_X2Y134_DLUT (
.I0(CLBLM_L_X8Y140_SLICE_X11Y140_BQ),
.I1(CLBLM_R_X3Y134_SLICE_X3Y134_AQ),
.I2(CLBLM_R_X7Y137_SLICE_X9Y137_D5Q),
.I3(1'b1),
.I4(CLBLM_R_X3Y135_SLICE_X2Y135_DQ),
.I5(CLBLM_R_X3Y134_SLICE_X3Y134_BQ),
.O5(CLBLM_R_X3Y134_SLICE_X2Y134_DO5),
.O6(CLBLM_R_X3Y134_SLICE_X2Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff9810ffff0000)
  ) CLBLM_R_X3Y134_SLICE_X2Y134_CLUT (
.I0(CLBLM_L_X8Y140_SLICE_X11Y140_BQ),
.I1(CLBLM_R_X3Y134_SLICE_X3Y134_AQ),
.I2(CLBLM_R_X7Y132_SLICE_X8Y132_D5Q),
.I3(CLBLM_R_X3Y132_SLICE_X2Y132_CO6),
.I4(CLBLM_R_X3Y134_SLICE_X2Y134_DO6),
.I5(CLBLM_R_X3Y134_SLICE_X3Y134_BQ),
.O5(CLBLM_R_X3Y134_SLICE_X2Y134_CO5),
.O6(CLBLM_R_X3Y134_SLICE_X2Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0fff4faf0faf0)
  ) CLBLM_R_X3Y134_SLICE_X2Y134_BLUT (
.I0(CLBLM_R_X3Y134_SLICE_X3Y134_BQ),
.I1(CLBLM_R_X7Y132_SLICE_X8Y132_D5Q),
.I2(CLBLM_R_X3Y134_SLICE_X3Y134_AQ),
.I3(CLBLM_R_X5Y135_SLICE_X6Y135_A5Q),
.I4(CLBLM_R_X3Y130_SLICE_X3Y130_AO6),
.I5(CLBLM_R_X3Y132_SLICE_X2Y132_CO6),
.O5(CLBLM_R_X3Y134_SLICE_X2Y134_BO5),
.O6(CLBLM_R_X3Y134_SLICE_X2Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha8080000a0a00000)
  ) CLBLM_R_X3Y134_SLICE_X2Y134_ALUT (
.I0(CLBLM_R_X3Y134_SLICE_X3Y134_BQ),
.I1(CLBLM_R_X3Y131_SLICE_X2Y131_AQ),
.I2(CLBLM_L_X8Y140_SLICE_X11Y140_BQ),
.I3(CLBLM_R_X3Y132_SLICE_X2Y132_CO6),
.I4(CLBLM_R_X3Y134_SLICE_X3Y134_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y134_SLICE_X2Y134_AO5),
.O6(CLBLM_R_X3Y134_SLICE_X2Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y134_SLICE_X3Y134_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y134_SLICE_X3Y134_AO5),
.Q(CLBLM_R_X3Y134_SLICE_X3Y134_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y134_SLICE_X3Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y134_SLICE_X3Y134_AO6),
.Q(CLBLM_R_X3Y134_SLICE_X3Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y134_SLICE_X3Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y134_SLICE_X3Y134_BO6),
.Q(CLBLM_R_X3Y134_SLICE_X3Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffdfffffffdffff)
  ) CLBLM_R_X3Y134_SLICE_X3Y134_DLUT (
.I0(CLBLM_L_X8Y140_SLICE_X11Y140_BQ),
.I1(CLBLM_R_X7Y132_SLICE_X8Y132_D5Q),
.I2(CLBLM_R_X3Y135_SLICE_X2Y135_DQ),
.I3(CLBLM_R_X3Y134_SLICE_X3Y134_BQ),
.I4(CLBLM_R_X3Y134_SLICE_X3Y134_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y134_SLICE_X3Y134_DO5),
.O6(CLBLM_R_X3Y134_SLICE_X3Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000555000005450)
  ) CLBLM_R_X3Y134_SLICE_X3Y134_CLUT (
.I0(CLBLM_L_X8Y140_SLICE_X11Y140_BQ),
.I1(CLBLM_R_X3Y130_SLICE_X3Y130_AO6),
.I2(CLBLM_R_X3Y134_SLICE_X3Y134_BQ),
.I3(CLBLM_R_X3Y132_SLICE_X2Y132_CO6),
.I4(CLBLM_R_X3Y134_SLICE_X3Y134_AQ),
.I5(CLBLM_R_X7Y132_SLICE_X8Y132_D5Q),
.O5(CLBLM_R_X3Y134_SLICE_X3Y134_CO5),
.O6(CLBLM_R_X3Y134_SLICE_X3Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f3f3ff00f1f1)
  ) CLBLM_R_X3Y134_SLICE_X3Y134_BLUT (
.I0(CLBLM_R_X3Y134_SLICE_X3Y134_DO6),
.I1(CLBLM_R_X5Y135_SLICE_X6Y135_A5Q),
.I2(CLBLM_R_X3Y134_SLICE_X2Y134_AO6),
.I3(CLBLM_R_X3Y140_SLICE_X3Y140_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X3Y134_SLICE_X3Y134_CO6),
.O5(CLBLM_R_X3Y134_SLICE_X3Y134_BO5),
.O6(CLBLM_R_X3Y134_SLICE_X3Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0e4e4fa50fa50)
  ) CLBLM_R_X3Y134_SLICE_X3Y134_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y134_SLICE_X2Y134_BO6),
.I2(CLBLM_R_X11Y141_SLICE_X14Y141_AQ),
.I3(CLBLM_L_X8Y139_SLICE_X11Y139_BQ),
.I4(CLBLM_R_X3Y133_SLICE_X2Y133_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y134_SLICE_X3Y134_AO5),
.O6(CLBLM_R_X3Y134_SLICE_X3Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y135_SLICE_X2Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y135_SLICE_X2Y135_AO6),
.Q(CLBLM_R_X3Y135_SLICE_X2Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y135_SLICE_X2Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y135_SLICE_X2Y135_BO6),
.Q(CLBLM_R_X3Y135_SLICE_X2Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y135_SLICE_X2Y135_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y135_SLICE_X2Y135_CO6),
.Q(CLBLM_R_X3Y135_SLICE_X2Y135_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y135_SLICE_X2Y135_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y135_SLICE_X2Y135_DO6),
.Q(CLBLM_R_X3Y135_SLICE_X2Y135_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000eccc2000)
  ) CLBLM_R_X3Y135_SLICE_X2Y135_DLUT (
.I0(CLBLM_L_X8Y140_SLICE_X11Y140_BQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y134_SLICE_X3Y134_AQ),
.I3(CLBLM_R_X7Y137_SLICE_X9Y137_D5Q),
.I4(CLBLM_R_X3Y136_SLICE_X3Y136_CQ),
.I5(CLBLM_R_X3Y134_SLICE_X3Y134_BQ),
.O5(CLBLM_R_X3Y135_SLICE_X2Y135_DO5),
.O6(CLBLM_R_X3Y135_SLICE_X2Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf0ccaaaaf0f0)
  ) CLBLM_R_X3Y135_SLICE_X2Y135_CLUT (
.I0(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.I1(CLBLM_R_X3Y135_SLICE_X2Y135_CQ),
.I2(CLBLL_L_X4Y133_SLICE_X4Y133_DQ),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X4Y136_SLICE_X4Y136_D5Q),
.O5(CLBLM_R_X3Y135_SLICE_X2Y135_CO5),
.O6(CLBLM_R_X3Y135_SLICE_X2Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000f0d8f0d8)
  ) CLBLM_R_X3Y135_SLICE_X2Y135_BLUT (
.I0(CLBLM_R_X7Y131_SLICE_X9Y131_D5Q),
.I1(CLBLM_R_X3Y135_SLICE_X2Y135_BQ),
.I2(CLBLM_R_X5Y139_SLICE_X7Y139_AQ),
.I3(CLBLM_L_X10Y140_SLICE_X13Y140_D5Q),
.I4(CLBLM_R_X3Y132_SLICE_X3Y132_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y135_SLICE_X2Y135_BO5),
.O6(CLBLM_R_X3Y135_SLICE_X2Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccfff00000)
  ) CLBLM_R_X3Y135_SLICE_X2Y135_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y132_SLICE_X9Y132_BQ),
.I2(CLBLM_R_X3Y135_SLICE_X2Y135_AQ),
.I3(CLBLM_R_X3Y137_SLICE_X2Y137_BO6),
.I4(CLBLL_L_X4Y135_SLICE_X5Y135_DO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y135_SLICE_X2Y135_AO5),
.O6(CLBLM_R_X3Y135_SLICE_X2Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y135_SLICE_X3Y135_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y135_SLICE_X3Y135_AO5),
.Q(CLBLM_R_X3Y135_SLICE_X3Y135_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y135_SLICE_X3Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y135_SLICE_X3Y135_AO6),
.Q(CLBLM_R_X3Y135_SLICE_X3Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y135_SLICE_X3Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y135_SLICE_X3Y135_BO6),
.Q(CLBLM_R_X3Y135_SLICE_X3Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y135_SLICE_X3Y135_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y135_SLICE_X3Y135_CO6),
.Q(CLBLM_R_X3Y135_SLICE_X3Y135_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y135_SLICE_X3Y135_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y135_SLICE_X3Y135_DO6),
.Q(CLBLM_R_X3Y135_SLICE_X3Y135_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff12ff0000120000)
  ) CLBLM_R_X3Y135_SLICE_X3Y135_DLUT (
.I0(CLBLL_L_X4Y138_SLICE_X4Y138_DO6),
.I1(CLBLM_R_X5Y130_SLICE_X7Y130_DQ),
.I2(CLBLM_R_X3Y135_SLICE_X3Y135_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y138_SLICE_X7Y138_AQ),
.I5(CLBLM_R_X3Y133_SLICE_X3Y133_BQ),
.O5(CLBLM_R_X3Y135_SLICE_X3Y135_DO5),
.O6(CLBLM_R_X3Y135_SLICE_X3Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hef45ef45fe54fe54)
  ) CLBLM_R_X3Y135_SLICE_X3Y135_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y130_SLICE_X7Y130_DQ),
.I2(CLBLM_R_X5Y135_SLICE_X6Y135_DO6),
.I3(CLBLM_R_X3Y135_SLICE_X3Y135_A5Q),
.I4(1'b1),
.I5(CLBLM_R_X3Y135_SLICE_X3Y135_CQ),
.O5(CLBLM_R_X3Y135_SLICE_X3Y135_CO5),
.O6(CLBLM_R_X3Y135_SLICE_X3Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaffaa3caacc)
  ) CLBLM_R_X3Y135_SLICE_X3Y135_BLUT (
.I0(CLBLM_R_X5Y134_SLICE_X7Y134_A5Q),
.I1(CLBLM_R_X3Y135_SLICE_X3Y135_BQ),
.I2(CLBLM_R_X3Y135_SLICE_X3Y135_CQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y135_SLICE_X6Y135_DO6),
.I5(CLBLM_R_X5Y130_SLICE_X7Y130_DQ),
.O5(CLBLM_R_X3Y135_SLICE_X3Y135_BO5),
.O6(CLBLM_R_X3Y135_SLICE_X3Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ccffaa00aaff)
  ) CLBLM_R_X3Y135_SLICE_X3Y135_ALUT (
.I0(CLBLM_R_X3Y140_SLICE_X3Y140_C5Q),
.I1(CLBLM_R_X3Y132_SLICE_X3Y132_DQ),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X12Y136_SLICE_X16Y136_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y135_SLICE_X3Y135_AO5),
.O6(CLBLM_R_X3Y135_SLICE_X3Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y136_SLICE_X2Y136_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y136_SLICE_X2Y136_AO5),
.Q(CLBLM_R_X3Y136_SLICE_X2Y136_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y136_SLICE_X2Y136_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y136_SLICE_X2Y136_BO5),
.Q(CLBLM_R_X3Y136_SLICE_X2Y136_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y136_SLICE_X2Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y136_SLICE_X2Y136_AO6),
.Q(CLBLM_R_X3Y136_SLICE_X2Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y136_SLICE_X2Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y136_SLICE_X2Y136_BO6),
.Q(CLBLM_R_X3Y136_SLICE_X2Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y136_SLICE_X2Y136_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y136_SLICE_X2Y136_CO6),
.Q(CLBLM_R_X3Y136_SLICE_X2Y136_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y136_SLICE_X2Y136_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y136_SLICE_X2Y136_DO6),
.Q(CLBLM_R_X3Y136_SLICE_X2Y136_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee2222fcfc3030)
  ) CLBLM_R_X3Y136_SLICE_X2Y136_DLUT (
.I0(CLBLM_R_X3Y132_SLICE_X2Y132_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X3Y136_SLICE_X2Y136_DQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y137_SLICE_X5Y137_B5Q),
.I5(CLBLM_R_X13Y134_SLICE_X18Y134_AO6),
.O5(CLBLM_R_X3Y136_SLICE_X2Y136_DO5),
.O6(CLBLM_R_X3Y136_SLICE_X2Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd0df000fd0df000)
  ) CLBLM_R_X3Y136_SLICE_X2Y136_CLUT (
.I0(CLBLL_L_X4Y135_SLICE_X4Y135_AQ),
.I1(CLBLM_R_X3Y136_SLICE_X2Y136_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y130_SLICE_X4Y130_BQ),
.I4(CLBLM_R_X3Y136_SLICE_X3Y136_DQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y136_SLICE_X2Y136_CO5),
.O6(CLBLM_R_X3Y136_SLICE_X2Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0a0acfc0cfc0)
  ) CLBLM_R_X3Y136_SLICE_X2Y136_BLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X3Y136_SLICE_X2Y136_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y136_SLICE_X4Y136_A5Q),
.I4(CLBLL_L_X4Y139_SLICE_X4Y139_CQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y136_SLICE_X2Y136_BO5),
.O6(CLBLM_R_X3Y136_SLICE_X2Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5a5aff00cccc)
  ) CLBLM_R_X3Y136_SLICE_X2Y136_ALUT (
.I0(CLBLM_R_X3Y138_SLICE_X3Y138_BO5),
.I1(CLBLM_R_X3Y136_SLICE_X3Y136_D5Q),
.I2(CLBLM_R_X3Y136_SLICE_X2Y136_AQ),
.I3(CLBLM_R_X3Y139_SLICE_X3Y139_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y136_SLICE_X2Y136_AO5),
.O6(CLBLM_R_X3Y136_SLICE_X2Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y136_SLICE_X3Y136_BO5),
.Q(CLBLM_R_X3Y136_SLICE_X3Y136_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y136_SLICE_X3Y136_CO5),
.Q(CLBLM_R_X3Y136_SLICE_X3Y136_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y136_SLICE_X3Y136_DO5),
.Q(CLBLM_R_X3Y136_SLICE_X3Y136_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y136_SLICE_X3Y136_AO6),
.Q(CLBLM_R_X3Y136_SLICE_X3Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y136_SLICE_X3Y136_BO6),
.Q(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y136_SLICE_X3Y136_CO6),
.Q(CLBLM_R_X3Y136_SLICE_X3Y136_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y136_SLICE_X3Y136_DO6),
.Q(CLBLM_R_X3Y136_SLICE_X3Y136_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0fa0afa0a)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_DLUT (
.I0(CLBLM_R_X5Y136_SLICE_X7Y136_C5Q),
.I1(CLBLL_L_X4Y134_SLICE_X4Y134_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y136_SLICE_X12Y136_CQ),
.I4(LIOB33_X0Y59_IOB_X0Y59_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y136_SLICE_X3Y136_DO5),
.O6(CLBLM_R_X3Y136_SLICE_X3Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc55aaf0f0cccc)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_CLUT (
.I0(CLBLM_R_X7Y136_SLICE_X9Y136_A5Q),
.I1(CLBLL_L_X4Y134_SLICE_X5Y134_DQ),
.I2(CLBLM_R_X7Y132_SLICE_X8Y132_BQ),
.I3(CLBLM_R_X3Y135_SLICE_X3Y135_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y136_SLICE_X3Y136_CO5),
.O6(CLBLM_R_X3Y136_SLICE_X3Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaff0055dddd8888)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y136_SLICE_X7Y136_C5Q),
.I2(1'b1),
.I3(CLBLM_L_X10Y140_SLICE_X13Y140_BQ),
.I4(CLBLL_L_X4Y133_SLICE_X5Y133_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y136_SLICE_X3Y136_BO5),
.O6(CLBLM_R_X3Y136_SLICE_X3Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0acca0cc0acca0)
  ) CLBLM_R_X3Y136_SLICE_X3Y136_ALUT (
.I0(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.I1(CLBLM_R_X3Y138_SLICE_X2Y138_BQ),
.I2(CLBLM_R_X3Y136_SLICE_X3Y136_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X8Y139_SLICE_X11Y139_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y136_SLICE_X3Y136_AO5),
.O6(CLBLM_R_X3Y136_SLICE_X3Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X2Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y137_SLICE_X2Y137_AO6),
.Q(CLBLM_R_X3Y137_SLICE_X2Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00000000)
  ) CLBLM_R_X3Y137_SLICE_X2Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X3Y136_SLICE_X3Y136_B5Q),
.I4(1'b1),
.I5(CLBLM_R_X3Y137_SLICE_X3Y137_BQ),
.O5(CLBLM_R_X3Y137_SLICE_X2Y137_DO5),
.O6(CLBLM_R_X3Y137_SLICE_X2Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0404040400000000)
  ) CLBLM_R_X3Y137_SLICE_X2Y137_CLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(CLBLM_R_X5Y137_SLICE_X7Y137_A5Q),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X3Y138_SLICE_X2Y138_AQ),
.O5(CLBLM_R_X3Y137_SLICE_X2Y137_CO5),
.O6(CLBLM_R_X3Y137_SLICE_X2Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffcdcccccc)
  ) CLBLM_R_X3Y137_SLICE_X2Y137_BLUT (
.I0(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.I1(CLBLL_L_X2Y133_SLICE_X1Y133_AO6),
.I2(CLBLL_L_X2Y138_SLICE_X1Y138_AO6),
.I3(CLBLM_R_X3Y139_SLICE_X3Y139_BQ),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_R_X3Y137_SLICE_X2Y137_CO6),
.O5(CLBLM_R_X3Y137_SLICE_X2Y137_BO5),
.O6(CLBLM_R_X3Y137_SLICE_X2Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ddddd0d0)
  ) CLBLM_R_X3Y137_SLICE_X2Y137_ALUT (
.I0(CLBLL_L_X4Y135_SLICE_X5Y135_CQ),
.I1(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I2(CLBLM_R_X3Y137_SLICE_X2Y137_AQ),
.I3(CLBLM_R_X3Y137_SLICE_X3Y137_BQ),
.I4(CLBLM_R_X3Y137_SLICE_X3Y137_A5Q),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X3Y137_SLICE_X2Y137_AO5),
.O6(CLBLM_R_X3Y137_SLICE_X2Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y137_SLICE_X3Y137_AO5),
.Q(CLBLM_R_X3Y137_SLICE_X3Y137_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y137_SLICE_X3Y137_BO5),
.Q(CLBLM_R_X3Y137_SLICE_X3Y137_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y137_SLICE_X3Y137_CO5),
.Q(CLBLM_R_X3Y137_SLICE_X3Y137_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y137_SLICE_X3Y137_DO5),
.Q(CLBLM_R_X3Y137_SLICE_X3Y137_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y137_SLICE_X3Y137_AO6),
.Q(CLBLM_R_X3Y137_SLICE_X3Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y137_SLICE_X3Y137_BO6),
.Q(CLBLM_R_X3Y137_SLICE_X3Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y137_SLICE_X3Y137_CO6),
.Q(CLBLM_R_X3Y137_SLICE_X3Y137_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y137_SLICE_X3Y137_DO6),
.Q(CLBLM_R_X3Y137_SLICE_X3Y137_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500e4e4e4e4)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y139_SLICE_X3Y139_A5Q),
.I2(CLBLM_R_X3Y137_SLICE_X3Y137_DQ),
.I3(CLBLM_L_X10Y140_SLICE_X13Y140_BQ),
.I4(CLBLM_R_X7Y139_SLICE_X8Y139_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y137_SLICE_X3Y137_DO5),
.O6(CLBLM_R_X3Y137_SLICE_X3Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000ccaaccaa)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_CLUT (
.I0(CLBLL_L_X4Y134_SLICE_X4Y134_C5Q),
.I1(CLBLM_R_X3Y137_SLICE_X3Y137_CQ),
.I2(CLBLL_L_X4Y139_SLICE_X4Y139_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y138_SLICE_X6Y138_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y137_SLICE_X3Y137_CO5),
.O6(CLBLM_R_X3Y137_SLICE_X3Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaffcc00cc)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_BLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_R_X5Y134_SLICE_X6Y134_AQ),
.I2(CLBLM_R_X3Y136_SLICE_X2Y136_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X3Y137_SLICE_X2Y137_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y137_SLICE_X3Y137_BO5),
.O6(CLBLM_R_X3Y137_SLICE_X3Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000ff0fcfc0cfc0)
  ) CLBLM_R_X3Y137_SLICE_X3Y137_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y136_SLICE_X2Y136_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X3Y135_SLICE_X3Y135_CQ),
.I4(CLBLM_L_X12Y136_SLICE_X16Y136_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y137_SLICE_X3Y137_AO5),
.O6(CLBLM_R_X3Y137_SLICE_X3Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y138_SLICE_X2Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y138_SLICE_X2Y138_AO6),
.Q(CLBLM_R_X3Y138_SLICE_X2Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y138_SLICE_X2Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y138_SLICE_X2Y138_BO6),
.Q(CLBLM_R_X3Y138_SLICE_X2Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y138_SLICE_X2Y138_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y138_SLICE_X2Y138_CO6),
.Q(CLBLM_R_X3Y138_SLICE_X2Y138_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010000000000)
  ) CLBLM_R_X3Y138_SLICE_X2Y138_DLUT (
.I0(CLBLM_R_X5Y137_SLICE_X7Y137_DO6),
.I1(CLBLM_R_X3Y137_SLICE_X3Y137_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y61_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_R_X5Y138_SLICE_X6Y138_B5Q),
.I5(CLBLM_R_X3Y141_SLICE_X2Y141_AQ),
.O5(CLBLM_R_X3Y138_SLICE_X2Y138_DO5),
.O6(CLBLM_R_X3Y138_SLICE_X2Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaffccaaaa00cc)
  ) CLBLM_R_X3Y138_SLICE_X2Y138_CLUT (
.I0(CLBLM_R_X3Y141_SLICE_X2Y141_AQ),
.I1(CLBLM_R_X3Y138_SLICE_X2Y138_CQ),
.I2(1'b1),
.I3(CLBLM_R_X13Y134_SLICE_X18Y134_AO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X3Y133_SLICE_X2Y133_BQ),
.O5(CLBLM_R_X3Y138_SLICE_X2Y138_CO5),
.O6(CLBLM_R_X3Y138_SLICE_X2Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaccaaf3aa33)
  ) CLBLM_R_X3Y138_SLICE_X2Y138_BLUT (
.I0(CLBLL_L_X4Y137_SLICE_X4Y137_CQ),
.I1(CLBLM_R_X3Y138_SLICE_X2Y138_BQ),
.I2(CLBLM_R_X3Y136_SLICE_X2Y136_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(LIOB33_X0Y55_IOB_X0Y55_I),
.I5(CLBLM_R_X3Y138_SLICE_X3Y138_BO6),
.O5(CLBLM_R_X3Y138_SLICE_X2Y138_BO5),
.O6(CLBLM_R_X3Y138_SLICE_X2Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ce02cc00cc00)
  ) CLBLM_R_X3Y138_SLICE_X2Y138_ALUT (
.I0(CLBLM_R_X3Y141_SLICE_X2Y141_CO6),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_R_X7Y135_SLICE_X9Y135_C5Q),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(CLBLM_R_X5Y137_SLICE_X7Y137_A5Q),
.O5(CLBLM_R_X3Y138_SLICE_X2Y138_AO5),
.O6(CLBLM_R_X3Y138_SLICE_X2Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y138_SLICE_X3Y138_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y138_SLICE_X3Y138_AO5),
.Q(CLBLM_R_X3Y138_SLICE_X3Y138_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y138_SLICE_X3Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y138_SLICE_X3Y138_AO6),
.Q(CLBLM_R_X3Y138_SLICE_X3Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff8000ffff0000)
  ) CLBLM_R_X3Y138_SLICE_X3Y138_DLUT (
.I0(CLBLL_L_X4Y138_SLICE_X5Y138_AQ),
.I1(CLBLM_R_X3Y138_SLICE_X3Y138_AQ),
.I2(CLBLM_R_X3Y136_SLICE_X2Y136_AQ),
.I3(CLBLM_R_X3Y138_SLICE_X3Y138_A5Q),
.I4(LIOB33_X0Y55_IOB_X0Y55_I),
.I5(CLBLM_R_X3Y138_SLICE_X2Y138_BQ),
.O5(CLBLM_R_X3Y138_SLICE_X3Y138_DO5),
.O6(CLBLM_R_X3Y138_SLICE_X3Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he6aa66aa66aa66aa)
  ) CLBLM_R_X3Y138_SLICE_X3Y138_CLUT (
.I0(CLBLL_L_X4Y138_SLICE_X5Y138_AQ),
.I1(CLBLM_R_X3Y138_SLICE_X3Y138_AQ),
.I2(CLBLM_R_X3Y136_SLICE_X2Y136_AQ),
.I3(CLBLM_R_X3Y138_SLICE_X3Y138_A5Q),
.I4(LIOB33_X0Y55_IOB_X0Y55_I),
.I5(CLBLM_R_X3Y138_SLICE_X2Y138_BQ),
.O5(CLBLM_R_X3Y138_SLICE_X3Y138_CO5),
.O6(CLBLM_R_X3Y138_SLICE_X3Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3fffffc0000000)
  ) CLBLM_R_X3Y138_SLICE_X3Y138_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y138_SLICE_X5Y138_AQ),
.I2(CLBLM_R_X3Y138_SLICE_X3Y138_AQ),
.I3(CLBLM_R_X3Y138_SLICE_X2Y138_BQ),
.I4(CLBLM_R_X3Y138_SLICE_X3Y138_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y138_SLICE_X3Y138_BO5),
.O6(CLBLM_R_X3Y138_SLICE_X3Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haf05fa508888dddd)
  ) CLBLM_R_X3Y138_SLICE_X3Y138_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y141_SLICE_X13Y141_BQ),
.I2(CLBLM_R_X3Y138_SLICE_X3Y138_AQ),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_AQ),
.I4(CLBLM_R_X3Y138_SLICE_X3Y138_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y138_SLICE_X3Y138_AO5),
.O6(CLBLM_R_X3Y138_SLICE_X3Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y139_SLICE_X2Y139_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y139_SLICE_X2Y139_CO5),
.Q(CLBLM_R_X3Y139_SLICE_X2Y139_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y139_SLICE_X2Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y139_SLICE_X2Y139_AO6),
.Q(CLBLM_R_X3Y139_SLICE_X2Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y139_SLICE_X2Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y139_SLICE_X2Y139_BO6),
.Q(CLBLM_R_X3Y139_SLICE_X2Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y139_SLICE_X2Y139_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y139_SLICE_X2Y139_CO6),
.Q(CLBLM_R_X3Y139_SLICE_X2Y139_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y139_SLICE_X2Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y139_SLICE_X2Y139_DO5),
.O6(CLBLM_R_X3Y139_SLICE_X2Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00ff00aaaa)
  ) CLBLM_R_X3Y139_SLICE_X2Y139_CLUT (
.I0(CLBLM_L_X8Y141_SLICE_X11Y141_BQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y133_SLICE_X5Y133_CQ),
.I3(CLBLM_R_X5Y139_SLICE_X6Y139_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y139_SLICE_X2Y139_CO5),
.O6(CLBLM_R_X3Y139_SLICE_X2Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aaaac300)
  ) CLBLM_R_X3Y139_SLICE_X2Y139_BLUT (
.I0(CLBLL_L_X4Y135_SLICE_X5Y135_CQ),
.I1(CLBLM_R_X3Y139_SLICE_X2Y139_BQ),
.I2(CLBLM_R_X3Y139_SLICE_X2Y139_AQ),
.I3(CLBLM_R_X3Y139_SLICE_X3Y139_CO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X8Y140_SLICE_X10Y140_DQ),
.O5(CLBLM_R_X3Y139_SLICE_X2Y139_BO5),
.O6(CLBLM_R_X3Y139_SLICE_X2Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfbbafaa15110500)
  ) CLBLM_R_X3Y139_SLICE_X2Y139_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X2Y134_SLICE_X1Y134_AO6),
.I2(CLBLM_R_X3Y139_SLICE_X2Y139_AQ),
.I3(CLBLM_R_X3Y139_SLICE_X3Y139_CO6),
.I4(CLBLM_L_X8Y140_SLICE_X10Y140_DQ),
.I5(CLBLM_R_X5Y136_SLICE_X6Y136_BQ),
.O5(CLBLM_R_X3Y139_SLICE_X2Y139_AO5),
.O6(CLBLM_R_X3Y139_SLICE_X2Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y139_SLICE_X3Y139_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y139_SLICE_X3Y139_AO5),
.Q(CLBLM_R_X3Y139_SLICE_X3Y139_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y139_SLICE_X3Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y139_SLICE_X3Y139_AO6),
.Q(CLBLM_R_X3Y139_SLICE_X3Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y139_SLICE_X3Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y141_SLICE_X3Y141_AO6),
.Q(CLBLM_R_X3Y139_SLICE_X3Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X3Y139_SLICE_X3Y139_DLUT (
.I0(CLBLM_R_X3Y137_SLICE_X3Y137_D5Q),
.I1(CLBLM_L_X8Y141_SLICE_X11Y141_BQ),
.I2(CLBLM_R_X3Y136_SLICE_X3Y136_C5Q),
.I3(CLBLM_R_X3Y139_SLICE_X3Y139_A5Q),
.I4(CLBLM_R_X3Y139_SLICE_X2Y139_C5Q),
.I5(CLBLL_L_X4Y134_SLICE_X5Y134_DQ),
.O5(CLBLM_R_X3Y139_SLICE_X3Y139_DO5),
.O6(CLBLM_R_X3Y139_SLICE_X3Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0ff00eee0ee00)
  ) CLBLM_R_X3Y139_SLICE_X3Y139_CLUT (
.I0(CLBLM_R_X3Y139_SLICE_X2Y139_AQ),
.I1(CLBLL_L_X4Y139_SLICE_X4Y139_BQ),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLL_L_X4Y141_SLICE_X5Y141_CO6),
.I4(CLBLM_R_X3Y135_SLICE_X2Y135_AQ),
.I5(CLBLM_R_X3Y139_SLICE_X2Y139_BQ),
.O5(CLBLM_R_X3Y139_SLICE_X3Y139_CO5),
.O6(CLBLM_R_X3Y139_SLICE_X3Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555544454444)
  ) CLBLM_R_X3Y139_SLICE_X3Y139_BLUT (
.I0(CLBLM_R_X3Y138_SLICE_X2Y138_DO6),
.I1(CLBLM_R_X3Y137_SLICE_X2Y137_BO6),
.I2(CLBLL_L_X4Y139_SLICE_X4Y139_BQ),
.I3(CLBLM_R_X3Y139_SLICE_X2Y139_BQ),
.I4(CLBLM_R_X3Y139_SLICE_X2Y139_AQ),
.I5(CLBLL_L_X4Y141_SLICE_X5Y141_CO6),
.O5(CLBLM_R_X3Y139_SLICE_X3Y139_BO5),
.O6(CLBLM_R_X3Y139_SLICE_X3Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3a3acacfa0afa0a)
  ) CLBLM_R_X3Y139_SLICE_X3Y139_ALUT (
.I0(CLBLM_R_X3Y139_SLICE_X2Y139_C5Q),
.I1(CLBLM_L_X10Y136_SLICE_X12Y136_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y137_SLICE_X4Y137_AQ),
.I4(CLBLM_R_X5Y140_SLICE_X6Y140_CQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y139_SLICE_X3Y139_AO5),
.O6(CLBLM_R_X3Y139_SLICE_X3Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y140_SLICE_X2Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y140_SLICE_X2Y140_DO5),
.O6(CLBLM_R_X3Y140_SLICE_X2Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y140_SLICE_X2Y140_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y140_SLICE_X2Y140_CO5),
.O6(CLBLM_R_X3Y140_SLICE_X2Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y140_SLICE_X2Y140_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y140_SLICE_X2Y140_BO5),
.O6(CLBLM_R_X3Y140_SLICE_X2Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y140_SLICE_X2Y140_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y140_SLICE_X2Y140_AO5),
.O6(CLBLM_R_X3Y140_SLICE_X2Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y140_SLICE_X3Y140_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y140_SLICE_X3Y140_CO5),
.Q(CLBLM_R_X3Y140_SLICE_X3Y140_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y140_SLICE_X3Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y140_SLICE_X3Y140_AO6),
.Q(CLBLM_R_X3Y140_SLICE_X3Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y140_SLICE_X3Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y140_SLICE_X3Y140_BO6),
.Q(CLBLM_R_X3Y140_SLICE_X3Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y140_SLICE_X3Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y140_SLICE_X3Y140_CO6),
.Q(CLBLM_R_X3Y140_SLICE_X3Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y140_SLICE_X3Y140_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y140_SLICE_X3Y140_DO6),
.Q(CLBLM_R_X3Y140_SLICE_X3Y140_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d888888d8d8888)
  ) CLBLM_R_X3Y140_SLICE_X3Y140_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y130_SLICE_X7Y130_CQ),
.I2(CLBLM_R_X3Y140_SLICE_X3Y140_DQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y141_SLICE_X7Y141_AO6),
.I5(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.O5(CLBLM_R_X3Y140_SLICE_X3Y140_DO5),
.O6(CLBLM_R_X3Y140_SLICE_X3Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0bb11bb11)
  ) CLBLM_R_X3Y140_SLICE_X3Y140_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y140_SLICE_X13Y140_BQ),
.I2(CLBLM_L_X8Y142_SLICE_X11Y142_AQ),
.I3(CLBLM_R_X3Y140_SLICE_X3Y140_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y140_SLICE_X3Y140_CO5),
.O6(CLBLM_R_X3Y140_SLICE_X3Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff33f0f0ff00)
  ) CLBLM_R_X3Y140_SLICE_X3Y140_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y135_SLICE_X2Y135_AQ),
.I2(CLBLM_R_X3Y138_SLICE_X3Y138_AQ),
.I3(CLBLM_R_X5Y133_SLICE_X7Y133_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y136_SLICE_X8Y136_AQ),
.O5(CLBLM_R_X3Y140_SLICE_X3Y140_BO5),
.O6(CLBLM_R_X3Y140_SLICE_X3Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaffaaf0aa3c)
  ) CLBLM_R_X3Y140_SLICE_X3Y140_ALUT (
.I0(CLBLM_R_X3Y135_SLICE_X3Y135_AQ),
.I1(CLBLL_L_X4Y140_SLICE_X4Y140_AO5),
.I2(CLBLM_R_X3Y140_SLICE_X3Y140_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.I5(CLBLM_R_X5Y142_SLICE_X6Y142_B5Q),
.O5(CLBLM_R_X3Y140_SLICE_X3Y140_AO5),
.O6(CLBLM_R_X3Y140_SLICE_X3Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y141_SLICE_X2Y141_BO5),
.Q(CLBLM_R_X3Y141_SLICE_X2Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y141_SLICE_X2Y141_AO6),
.Q(CLBLM_R_X3Y141_SLICE_X2Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y141_SLICE_X2Y141_DO5),
.O6(CLBLM_R_X3Y141_SLICE_X2Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000010005)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_CLUT (
.I0(CLBLM_R_X7Y140_SLICE_X9Y140_BQ),
.I1(CLBLM_R_X3Y141_SLICE_X2Y141_AQ),
.I2(CLBLM_R_X3Y135_SLICE_X2Y135_AQ),
.I3(CLBLL_L_X2Y138_SLICE_X1Y138_AO5),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_R_X7Y141_SLICE_X8Y141_BO6),
.O5(CLBLM_R_X3Y141_SLICE_X2Y141_CO5),
.O6(CLBLM_R_X3Y141_SLICE_X2Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h44444444f8f00800)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_BLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(CLBLL_L_X2Y138_SLICE_X1Y138_AO5),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLL_L_X4Y135_SLICE_X4Y135_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y141_SLICE_X2Y141_BO5),
.O6(CLBLM_R_X3Y141_SLICE_X2Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00202055555555)
  ) CLBLM_R_X3Y141_SLICE_X2Y141_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLL_L_X2Y138_SLICE_X1Y138_AO5),
.I2(CLBLM_R_X3Y141_SLICE_X2Y141_AQ),
.I3(CLBLL_L_X4Y142_SLICE_X5Y142_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y141_SLICE_X2Y141_AO5),
.O6(CLBLM_R_X3Y141_SLICE_X2Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y141_SLICE_X3Y141_DO5),
.O6(CLBLM_R_X3Y141_SLICE_X3Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y141_SLICE_X3Y141_CO5),
.O6(CLBLM_R_X3Y141_SLICE_X3Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333000033330000)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y136_SLICE_X2Y136_B5Q),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X4Y130_SLICE_X4Y130_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y141_SLICE_X3Y141_BO5),
.O6(CLBLM_R_X3Y141_SLICE_X3Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf4f00400aa00aa00)
  ) CLBLM_R_X3Y141_SLICE_X3Y141_ALUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X2Y138_SLICE_X1Y138_AO5),
.I4(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y141_SLICE_X3Y141_AO5),
.O6(CLBLM_R_X3Y141_SLICE_X3Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X6Y127_DO6),
.Q(CLBLM_R_X5Y126_SLICE_X6Y126_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y126_SLICE_X6Y126_AO6),
.Q(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_DO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_CO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4444444444444444)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_BLUT (
.I0(CLBLM_R_X5Y128_SLICE_X6Y128_DO6),
.I1(LIOB33_X0Y53_IOB_X0Y54_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_BO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff000a0a0a0a)
  ) CLBLM_R_X5Y126_SLICE_X6Y126_ALUT (
.I0(CLBLM_R_X5Y126_SLICE_X6Y126_BO6),
.I1(1'b1),
.I2(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.I3(CLBLM_R_X5Y137_SLICE_X6Y137_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y126_SLICE_X6Y126_AO5),
.O6(CLBLM_R_X5Y126_SLICE_X6Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_DO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_CO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_BO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y126_SLICE_X7Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y126_SLICE_X7Y126_AO5),
.O6(CLBLM_R_X5Y126_SLICE_X7Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X6Y127_AO6),
.Q(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X6Y127_BO6),
.Q(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y127_SLICE_X6Y127_CO6),
.Q(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff0080808080)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_DLUT (
.I0(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.I2(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.I3(CLBLL_L_X4Y130_SLICE_X4Y130_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_DO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff22ff8800220088)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_CLUT (
.I0(CLBLM_R_X5Y126_SLICE_X6Y126_BO6),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.I5(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_CO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3fcffff030c0f0f)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y127_SLICE_X6Y127_DO5),
.I4(CLBLM_R_X5Y126_SLICE_X6Y126_BO6),
.I5(CLBLM_L_X8Y131_SLICE_X10Y131_CQ),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_BO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8bb8bbbbb8b8bbbb)
  ) CLBLM_R_X5Y127_SLICE_X6Y127_ALUT (
.I0(CLBLM_R_X5Y135_SLICE_X7Y135_DQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.I3(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.I4(CLBLM_R_X5Y126_SLICE_X6Y126_BO6),
.I5(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.O5(CLBLM_R_X5Y127_SLICE_X6Y127_AO5),
.O6(CLBLM_R_X5Y127_SLICE_X6Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_DO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_CO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_BO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y127_SLICE_X7Y127_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y127_SLICE_X7Y127_AO5),
.O6(CLBLM_R_X5Y127_SLICE_X7Y127_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X6Y128_AO6),
.Q(CLBLM_R_X5Y128_SLICE_X6Y128_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y128_SLICE_X6Y128_BO6),
.Q(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_DLUT (
.I0(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_AQ),
.I2(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.I3(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.I4(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.I5(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.O5(CLBLM_R_X5Y128_SLICE_X6Y128_DO5),
.O6(CLBLM_R_X5Y128_SLICE_X6Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000088000000)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_CLUT (
.I0(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.I1(CLBLM_R_X5Y127_SLICE_X6Y127_BQ),
.I2(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.I3(CLBLM_R_X5Y127_SLICE_X6Y127_CQ),
.I4(CLBLM_R_X5Y127_SLICE_X6Y127_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X6Y128_CO5),
.O6(CLBLM_R_X5Y128_SLICE_X6Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1b1e4e4a0a0a0a0)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.I2(CLBLM_R_X5Y126_SLICE_X6Y126_AQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y128_SLICE_X6Y128_CO5),
.I5(LIOB33_X0Y53_IOB_X0Y54_I),
.O5(CLBLM_R_X5Y128_SLICE_X6Y128_BO5),
.O6(CLBLM_R_X5Y128_SLICE_X6Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8b888b88b888b888)
  ) CLBLM_R_X5Y128_SLICE_X6Y128_ALUT (
.I0(CLBLM_R_X5Y142_SLICE_X6Y142_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y128_SLICE_X6Y128_AQ),
.I3(LIOB33_X0Y53_IOB_X0Y54_I),
.I4(1'b1),
.I5(CLBLM_R_X5Y128_SLICE_X6Y128_CO6),
.O5(CLBLM_R_X5Y128_SLICE_X6Y128_AO5),
.O6(CLBLM_R_X5Y128_SLICE_X6Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X7Y128_DO5),
.O6(CLBLM_R_X5Y128_SLICE_X7Y128_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X7Y128_CO5),
.O6(CLBLM_R_X5Y128_SLICE_X7Y128_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X7Y128_BO5),
.O6(CLBLM_R_X5Y128_SLICE_X7Y128_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y128_SLICE_X7Y128_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y128_SLICE_X7Y128_AO5),
.O6(CLBLM_R_X5Y128_SLICE_X7Y128_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X6Y129_AO6),
.Q(CLBLM_R_X5Y129_SLICE_X6Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y129_SLICE_X6Y129_DO5),
.O6(CLBLM_R_X5Y129_SLICE_X6Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y129_SLICE_X6Y129_CO5),
.O6(CLBLM_R_X5Y129_SLICE_X6Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y129_SLICE_X6Y129_BO5),
.O6(CLBLM_R_X5Y129_SLICE_X6Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00f0aaaa000f)
  ) CLBLM_R_X5Y129_SLICE_X6Y129_ALUT (
.I0(CLBLM_R_X5Y133_SLICE_X6Y133_B5Q),
.I1(1'b1),
.I2(CLBLM_R_X5Y129_SLICE_X6Y129_AQ),
.I3(CLBLM_R_X5Y130_SLICE_X6Y130_B5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y130_SLICE_X6Y130_CO6),
.O5(CLBLM_R_X5Y129_SLICE_X6Y129_AO5),
.O6(CLBLM_R_X5Y129_SLICE_X6Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X7Y129_BO5),
.Q(CLBLM_R_X5Y129_SLICE_X7Y129_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X7Y129_AO6),
.Q(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y129_SLICE_X7Y129_BO6),
.Q(CLBLM_R_X5Y129_SLICE_X7Y129_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y129_SLICE_X7Y129_DO5),
.O6(CLBLM_R_X5Y129_SLICE_X7Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y129_SLICE_X7Y129_CO5),
.O6(CLBLM_R_X5Y129_SLICE_X7Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee2222f3c0f3c0)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_BLUT (
.I0(RIOB33_X105Y107_IOB_X1Y108_I),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.I3(RIOB33_X105Y123_IOB_X1Y123_I),
.I4(CLBLM_L_X8Y133_SLICE_X11Y133_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y129_SLICE_X7Y129_BO5),
.O6(CLBLM_R_X5Y129_SLICE_X7Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccaaccf0ccf0)
  ) CLBLM_R_X5Y129_SLICE_X7Y129_ALUT (
.I0(CLBLM_R_X5Y131_SLICE_X7Y131_CQ),
.I1(CLBLM_R_X5Y129_SLICE_X7Y129_BQ),
.I2(CLBLM_R_X5Y129_SLICE_X7Y129_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(CLBLM_R_X13Y134_SLICE_X18Y134_AO6),
.O5(CLBLM_R_X5Y129_SLICE_X7Y129_AO5),
.O6(CLBLM_R_X5Y129_SLICE_X7Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X6Y130_BO5),
.Q(CLBLM_R_X5Y130_SLICE_X6Y130_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X6Y130_AO6),
.Q(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X6Y130_BO6),
.Q(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5ff55ff5affaaffa)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_DLUT (
.I0(CLBLL_L_X4Y130_SLICE_X4Y130_BQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.I3(CLBLL_L_X4Y130_SLICE_X5Y130_B5Q),
.I4(1'b1),
.I5(CLBLM_R_X5Y126_SLICE_X6Y126_A5Q),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_DO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffffffffffff)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_CLUT (
.I0(CLBLM_R_X3Y131_SLICE_X3Y131_AQ),
.I1(CLBLM_R_X7Y131_SLICE_X8Y131_A5Q),
.I2(CLBLL_L_X4Y134_SLICE_X4Y134_CQ),
.I3(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I4(CLBLL_L_X4Y130_SLICE_X5Y130_AQ),
.I5(CLBLM_R_X5Y130_SLICE_X7Y130_BQ),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_CO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa5050dd88dd88)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.I2(CLBLL_L_X4Y130_SLICE_X4Y130_BQ),
.I3(CLBLM_R_X5Y133_SLICE_X6Y133_AQ),
.I4(CLBLM_L_X8Y132_SLICE_X10Y132_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_BO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f04400f0f00000)
  ) CLBLM_R_X5Y130_SLICE_X6Y130_ALUT (
.I0(CLBLL_L_X4Y130_SLICE_X5Y130_DO6),
.I1(CLBLM_R_X3Y131_SLICE_X3Y131_AQ),
.I2(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.I3(CLBLM_R_X7Y131_SLICE_X8Y131_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y131_SLICE_X6Y131_CO5),
.O5(CLBLM_R_X5Y130_SLICE_X6Y130_AO5),
.O6(CLBLM_R_X5Y130_SLICE_X6Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X7Y130_DO5),
.Q(CLBLM_R_X5Y130_SLICE_X7Y130_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X7Y130_AO6),
.Q(CLBLM_R_X5Y130_SLICE_X7Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X7Y130_BO6),
.Q(CLBLM_R_X5Y130_SLICE_X7Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X7Y130_CO6),
.Q(CLBLM_R_X5Y130_SLICE_X7Y130_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y130_SLICE_X7Y130_DO6),
.Q(CLBLM_R_X5Y130_SLICE_X7Y130_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00aaaacccc)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_DLUT (
.I0(CLBLM_L_X10Y135_SLICE_X13Y135_AQ),
.I1(CLBLM_R_X7Y131_SLICE_X8Y131_C5Q),
.I2(CLBLL_L_X4Y136_SLICE_X4Y136_AQ),
.I3(CLBLM_R_X5Y133_SLICE_X7Y133_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_DO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbf15ae04bf15ae04)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y130_SLICE_X7Y130_CQ),
.I2(CLBLM_R_X5Y139_SLICE_X7Y139_B5Q),
.I3(CLBLM_L_X8Y135_SLICE_X10Y135_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_CO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f606f000fc0c)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_BLUT (
.I0(CLBLL_L_X4Y134_SLICE_X4Y134_CQ),
.I1(CLBLM_R_X5Y130_SLICE_X7Y130_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y134_SLICE_X4Y134_A5Q),
.I4(CLBLM_R_X5Y130_SLICE_X6Y130_B5Q),
.I5(CLBLM_R_X7Y131_SLICE_X8Y131_A5Q),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_BO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0ccccfa50)
  ) CLBLM_R_X5Y130_SLICE_X7Y130_ALUT (
.I0(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.I1(CLBLM_R_X5Y128_SLICE_X6Y128_BQ),
.I2(CLBLM_R_X5Y130_SLICE_X7Y130_AQ),
.I3(CLBLL_L_X4Y130_SLICE_X5Y130_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y135_SLICE_X9Y135_C5Q),
.O5(CLBLM_R_X5Y130_SLICE_X7Y130_AO5),
.O6(CLBLM_R_X5Y130_SLICE_X7Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X6Y131_AO6),
.Q(CLBLM_R_X5Y131_SLICE_X6Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X6Y131_BO6),
.Q(CLBLM_R_X5Y131_SLICE_X6Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffff6fff6)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_DLUT (
.I0(CLBLL_L_X4Y130_SLICE_X5Y130_AQ),
.I1(CLBLL_L_X4Y134_SLICE_X4Y134_A5Q),
.I2(CLBLL_L_X4Y131_SLICE_X5Y131_CO6),
.I3(CLBLM_R_X5Y131_SLICE_X6Y131_CO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y131_SLICE_X5Y131_DO6),
.O5(CLBLM_R_X5Y131_SLICE_X6Y131_DO5),
.O6(CLBLM_R_X5Y131_SLICE_X6Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6f6ff6f6cc00cc00)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_CLUT (
.I0(CLBLM_R_X7Y134_SLICE_X8Y134_AQ),
.I1(CLBLM_R_X5Y130_SLICE_X7Y130_BQ),
.I2(CLBLM_R_X7Y131_SLICE_X8Y131_A5Q),
.I3(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I4(CLBLM_L_X8Y132_SLICE_X10Y132_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y131_SLICE_X6Y131_CO5),
.O6(CLBLM_R_X5Y131_SLICE_X6Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafffffa0a0f0f0a)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_BLUT (
.I0(CLBLM_R_X5Y131_SLICE_X6Y131_DO6),
.I1(1'b1),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y135_SLICE_X10Y135_CQ),
.I4(CLBLM_R_X5Y129_SLICE_X6Y129_AQ),
.I5(CLBLL_L_X4Y131_SLICE_X4Y131_AQ),
.O5(CLBLM_R_X5Y131_SLICE_X6Y131_BO5),
.O6(CLBLM_R_X5Y131_SLICE_X6Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafc30aaaafc30)
  ) CLBLM_R_X5Y131_SLICE_X6Y131_ALUT (
.I0(CLBLM_R_X3Y131_SLICE_X3Y131_B5Q),
.I1(CLBLM_R_X11Y131_SLICE_X14Y131_BO6),
.I2(CLBLM_R_X5Y131_SLICE_X6Y131_AQ),
.I3(CLBLL_L_X4Y131_SLICE_X4Y131_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y131_SLICE_X6Y131_AO5),
.O6(CLBLM_R_X5Y131_SLICE_X6Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X7Y131_DO5),
.Q(CLBLM_R_X5Y131_SLICE_X7Y131_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X7Y131_AO6),
.Q(CLBLM_R_X5Y131_SLICE_X7Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X7Y131_BO6),
.Q(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X7Y131_CO6),
.Q(CLBLM_R_X5Y131_SLICE_X7Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y131_SLICE_X7Y131_DO6),
.Q(CLBLM_R_X5Y131_SLICE_X7Y131_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44f5f5a0a0)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y132_SLICE_X6Y132_AQ),
.I2(CLBLM_R_X5Y131_SLICE_X7Y131_DQ),
.I3(CLBLL_L_X4Y134_SLICE_X4Y134_DQ),
.I4(CLBLM_R_X7Y130_SLICE_X9Y130_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y131_SLICE_X7Y131_DO5),
.O6(CLBLM_R_X5Y131_SLICE_X7Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffee5544afae0504)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y131_SLICE_X7Y131_CQ),
.I2(CLBLL_L_X4Y135_SLICE_X5Y135_CQ),
.I3(CLBLL_L_X4Y140_SLICE_X5Y140_CQ),
.I4(CLBLM_R_X7Y138_SLICE_X9Y138_B5Q),
.I5(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.O5(CLBLM_R_X5Y131_SLICE_X7Y131_CO5),
.O6(CLBLM_R_X5Y131_SLICE_X7Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0afa0af303fc0c)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_BLUT (
.I0(CLBLM_R_X5Y136_SLICE_X7Y136_DQ),
.I1(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.I4(CLBLM_R_X7Y130_SLICE_X8Y130_CO6),
.I5(CLBLM_R_X5Y133_SLICE_X6Y133_A5Q),
.O5(CLBLM_R_X5Y131_SLICE_X7Y131_BO5),
.O6(CLBLM_R_X5Y131_SLICE_X7Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcff5400fc0054)
  ) CLBLM_R_X5Y131_SLICE_X7Y131_ALUT (
.I0(CLBLL_L_X4Y135_SLICE_X4Y135_D5Q),
.I1(CLBLM_R_X5Y131_SLICE_X7Y131_DQ),
.I2(CLBLM_R_X5Y131_SLICE_X7Y131_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y133_SLICE_X7Y133_AQ),
.I5(CLBLL_L_X4Y133_SLICE_X5Y133_B5Q),
.O5(CLBLM_R_X5Y131_SLICE_X7Y131_AO5),
.O6(CLBLM_R_X5Y131_SLICE_X7Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y132_SLICE_X6Y132_AO6),
.Q(CLBLM_R_X5Y132_SLICE_X6Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y132_SLICE_X6Y132_BO6),
.Q(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7fdf7fdfbfefbfe)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_DLUT (
.I0(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I1(CLBLM_R_X5Y133_SLICE_X7Y133_BQ),
.I2(CLBLM_R_X5Y130_SLICE_X6Y130_DO6),
.I3(CLBLL_L_X4Y130_SLICE_X4Y130_B5Q),
.I4(1'b1),
.I5(CLBLM_R_X11Y140_SLICE_X15Y140_BQ),
.O5(CLBLM_R_X5Y132_SLICE_X6Y132_DO5),
.O6(CLBLM_R_X5Y132_SLICE_X6Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff7fdfffffbfe)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_CLUT (
.I0(CLBLL_L_X4Y130_SLICE_X4Y130_DQ),
.I1(CLBLL_L_X4Y132_SLICE_X5Y132_A5Q),
.I2(CLBLM_R_X5Y132_SLICE_X7Y132_DO6),
.I3(CLBLM_R_X5Y132_SLICE_X7Y132_CQ),
.I4(CLBLM_R_X5Y132_SLICE_X6Y132_DO6),
.I5(CLBLL_L_X4Y133_SLICE_X4Y133_D5Q),
.O5(CLBLM_R_X5Y132_SLICE_X6Y132_CO5),
.O6(CLBLM_R_X5Y132_SLICE_X6Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fffff0f06666)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_BLUT (
.I0(CLBLM_R_X5Y133_SLICE_X6Y133_DO6),
.I1(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.I2(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y130_SLICE_X7Y130_DQ),
.O5(CLBLM_R_X5Y132_SLICE_X6Y132_BO5),
.O6(CLBLM_R_X5Y132_SLICE_X6Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fffff0f07788)
  ) CLBLM_R_X5Y132_SLICE_X6Y132_ALUT (
.I0(CLBLM_R_X5Y133_SLICE_X6Y133_DO6),
.I1(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.I2(CLBLM_R_X5Y132_SLICE_X7Y132_C5Q),
.I3(CLBLM_R_X5Y132_SLICE_X6Y132_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y130_SLICE_X7Y130_DQ),
.O5(CLBLM_R_X5Y132_SLICE_X6Y132_AO5),
.O6(CLBLM_R_X5Y132_SLICE_X6Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y132_SLICE_X7Y132_CO5),
.Q(CLBLM_R_X5Y132_SLICE_X7Y132_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y132_SLICE_X7Y132_AO6),
.Q(CLBLM_R_X5Y132_SLICE_X7Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y132_SLICE_X7Y132_BO6),
.Q(CLBLM_R_X5Y132_SLICE_X7Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y132_SLICE_X7Y132_CO6),
.Q(CLBLM_R_X5Y132_SLICE_X7Y132_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5ff55ff5affaaffa)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_DLUT (
.I0(CLBLM_R_X5Y134_SLICE_X6Y134_B5Q),
.I1(1'b1),
.I2(CLBLM_R_X5Y133_SLICE_X7Y133_CQ),
.I3(CLBLM_R_X7Y133_SLICE_X9Y133_DQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y131_SLICE_X4Y131_D5Q),
.O5(CLBLM_R_X5Y132_SLICE_X7Y132_DO5),
.O6(CLBLM_R_X5Y132_SLICE_X7Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d8f5a0f5a0)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y136_SLICE_X7Y136_DQ),
.I2(CLBLL_L_X4Y132_SLICE_X5Y132_A5Q),
.I3(CLBLL_L_X4Y134_SLICE_X4Y134_DQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y132_SLICE_X7Y132_CO5),
.O6(CLBLM_R_X5Y132_SLICE_X7Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f05544f0f05544)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_BLUT (
.I0(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.I1(CLBLM_R_X5Y132_SLICE_X7Y132_BQ),
.I2(CLBLM_L_X8Y140_SLICE_X11Y140_BQ),
.I3(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y132_SLICE_X7Y132_BO5),
.O6(CLBLM_R_X5Y132_SLICE_X7Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffa5550bbba1110)
  ) CLBLM_R_X5Y132_SLICE_X7Y132_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y135_SLICE_X4Y135_D5Q),
.I2(CLBLM_R_X5Y132_SLICE_X7Y132_AQ),
.I3(CLBLM_R_X5Y134_SLICE_X7Y134_DQ),
.I4(CLBLM_L_X8Y131_SLICE_X11Y131_C5Q),
.I5(CLBLM_R_X5Y133_SLICE_X7Y133_AQ),
.O5(CLBLM_R_X5Y132_SLICE_X7Y132_AO5),
.O6(CLBLM_R_X5Y132_SLICE_X7Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X6Y133_AO5),
.Q(CLBLM_R_X5Y133_SLICE_X6Y133_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X6Y133_BO5),
.Q(CLBLM_R_X5Y133_SLICE_X6Y133_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X6Y133_AO6),
.Q(CLBLM_R_X5Y133_SLICE_X6Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X6Y133_BO6),
.Q(CLBLM_R_X5Y133_SLICE_X6Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_DLUT (
.I0(CLBLL_L_X4Y137_SLICE_X5Y137_C5Q),
.I1(CLBLM_R_X5Y134_SLICE_X6Y134_CQ),
.I2(CLBLL_L_X4Y138_SLICE_X5Y138_DQ),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_BQ),
.I4(CLBLM_R_X3Y135_SLICE_X3Y135_BQ),
.I5(CLBLM_R_X3Y135_SLICE_X3Y135_CQ),
.O5(CLBLM_R_X5Y133_SLICE_X6Y133_DO5),
.O6(CLBLM_R_X5Y133_SLICE_X6Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3aca3ac0000aaaa)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_CLUT (
.I0(CLBLM_R_X7Y132_SLICE_X9Y132_DQ),
.I1(LIOB33_X0Y59_IOB_X0Y60_I),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y134_SLICE_X6Y134_C5Q),
.I4(CLBLM_R_X11Y134_SLICE_X14Y134_AO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y133_SLICE_X6Y133_CO5),
.O6(CLBLM_R_X5Y133_SLICE_X6Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0f5f50505)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_BLUT (
.I0(CLBLM_R_X7Y135_SLICE_X8Y135_AQ),
.I1(CLBLM_R_X7Y139_SLICE_X9Y139_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y133_SLICE_X5Y133_B5Q),
.I4(CLBLL_L_X4Y132_SLICE_X5Y132_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y133_SLICE_X6Y133_BO5),
.O6(CLBLM_R_X5Y133_SLICE_X6Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaccccf0f0aaaa)
  ) CLBLM_R_X5Y133_SLICE_X6Y133_ALUT (
.I0(CLBLM_R_X7Y133_SLICE_X9Y133_A5Q),
.I1(CLBLM_R_X5Y134_SLICE_X7Y134_D5Q),
.I2(CLBLM_R_X5Y137_SLICE_X6Y137_CQ),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y133_SLICE_X6Y133_AO5),
.O6(CLBLM_R_X5Y133_SLICE_X6Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X7Y133_AO5),
.Q(CLBLM_R_X5Y133_SLICE_X7Y133_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X7Y133_BO5),
.Q(CLBLM_R_X5Y133_SLICE_X7Y133_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X7Y133_CO5),
.Q(CLBLM_R_X5Y133_SLICE_X7Y133_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X7Y133_AO6),
.Q(CLBLM_R_X5Y133_SLICE_X7Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X7Y133_BO6),
.Q(CLBLM_R_X5Y133_SLICE_X7Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X7Y133_CO6),
.Q(CLBLM_R_X5Y133_SLICE_X7Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X7Y133_DO6),
.Q(CLBLM_R_X5Y133_SLICE_X7Y133_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55ff55fb51ff55)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y130_SLICE_X9Y130_BQ),
.I2(CLBLM_R_X3Y135_SLICE_X3Y135_BQ),
.I3(CLBLL_L_X4Y132_SLICE_X4Y132_AQ),
.I4(CLBLL_L_X4Y138_SLICE_X5Y138_DQ),
.I5(CLBLM_R_X3Y135_SLICE_X3Y135_CQ),
.O5(CLBLM_R_X5Y133_SLICE_X7Y133_DO5),
.O6(CLBLM_R_X5Y133_SLICE_X7Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa5500e4e4e4e4)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y134_SLICE_X3Y134_A5Q),
.I2(CLBLM_R_X7Y134_SLICE_X8Y134_C5Q),
.I3(CLBLM_R_X5Y135_SLICE_X6Y135_A5Q),
.I4(CLBLM_R_X5Y133_SLICE_X7Y133_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y133_SLICE_X7Y133_CO5),
.O6(CLBLM_R_X5Y133_SLICE_X7Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaacccccccc00ff)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_BLUT (
.I0(CLBLM_R_X7Y133_SLICE_X8Y133_CQ),
.I1(CLBLL_L_X4Y131_SLICE_X4Y131_D5Q),
.I2(1'b1),
.I3(CLBLM_L_X10Y140_SLICE_X13Y140_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y133_SLICE_X7Y133_BO5),
.O6(CLBLM_R_X5Y133_SLICE_X7Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afa0cfcfc0c0)
  ) CLBLM_R_X5Y133_SLICE_X7Y133_ALUT (
.I0(CLBLM_R_X5Y135_SLICE_X6Y135_A5Q),
.I1(CLBLM_R_X5Y134_SLICE_X7Y134_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(RIOB33_X105Y109_IOB_X1Y109_I),
.I4(CLBLM_L_X10Y131_SLICE_X12Y131_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y133_SLICE_X7Y133_AO5),
.O6(CLBLM_R_X5Y133_SLICE_X7Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X6Y134_AO5),
.Q(CLBLM_R_X5Y134_SLICE_X6Y134_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X6Y134_BO5),
.Q(CLBLM_R_X5Y134_SLICE_X6Y134_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y133_SLICE_X6Y133_CO6),
.Q(CLBLM_R_X5Y134_SLICE_X6Y134_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X6Y134_AO6),
.Q(CLBLM_R_X5Y134_SLICE_X6Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X6Y134_BO6),
.Q(CLBLM_R_X5Y134_SLICE_X6Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X6Y134_CO6),
.Q(CLBLM_R_X5Y134_SLICE_X6Y134_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X6Y134_DO6),
.Q(CLBLM_R_X5Y134_SLICE_X6Y134_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heffefefe45545454)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y130_SLICE_X7Y130_DQ),
.I2(CLBLM_R_X5Y134_SLICE_X6Y134_DQ),
.I3(CLBLM_R_X5Y135_SLICE_X6Y135_CO6),
.I4(CLBLM_R_X5Y132_SLICE_X6Y132_AQ),
.I5(CLBLM_R_X5Y133_SLICE_X7Y133_BQ),
.O5(CLBLM_R_X5Y134_SLICE_X6Y134_DO5),
.O6(CLBLM_R_X5Y134_SLICE_X6Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00eeeedddd)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_CLUT (
.I0(CLBLM_R_X5Y134_SLICE_X6Y134_CQ),
.I1(CLBLM_R_X5Y130_SLICE_X7Y130_DQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y133_SLICE_X4Y133_A5Q),
.I4(CLBLM_R_X5Y137_SLICE_X6Y137_DO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y134_SLICE_X6Y134_CO5),
.O6(CLBLM_R_X5Y134_SLICE_X6Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afa0fcfc0c0c)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_BLUT (
.I0(CLBLM_R_X7Y142_SLICE_X9Y142_CQ),
.I1(CLBLL_L_X4Y131_SLICE_X4Y131_D5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y133_SLICE_X6Y133_B5Q),
.I4(CLBLM_R_X7Y137_SLICE_X8Y137_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X6Y134_BO5),
.O6(CLBLM_R_X5Y134_SLICE_X6Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0f000fcc0fcc0f)
  ) CLBLM_R_X5Y134_SLICE_X6Y134_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y132_SLICE_X12Y132_AQ),
.I2(CLBLM_R_X11Y142_SLICE_X14Y142_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y135_SLICE_X4Y135_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X6Y134_AO5),
.O6(CLBLM_R_X5Y134_SLICE_X6Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X7Y134_AO5),
.Q(CLBLM_R_X5Y134_SLICE_X7Y134_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X7Y134_DO5),
.Q(CLBLM_R_X5Y134_SLICE_X7Y134_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X7Y134_AO6),
.Q(CLBLM_R_X5Y134_SLICE_X7Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X7Y134_BO6),
.Q(CLBLM_R_X5Y134_SLICE_X7Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X7Y134_CO6),
.Q(CLBLM_R_X5Y134_SLICE_X7Y134_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y134_SLICE_X7Y134_DO6),
.Q(CLBLM_R_X5Y134_SLICE_X7Y134_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888ee44ee44)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y141_SLICE_X8Y141_A5Q),
.I2(1'b1),
.I3(CLBLM_L_X10Y133_SLICE_X13Y133_AQ),
.I4(CLBLM_R_X5Y134_SLICE_X6Y134_DQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X7Y134_DO5),
.O6(CLBLM_R_X5Y134_SLICE_X7Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaffffcccc)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_CLUT (
.I0(CLBLL_L_X4Y132_SLICE_X5Y132_C5Q),
.I1(CLBLM_L_X8Y134_SLICE_X10Y134_BO6),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_L_X8Y139_SLICE_X11Y139_BQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y134_SLICE_X7Y134_CO5),
.O6(CLBLM_R_X5Y134_SLICE_X7Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f1f1ff00f1f1)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_BLUT (
.I0(CLBLL_L_X4Y134_SLICE_X5Y134_CQ),
.I1(CLBLM_R_X5Y134_SLICE_X7Y134_BQ),
.I2(CLBLL_L_X4Y139_SLICE_X5Y139_CQ),
.I3(CLBLM_L_X8Y133_SLICE_X10Y133_C5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X7Y134_BO5),
.O6(CLBLM_R_X5Y134_SLICE_X7Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa33aa33f055f0aa)
  ) CLBLM_R_X5Y134_SLICE_X7Y134_ALUT (
.I0(CLBLM_R_X5Y134_SLICE_X6Y134_DQ),
.I1(CLBLM_L_X10Y140_SLICE_X13Y140_BQ),
.I2(CLBLL_L_X4Y131_SLICE_X5Y131_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y134_SLICE_X7Y134_AO5),
.O6(CLBLM_R_X5Y134_SLICE_X7Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y135_SLICE_X6Y135_AO5),
.Q(CLBLM_R_X5Y135_SLICE_X6Y135_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y135_SLICE_X6Y135_BO5),
.Q(CLBLM_R_X5Y135_SLICE_X6Y135_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y135_SLICE_X6Y135_AO6),
.Q(CLBLM_R_X5Y135_SLICE_X6Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y135_SLICE_X6Y135_BO6),
.Q(CLBLM_R_X5Y135_SLICE_X6Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha000a000a000a000)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_DLUT (
.I0(CLBLL_L_X4Y137_SLICE_X5Y137_C5Q),
.I1(1'b1),
.I2(CLBLL_L_X4Y138_SLICE_X5Y138_DQ),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y135_SLICE_X6Y135_DO5),
.O6(CLBLM_R_X5Y135_SLICE_X6Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h800000006aaaaaaa)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_CLUT (
.I0(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.I1(CLBLM_R_X3Y135_SLICE_X3Y135_BQ),
.I2(CLBLM_R_X5Y134_SLICE_X6Y134_CQ),
.I3(CLBLM_R_X3Y135_SLICE_X3Y135_CQ),
.I4(CLBLM_R_X5Y135_SLICE_X6Y135_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y135_SLICE_X6Y135_CO5),
.O6(CLBLM_R_X5Y135_SLICE_X6Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc3030b8b8b8b8)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_BLUT (
.I0(CLBLL_L_X4Y134_SLICE_X5Y134_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y135_SLICE_X10Y135_DQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y135_SLICE_X6Y135_BO5),
.O6(CLBLM_R_X5Y135_SLICE_X6Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33cc00b8b8b8b8)
  ) CLBLM_R_X5Y135_SLICE_X6Y135_ALUT (
.I0(CLBLL_L_X4Y135_SLICE_X4Y135_CQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y137_SLICE_X9Y137_D5Q),
.I3(CLBLM_R_X5Y135_SLICE_X7Y135_BQ),
.I4(CLBLM_R_X3Y135_SLICE_X3Y135_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y135_SLICE_X6Y135_AO5),
.O6(CLBLM_R_X5Y135_SLICE_X6Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y135_SLICE_X7Y135_BO5),
.Q(CLBLM_R_X5Y135_SLICE_X7Y135_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y135_SLICE_X7Y135_DO5),
.Q(CLBLM_R_X5Y135_SLICE_X7Y135_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y135_SLICE_X7Y135_AO6),
.Q(CLBLM_R_X5Y135_SLICE_X7Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y135_SLICE_X7Y135_BO6),
.Q(CLBLM_R_X5Y135_SLICE_X7Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y135_SLICE_X7Y135_CO6),
.Q(CLBLM_R_X5Y135_SLICE_X7Y135_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y135_SLICE_X7Y135_DO6),
.Q(CLBLM_R_X5Y135_SLICE_X7Y135_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff003c3caaaacccc)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_DLUT (
.I0(CLBLM_R_X5Y139_SLICE_X7Y139_AQ),
.I1(CLBLL_L_X4Y137_SLICE_X5Y137_C5Q),
.I2(CLBLL_L_X4Y132_SLICE_X5Y132_D5Q),
.I3(CLBLM_R_X7Y132_SLICE_X8Y132_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y135_SLICE_X7Y135_DO5),
.O6(CLBLM_R_X5Y135_SLICE_X7Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccf000faaa)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_CLUT (
.I0(CLBLM_R_X5Y139_SLICE_X7Y139_B5Q),
.I1(CLBLM_L_X8Y135_SLICE_X10Y135_AQ),
.I2(CLBLL_L_X4Y136_SLICE_X4Y136_AQ),
.I3(CLBLL_L_X4Y136_SLICE_X4Y136_CQ),
.I4(CLBLM_R_X11Y140_SLICE_X15Y140_CO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y135_SLICE_X7Y135_CO5),
.O6(CLBLM_R_X5Y135_SLICE_X7Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0fcc0faa0faa0f)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_BLUT (
.I0(CLBLM_R_X3Y137_SLICE_X3Y137_A5Q),
.I1(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.I2(CLBLL_L_X4Y131_SLICE_X5Y131_B5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y135_SLICE_X7Y135_BO5),
.O6(CLBLM_R_X5Y135_SLICE_X7Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heefc2230eefc2230)
  ) CLBLM_R_X5Y135_SLICE_X7Y135_ALUT (
.I0(CLBLM_R_X5Y131_SLICE_X7Y131_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y135_SLICE_X7Y135_AQ),
.I3(CLBLM_R_X11Y131_SLICE_X14Y131_BO6),
.I4(CLBLM_R_X5Y135_SLICE_X6Y135_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y135_SLICE_X7Y135_AO5),
.O6(CLBLM_R_X5Y135_SLICE_X7Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X6Y136_BO5),
.Q(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X6Y136_AO6),
.Q(CLBLM_R_X5Y136_SLICE_X6Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X6Y136_BO6),
.Q(CLBLM_R_X5Y136_SLICE_X6Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X6Y136_CO6),
.Q(CLBLM_R_X5Y136_SLICE_X6Y136_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X6Y136_DO6),
.Q(CLBLM_R_X5Y136_SLICE_X6Y136_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88ddd88d88)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y136_SLICE_X6Y136_CQ),
.I2(CLBLM_R_X3Y136_SLICE_X2Y136_CQ),
.I3(CLBLL_L_X4Y136_SLICE_X4Y136_B5Q),
.I4(CLBLL_L_X4Y134_SLICE_X4Y134_C5Q),
.I5(CLBLL_L_X4Y135_SLICE_X4Y135_AQ),
.O5(CLBLM_R_X5Y136_SLICE_X6Y136_DO5),
.O6(CLBLM_R_X5Y136_SLICE_X6Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe54ae04fe54ae04)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y134_SLICE_X4Y134_BQ),
.I2(CLBLM_L_X12Y132_SLICE_X16Y132_AO6),
.I3(CLBLM_R_X7Y135_SLICE_X9Y135_BQ),
.I4(CLBLM_R_X5Y136_SLICE_X6Y136_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y136_SLICE_X6Y136_CO5),
.O6(CLBLM_R_X5Y136_SLICE_X6Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888bbbbcc00ff33)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_BLUT (
.I0(CLBLM_R_X5Y141_SLICE_X6Y141_DQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLL_L_X4Y133_SLICE_X4Y133_CQ),
.I4(CLBLM_L_X10Y140_SLICE_X13Y140_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y136_SLICE_X6Y136_BO5),
.O6(CLBLM_R_X5Y136_SLICE_X6Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00aaf0aaf0)
  ) CLBLM_R_X5Y136_SLICE_X6Y136_ALUT (
.I0(CLBLM_R_X5Y134_SLICE_X6Y134_B5Q),
.I1(1'b1),
.I2(CLBLM_R_X5Y136_SLICE_X6Y136_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y136_SLICE_X7Y136_AQ),
.I5(CLBLM_R_X11Y131_SLICE_X14Y131_BO6),
.O5(CLBLM_R_X5Y136_SLICE_X6Y136_AO5),
.O6(CLBLM_R_X5Y136_SLICE_X6Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X7Y136_CO5),
.Q(CLBLM_R_X5Y136_SLICE_X7Y136_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X7Y136_DO5),
.Q(CLBLM_R_X5Y136_SLICE_X7Y136_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X7Y136_AO6),
.Q(CLBLM_R_X5Y136_SLICE_X7Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X7Y136_BO6),
.Q(CLBLM_R_X5Y136_SLICE_X7Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X7Y136_CO6),
.Q(CLBLM_R_X5Y136_SLICE_X7Y136_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y136_SLICE_X7Y136_DO6),
.Q(CLBLM_R_X5Y136_SLICE_X7Y136_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa50ffaa5500)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(CLBLL_L_X4Y136_SLICE_X5Y136_DQ),
.I3(CLBLM_R_X3Y141_SLICE_X2Y141_BQ),
.I4(CLBLM_R_X7Y136_SLICE_X8Y136_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y136_SLICE_X7Y136_DO5),
.O6(CLBLM_R_X5Y136_SLICE_X7Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0dddd8888)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y136_SLICE_X9Y136_CQ),
.I2(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.I3(CLBLM_R_X5Y134_SLICE_X7Y134_CQ),
.I4(RIOB33_X105Y117_IOB_X1Y117_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y136_SLICE_X7Y136_CO5),
.O6(CLBLM_R_X5Y136_SLICE_X7Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfafcfc0c0a0c0c)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_BLUT (
.I0(CLBLM_R_X7Y136_SLICE_X8Y136_CQ),
.I1(CLBLM_R_X5Y136_SLICE_X7Y136_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y135_SLICE_X9Y135_C5Q),
.I4(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.I5(CLBLM_R_X11Y136_SLICE_X15Y136_AQ),
.O5(CLBLM_R_X5Y136_SLICE_X7Y136_BO5),
.O6(CLBLM_R_X5Y136_SLICE_X7Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefeaafe54540054)
  ) CLBLM_R_X5Y136_SLICE_X7Y136_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y133_SLICE_X8Y133_CQ),
.I2(CLBLM_R_X5Y136_SLICE_X7Y136_AQ),
.I3(CLBLL_L_X4Y135_SLICE_X4Y135_D5Q),
.I4(CLBLM_R_X5Y133_SLICE_X7Y133_AQ),
.I5(CLBLL_L_X4Y142_SLICE_X4Y142_A5Q),
.O5(CLBLM_R_X5Y136_SLICE_X7Y136_AO5),
.O6(CLBLM_R_X5Y136_SLICE_X7Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y137_SLICE_X6Y137_AO6),
.Q(CLBLM_R_X5Y137_SLICE_X6Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y137_SLICE_X6Y137_BO6),
.Q(CLBLM_R_X5Y137_SLICE_X6Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y137_SLICE_X6Y137_CO6),
.Q(CLBLM_R_X5Y137_SLICE_X6Y137_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffff7f7f7f7f)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_DLUT (
.I0(CLBLM_R_X3Y135_SLICE_X3Y135_CQ),
.I1(CLBLM_R_X3Y135_SLICE_X3Y135_BQ),
.I2(CLBLL_L_X4Y138_SLICE_X5Y138_DQ),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_BQ),
.I4(CLBLL_L_X4Y137_SLICE_X5Y137_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y137_SLICE_X6Y137_DO5),
.O6(CLBLM_R_X5Y137_SLICE_X6Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfa50ccccff00)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_CLUT (
.I0(CLBLL_L_X4Y135_SLICE_X4Y135_AQ),
.I1(CLBLM_R_X7Y137_SLICE_X8Y137_C5Q),
.I2(CLBLM_L_X12Y136_SLICE_X16Y136_A5Q),
.I3(CLBLM_R_X5Y136_SLICE_X6Y136_DQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X3Y136_SLICE_X2Y136_CQ),
.O5(CLBLM_R_X5Y137_SLICE_X6Y137_CO5),
.O6(CLBLM_R_X5Y137_SLICE_X6Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd888d8ddd88dd88)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.I2(CLBLL_L_X4Y131_SLICE_X5Y131_B5Q),
.I3(CLBLM_R_X5Y137_SLICE_X6Y137_CQ),
.I4(CLBLL_L_X4Y135_SLICE_X4Y135_AQ),
.I5(CLBLM_R_X3Y136_SLICE_X2Y136_CQ),
.O5(CLBLM_R_X5Y137_SLICE_X6Y137_BO5),
.O6(CLBLM_R_X5Y137_SLICE_X6Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cf404fc0cfe0e)
  ) CLBLM_R_X5Y137_SLICE_X6Y137_ALUT (
.I0(CLBLM_R_X3Y136_SLICE_X2Y136_CQ),
.I1(CLBLM_R_X5Y137_SLICE_X6Y137_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y134_SLICE_X5Y134_CQ),
.I4(CLBLL_L_X4Y135_SLICE_X4Y135_AQ),
.I5(CLBLM_R_X11Y142_SLICE_X14Y142_AQ),
.O5(CLBLM_R_X5Y137_SLICE_X6Y137_AO5),
.O6(CLBLM_R_X5Y137_SLICE_X6Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y137_SLICE_X7Y137_AO5),
.Q(CLBLM_R_X5Y137_SLICE_X7Y137_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y137_SLICE_X7Y137_BO5),
.Q(CLBLM_R_X5Y137_SLICE_X7Y137_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y137_SLICE_X7Y137_AO6),
.Q(CLBLM_R_X5Y137_SLICE_X7Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y137_SLICE_X7Y137_BO6),
.Q(CLBLM_R_X5Y137_SLICE_X7Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffaa)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_DLUT (
.I0(CLBLM_L_X8Y137_SLICE_X10Y137_CQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X3Y141_SLICE_X2Y141_BQ),
.I4(CLBLL_L_X4Y132_SLICE_X5Y132_C5Q),
.I5(CLBLM_R_X5Y136_SLICE_X7Y136_D5Q),
.O5(CLBLM_R_X5Y137_SLICE_X7Y137_DO5),
.O6(CLBLM_R_X5Y137_SLICE_X7Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffaa)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_CLUT (
.I0(CLBLM_R_X5Y134_SLICE_X7Y134_A5Q),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X7Y138_SLICE_X8Y138_DQ),
.I4(CLBLM_R_X5Y135_SLICE_X7Y135_DQ),
.I5(CLBLM_R_X7Y133_SLICE_X9Y133_BQ),
.O5(CLBLM_R_X5Y137_SLICE_X7Y137_CO5),
.O6(CLBLM_R_X5Y137_SLICE_X7Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0a0afc0cfc0c)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_BLUT (
.I0(CLBLL_L_X4Y137_SLICE_X4Y137_DO6),
.I1(CLBLM_L_X8Y139_SLICE_X10Y139_AO6),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y136_SLICE_X7Y136_D5Q),
.I4(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y137_SLICE_X7Y137_BO5),
.O6(CLBLM_R_X5Y137_SLICE_X7Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0eeee4444)
  ) CLBLM_R_X5Y137_SLICE_X7Y137_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y137_SLICE_X8Y137_D5Q),
.I2(CLBLL_L_X4Y140_SLICE_X5Y140_AQ),
.I3(CLBLL_L_X4Y134_SLICE_X4Y134_C5Q),
.I4(CLBLM_L_X8Y137_SLICE_X10Y137_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y137_SLICE_X7Y137_AO5),
.O6(CLBLM_R_X5Y137_SLICE_X7Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y138_SLICE_X6Y138_BO5),
.Q(CLBLM_R_X5Y138_SLICE_X6Y138_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y138_SLICE_X6Y138_AO6),
.Q(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y138_SLICE_X6Y138_BO6),
.Q(CLBLM_R_X5Y138_SLICE_X6Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y138_SLICE_X6Y138_CO6),
.Q(CLBLM_R_X5Y138_SLICE_X6Y138_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f00100cc00cc00)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_DLUT (
.I0(CLBLM_R_X5Y137_SLICE_X6Y137_DO5),
.I1(CLBLL_L_X4Y137_SLICE_X5Y137_C5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_BQ),
.I4(CLBLM_R_X5Y137_SLICE_X6Y137_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y138_SLICE_X6Y138_DO5),
.O6(CLBLM_R_X5Y138_SLICE_X6Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b888b8b8b8bbb8)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_CLUT (
.I0(CLBLM_R_X5Y140_SLICE_X6Y140_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y137_SLICE_X6Y137_AQ),
.I3(CLBLM_R_X3Y136_SLICE_X2Y136_CQ),
.I4(CLBLL_L_X4Y135_SLICE_X4Y135_AQ),
.I5(CLBLM_L_X10Y140_SLICE_X13Y140_BQ),
.O5(CLBLM_R_X5Y138_SLICE_X6Y138_CO5),
.O6(CLBLM_R_X5Y138_SLICE_X6Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa3caa3cccffcc00)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_BLUT (
.I0(CLBLM_L_X8Y140_SLICE_X10Y140_DQ),
.I1(CLBLM_R_X7Y130_SLICE_X9Y130_BQ),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X2Y138_SLICE_X1Y138_BO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y138_SLICE_X6Y138_BO5),
.O6(CLBLM_R_X5Y138_SLICE_X6Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0cc00ccf5cc00)
  ) CLBLM_R_X5Y138_SLICE_X6Y138_ALUT (
.I0(CLBLM_R_X5Y139_SLICE_X7Y139_CQ),
.I1(CLBLM_R_X7Y133_SLICE_X9Y133_CQ),
.I2(CLBLM_R_X5Y138_SLICE_X7Y138_DO6),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.I5(CLBLL_L_X4Y138_SLICE_X5Y138_B5Q),
.O5(CLBLM_R_X5Y138_SLICE_X6Y138_AO5),
.O6(CLBLM_R_X5Y138_SLICE_X6Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y138_SLICE_X7Y138_AO6),
.Q(CLBLM_R_X5Y138_SLICE_X7Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbfffffffffff)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_DLUT (
.I0(CLBLM_R_X3Y135_SLICE_X3Y135_DQ),
.I1(CLBLM_R_X5Y140_SLICE_X6Y140_CQ),
.I2(CLBLM_R_X7Y138_SLICE_X9Y138_B5Q),
.I3(CLBLM_R_X5Y134_SLICE_X6Y134_DQ),
.I4(CLBLM_R_X5Y138_SLICE_X7Y138_BO5),
.I5(CLBLM_R_X5Y137_SLICE_X7Y137_BQ),
.O5(CLBLM_R_X5Y138_SLICE_X7Y138_DO5),
.O6(CLBLM_R_X5Y138_SLICE_X7Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffff7fff)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_CLUT (
.I0(CLBLM_R_X7Y130_SLICE_X9Y130_BQ),
.I1(CLBLL_L_X4Y137_SLICE_X5Y137_C5Q),
.I2(CLBLM_R_X5Y134_SLICE_X6Y134_DQ),
.I3(CLBLM_R_X5Y140_SLICE_X6Y140_CQ),
.I4(CLBLM_R_X5Y138_SLICE_X7Y138_BO5),
.I5(CLBLM_R_X5Y137_SLICE_X6Y137_DO5),
.O5(CLBLM_R_X5Y138_SLICE_X7Y138_CO5),
.O6(CLBLM_R_X5Y138_SLICE_X7Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffee5fff5fff)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_BLUT (
.I0(CLBLM_R_X5Y132_SLICE_X6Y132_AQ),
.I1(CLBLM_R_X5Y137_SLICE_X7Y137_BQ),
.I2(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.I3(CLBLM_R_X5Y134_SLICE_X6Y134_CQ),
.I4(CLBLM_R_X7Y138_SLICE_X9Y138_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y138_SLICE_X7Y138_BO5),
.O6(CLBLM_R_X5Y138_SLICE_X7Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ee22ff33ff33)
  ) CLBLM_R_X5Y138_SLICE_X7Y138_ALUT (
.I0(CLBLM_R_X5Y138_SLICE_X7Y138_DO6),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLM_L_X8Y137_SLICE_X10Y137_C5Q),
.I4(1'b1),
.I5(CLBLM_R_X5Y139_SLICE_X7Y139_CQ),
.O5(CLBLM_R_X5Y138_SLICE_X7Y138_AO5),
.O6(CLBLM_R_X5Y138_SLICE_X7Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y139_SLICE_X6Y139_CO5),
.Q(CLBLM_R_X5Y139_SLICE_X6Y139_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y139_SLICE_X6Y139_AO6),
.Q(CLBLM_R_X5Y139_SLICE_X6Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y139_SLICE_X6Y139_BO6),
.Q(CLBLM_R_X5Y139_SLICE_X6Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y139_SLICE_X6Y139_CO6),
.Q(CLBLM_R_X5Y139_SLICE_X6Y139_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a2a0a2a0a2a0a2)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_DLUT (
.I0(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.I1(CLBLL_L_X4Y138_SLICE_X5Y138_B5Q),
.I2(CLBLM_R_X5Y138_SLICE_X7Y138_DO6),
.I3(CLBLM_R_X5Y139_SLICE_X7Y139_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y139_SLICE_X6Y139_DO5),
.O6(CLBLM_R_X5Y139_SLICE_X6Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacacacc0cfcfc0)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_CLUT (
.I0(CLBLM_R_X5Y140_SLICE_X7Y140_AQ),
.I1(CLBLL_L_X4Y130_SLICE_X5Y130_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y132_SLICE_X6Y132_AQ),
.I4(CLBLM_R_X7Y140_SLICE_X8Y140_DQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y139_SLICE_X6Y139_CO5),
.O6(CLBLM_R_X5Y139_SLICE_X6Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00bbbbbbbb)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_BLUT (
.I0(CLBLM_R_X5Y139_SLICE_X6Y139_DO6),
.I1(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y136_SLICE_X9Y136_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y139_SLICE_X6Y139_BO5),
.O6(CLBLM_R_X5Y139_SLICE_X6Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8bbb8bbb888b888)
  ) CLBLM_R_X5Y139_SLICE_X6Y139_ALUT (
.I0(CLBLM_R_X11Y140_SLICE_X15Y140_BQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y139_SLICE_X6Y139_AQ),
.I3(CLBLM_L_X12Y132_SLICE_X16Y132_AO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y139_SLICE_X5Y139_AQ),
.O5(CLBLM_R_X5Y139_SLICE_X6Y139_AO5),
.O6(CLBLM_R_X5Y139_SLICE_X6Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y139_SLICE_X7Y139_AO5),
.Q(CLBLM_R_X5Y139_SLICE_X7Y139_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y139_SLICE_X7Y139_BO5),
.Q(CLBLM_R_X5Y139_SLICE_X7Y139_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y139_SLICE_X7Y139_AO6),
.Q(CLBLM_R_X5Y139_SLICE_X7Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y139_SLICE_X7Y139_BO6),
.Q(CLBLM_R_X5Y139_SLICE_X7Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y139_SLICE_X7Y139_CO6),
.Q(CLBLM_R_X5Y139_SLICE_X7Y139_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_DLUT (
.I0(CLBLM_R_X5Y140_SLICE_X7Y140_AQ),
.I1(CLBLM_R_X7Y140_SLICE_X8Y140_B5Q),
.I2(CLBLM_L_X8Y133_SLICE_X11Y133_BQ),
.I3(CLBLM_R_X3Y136_SLICE_X3Y136_CQ),
.I4(CLBLM_R_X7Y139_SLICE_X8Y139_CO6),
.I5(CLBLM_R_X5Y139_SLICE_X6Y139_C5Q),
.O5(CLBLM_R_X5Y139_SLICE_X7Y139_DO5),
.O6(CLBLM_R_X5Y139_SLICE_X7Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000440044)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_CLUT (
.I0(CLBLM_R_X5Y137_SLICE_X6Y137_DO5),
.I1(CLBLL_L_X4Y137_SLICE_X5Y137_C5Q),
.I2(1'b1),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_BQ),
.I4(CLBLM_R_X5Y137_SLICE_X7Y137_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y139_SLICE_X7Y139_CO5),
.O6(CLBLM_R_X5Y139_SLICE_X7Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0fafa0a0a)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_BLUT (
.I0(CLBLM_R_X3Y139_SLICE_X3Y139_DO6),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_C5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y136_SLICE_X8Y136_C5Q),
.I4(CLBLM_R_X5Y138_SLICE_X6Y138_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y139_SLICE_X7Y139_BO5),
.O6(CLBLM_R_X5Y139_SLICE_X7Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afa0c0cfcfc0)
  ) CLBLM_R_X5Y139_SLICE_X7Y139_ALUT (
.I0(CLBLM_R_X3Y136_SLICE_X2Y136_B5Q),
.I1(CLBLM_L_X8Y140_SLICE_X11Y140_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y137_SLICE_X7Y137_BQ),
.I4(CLBLM_L_X8Y131_SLICE_X11Y131_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y139_SLICE_X7Y139_AO5),
.O6(CLBLM_R_X5Y139_SLICE_X7Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y140_SLICE_X6Y140_BO6),
.Q(CLBLM_R_X5Y140_SLICE_X6Y140_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y140_SLICE_X6Y140_AO6),
.Q(CLBLM_R_X5Y140_SLICE_X6Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y140_SLICE_X6Y140_CO6),
.Q(CLBLM_R_X5Y140_SLICE_X6Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y140_SLICE_X6Y140_DO5),
.O6(CLBLM_R_X5Y140_SLICE_X6Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbebe0000bebe)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_CLUT (
.I0(CLBLM_R_X5Y130_SLICE_X7Y130_DQ),
.I1(CLBLM_R_X5Y140_SLICE_X6Y140_CQ),
.I2(CLBLM_R_X5Y140_SLICE_X7Y140_DO6),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y141_SLICE_X6Y141_BQ),
.O5(CLBLM_R_X5Y140_SLICE_X6Y140_CO5),
.O6(CLBLM_R_X5Y140_SLICE_X6Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0e4a0e4fffff0f0)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y139_SLICE_X7Y139_DO6),
.I2(CLBLM_R_X5Y131_SLICE_X6Y131_BQ),
.I3(CLBLM_R_X5Y137_SLICE_X7Y137_CO6),
.I4(CLBLM_L_X10Y137_SLICE_X13Y137_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y140_SLICE_X6Y140_BO5),
.O6(CLBLM_R_X5Y140_SLICE_X6Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa800a8fffc00fc)
  ) CLBLM_R_X5Y140_SLICE_X6Y140_ALUT (
.I0(CLBLM_R_X5Y133_SLICE_X7Y133_AQ),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_DQ),
.I2(CLBLM_R_X5Y140_SLICE_X6Y140_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y139_SLICE_X5Y139_C5Q),
.I5(CLBLL_L_X4Y135_SLICE_X4Y135_D5Q),
.O5(CLBLM_R_X5Y140_SLICE_X6Y140_AO5),
.O6(CLBLM_R_X5Y140_SLICE_X6Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y140_SLICE_X7Y140_AO5),
.Q(CLBLM_R_X5Y140_SLICE_X7Y140_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y140_SLICE_X7Y140_BO5),
.Q(CLBLM_R_X5Y140_SLICE_X7Y140_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y140_SLICE_X7Y140_AO6),
.Q(CLBLM_R_X5Y140_SLICE_X7Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y140_SLICE_X7Y140_BO6),
.Q(CLBLM_R_X5Y140_SLICE_X7Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y140_SLICE_X7Y140_CO6),
.Q(CLBLM_R_X5Y140_SLICE_X7Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000080800000000)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_DLUT (
.I0(CLBLL_L_X4Y137_SLICE_X5Y137_C5Q),
.I1(CLBLM_R_X7Y130_SLICE_X9Y130_BQ),
.I2(CLBLM_R_X5Y137_SLICE_X6Y137_DO5),
.I3(1'b1),
.I4(CLBLM_R_X5Y138_SLICE_X7Y138_BO5),
.I5(CLBLM_R_X5Y134_SLICE_X6Y134_DQ),
.O5(CLBLM_R_X5Y140_SLICE_X7Y140_DO5),
.O6(CLBLM_R_X5Y140_SLICE_X7Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0c0c5c0c5)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_CLUT (
.I0(CLBLL_L_X4Y137_SLICE_X5Y137_C5Q),
.I1(CLBLM_R_X5Y135_SLICE_X7Y135_D5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_BQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y137_SLICE_X6Y137_DO5),
.O5(CLBLM_R_X5Y140_SLICE_X7Y140_CO5),
.O6(CLBLM_R_X5Y140_SLICE_X7Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33cc00efef2323)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_BLUT (
.I0(CLBLM_R_X5Y138_SLICE_X7Y138_DO6),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y140_SLICE_X7Y140_CQ),
.I3(CLBLL_L_X4Y142_SLICE_X5Y142_A5Q),
.I4(CLBLM_L_X10Y134_SLICE_X12Y134_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y140_SLICE_X7Y140_BO5),
.O6(CLBLM_R_X5Y140_SLICE_X7Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5c5cacafc0cfc0c)
  ) CLBLM_R_X5Y140_SLICE_X7Y140_ALUT (
.I0(CLBLL_L_X4Y138_SLICE_X5Y138_DQ),
.I1(CLBLM_R_X5Y140_SLICE_X7Y140_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X3Y140_SLICE_X3Y140_DQ),
.I4(CLBLM_L_X10Y140_SLICE_X12Y140_DQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y140_SLICE_X7Y140_AO5),
.O6(CLBLM_R_X5Y140_SLICE_X7Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y141_SLICE_X6Y141_AO6),
.Q(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y141_SLICE_X6Y141_BO6),
.Q(CLBLM_R_X5Y141_SLICE_X6Y141_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y141_SLICE_X6Y141_CO6),
.Q(CLBLM_R_X5Y141_SLICE_X6Y141_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y141_SLICE_X6Y141_DO6),
.Q(CLBLM_R_X5Y141_SLICE_X6Y141_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff480048ffc000c0)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_DLUT (
.I0(CLBLL_L_X4Y140_SLICE_X4Y140_BO5),
.I1(CLBLM_R_X5Y141_SLICE_X7Y141_AO6),
.I2(CLBLM_R_X5Y141_SLICE_X6Y141_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y140_SLICE_X8Y140_CQ),
.I5(CLBLL_L_X4Y142_SLICE_X5Y142_A5Q),
.O5(CLBLM_R_X5Y141_SLICE_X6Y141_DO5),
.O6(CLBLM_R_X5Y141_SLICE_X6Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0001010303)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_CLUT (
.I0(CLBLM_R_X5Y141_SLICE_X6Y141_BQ),
.I1(CLBLM_R_X5Y139_SLICE_X7Y139_BQ),
.I2(CLBLM_R_X5Y142_SLICE_X6Y142_BQ),
.I3(CLBLM_L_X8Y142_SLICE_X10Y142_A5Q),
.I4(CLBLM_R_X5Y141_SLICE_X6Y141_CQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y141_SLICE_X6Y141_CO5),
.O6(CLBLM_R_X5Y141_SLICE_X6Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcfcfcfcacfca)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_BLUT (
.I0(CLBLM_R_X5Y141_SLICE_X6Y141_CQ),
.I1(CLBLM_L_X10Y140_SLICE_X13Y140_DQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y139_SLICE_X7Y139_BQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y142_SLICE_X6Y142_BQ),
.O5(CLBLM_R_X5Y141_SLICE_X6Y141_BO5),
.O6(CLBLM_R_X5Y141_SLICE_X6Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccaaccffccff)
  ) CLBLM_R_X5Y141_SLICE_X6Y141_ALUT (
.I0(CLBLM_R_X5Y138_SLICE_X7Y138_DO6),
.I1(CLBLM_R_X5Y142_SLICE_X6Y142_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y138_SLICE_X5Y138_B5Q),
.O5(CLBLM_R_X5Y141_SLICE_X6Y141_AO5),
.O6(CLBLM_R_X5Y141_SLICE_X6Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdcdcdcdcfcfcfcfc)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_DLUT (
.I0(CLBLM_R_X5Y143_SLICE_X7Y143_AQ),
.I1(CLBLL_L_X4Y143_SLICE_X5Y143_DO6),
.I2(CLBLM_L_X10Y137_SLICE_X12Y137_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y142_SLICE_X5Y142_A5Q),
.O5(CLBLM_R_X5Y141_SLICE_X7Y141_DO5),
.O6(CLBLM_R_X5Y141_SLICE_X7Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffeffffff)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_CLUT (
.I0(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.I1(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.I2(CLBLM_R_X11Y139_SLICE_X14Y139_AO5),
.I3(CLBLL_L_X4Y142_SLICE_X5Y142_A5Q),
.I4(CLBLM_R_X5Y141_SLICE_X6Y141_DQ),
.I5(CLBLL_L_X4Y140_SLICE_X4Y140_CO5),
.O5(CLBLM_R_X5Y141_SLICE_X7Y141_CO5),
.O6(CLBLM_R_X5Y141_SLICE_X7Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4455000040500000)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_BLUT (
.I0(CLBLM_R_X5Y141_SLICE_X7Y141_DO6),
.I1(CLBLM_R_X3Y135_SLICE_X2Y135_AQ),
.I2(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.I3(CLBLM_L_X8Y136_SLICE_X10Y136_BQ),
.I4(CLBLL_L_X4Y140_SLICE_X4Y140_BO5),
.I5(CLBLM_L_X10Y137_SLICE_X12Y137_AQ),
.O5(CLBLM_R_X5Y141_SLICE_X7Y141_BO5),
.O6(CLBLM_R_X5Y141_SLICE_X7Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00fd00f70a0a0a0a)
  ) CLBLM_R_X5Y141_SLICE_X7Y141_ALUT (
.I0(CLBLM_L_X8Y136_SLICE_X10Y136_BQ),
.I1(CLBLM_R_X7Y141_SLICE_X9Y141_A5Q),
.I2(CLBLM_R_X3Y135_SLICE_X2Y135_AQ),
.I3(CLBLM_R_X5Y141_SLICE_X7Y141_BO6),
.I4(CLBLM_L_X10Y130_SLICE_X12Y130_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y141_SLICE_X7Y141_AO5),
.O6(CLBLM_R_X5Y141_SLICE_X7Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X6Y142_BO5),
.Q(CLBLM_R_X5Y142_SLICE_X6Y142_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X6Y142_AO6),
.Q(CLBLM_R_X5Y142_SLICE_X6Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X6Y142_BO6),
.Q(CLBLM_R_X5Y142_SLICE_X6Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X6Y142_CO6),
.Q(CLBLM_R_X5Y142_SLICE_X6Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y142_SLICE_X6Y142_DO5),
.O6(CLBLM_R_X5Y142_SLICE_X6Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff9cff00009c0000)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_CLUT (
.I0(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.I1(CLBLM_R_X5Y142_SLICE_X6Y142_CQ),
.I2(CLBLM_R_X5Y142_SLICE_X7Y142_BO6),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y141_SLICE_X7Y141_AO6),
.I5(CLBLM_R_X5Y130_SLICE_X6Y130_AQ),
.O5(CLBLM_R_X5Y142_SLICE_X6Y142_CO5),
.O6(CLBLM_R_X5Y142_SLICE_X6Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0f3f38888bbbb)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_BLUT (
.I0(CLBLL_L_X4Y143_SLICE_X5Y143_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y140_SLICE_X8Y140_DQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y139_SLICE_X5Y139_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y142_SLICE_X6Y142_BO5),
.O6(CLBLM_R_X5Y142_SLICE_X6Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddd88888ddd8ddd8)
  ) CLBLM_R_X5Y142_SLICE_X6Y142_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y142_SLICE_X10Y142_AQ),
.I2(CLBLM_R_X5Y142_SLICE_X6Y142_AQ),
.I3(CLBLM_R_X5Y135_SLICE_X6Y135_B5Q),
.I4(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I5(CLBLL_L_X4Y135_SLICE_X5Y135_CQ),
.O5(CLBLM_R_X5Y142_SLICE_X6Y142_AO5),
.O6(CLBLM_R_X5Y142_SLICE_X6Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y142_SLICE_X7Y142_AO6),
.Q(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y142_SLICE_X7Y142_DO5),
.O6(CLBLM_R_X5Y142_SLICE_X7Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y142_SLICE_X7Y142_CO5),
.O6(CLBLM_R_X5Y142_SLICE_X7Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000200055ffffff)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_BLUT (
.I0(CLBLM_R_X5Y141_SLICE_X6Y141_DQ),
.I1(CLBLL_L_X4Y140_SLICE_X4Y140_CO5),
.I2(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.I3(CLBLL_L_X4Y142_SLICE_X5Y142_A5Q),
.I4(CLBLL_L_X4Y140_SLICE_X4Y140_BO5),
.I5(1'b1),
.O5(CLBLM_R_X5Y142_SLICE_X7Y142_BO5),
.O6(CLBLM_R_X5Y142_SLICE_X7Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccca0f50000)
  ) CLBLM_R_X5Y142_SLICE_X7Y142_ALUT (
.I0(CLBLM_R_X5Y142_SLICE_X7Y142_BO5),
.I1(CLBLL_L_X4Y137_SLICE_X5Y137_A5Q),
.I2(CLBLM_R_X5Y142_SLICE_X7Y142_AQ),
.I3(CLBLM_R_X5Y142_SLICE_X7Y142_BO6),
.I4(CLBLM_R_X5Y141_SLICE_X7Y141_AO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X5Y142_SLICE_X7Y142_AO5),
.O6(CLBLM_R_X5Y142_SLICE_X7Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y143_SLICE_X6Y143_DO5),
.O6(CLBLM_R_X5Y143_SLICE_X6Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y143_SLICE_X6Y143_CO5),
.O6(CLBLM_R_X5Y143_SLICE_X6Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y143_SLICE_X6Y143_BO5),
.O6(CLBLM_R_X5Y143_SLICE_X6Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y143_SLICE_X6Y143_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y143_SLICE_X6Y143_AO5),
.O6(CLBLM_R_X5Y143_SLICE_X6Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y143_SLICE_X7Y143_AO6),
.Q(CLBLM_R_X5Y143_SLICE_X7Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y143_SLICE_X7Y143_DO5),
.O6(CLBLM_R_X5Y143_SLICE_X7Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y143_SLICE_X7Y143_CO5),
.O6(CLBLM_R_X5Y143_SLICE_X7Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y143_SLICE_X7Y143_BO5),
.O6(CLBLM_R_X5Y143_SLICE_X7Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcffccccc03300000)
  ) CLBLM_R_X5Y143_SLICE_X7Y143_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X5Y143_SLICE_X7Y143_AQ),
.I3(CLBLL_L_X4Y143_SLICE_X5Y143_CO6),
.I4(CLBLM_R_X5Y141_SLICE_X7Y141_AO6),
.I5(CLBLM_R_X7Y138_SLICE_X9Y138_BQ),
.O5(CLBLM_R_X5Y143_SLICE_X7Y143_AO5),
.O6(CLBLM_R_X5Y143_SLICE_X7Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X7Y134_SLICE_X8Y134_AQ),
.Q(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_DO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_CO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_BO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y129_SLICE_X8Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X8Y129_AO5),
.O6(CLBLM_R_X7Y129_SLICE_X8Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_DO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_CO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_BO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y129_SLICE_X9Y129_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y129_SLICE_X9Y129_AO5),
.O6(CLBLM_R_X7Y129_SLICE_X9Y129_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X8Y130_AO6),
.Q(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X8Y130_BO6),
.Q(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_DLUT (
.I0(CLBLM_R_X7Y134_SLICE_X9Y134_BQ),
.I1(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.I2(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.I3(CLBLM_R_X7Y138_SLICE_X8Y138_CQ),
.I4(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.I5(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.O5(CLBLM_R_X7Y130_SLICE_X8Y130_DO5),
.O6(CLBLM_R_X7Y130_SLICE_X8Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800000080000000)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_CLUT (
.I0(CLBLM_R_X7Y134_SLICE_X9Y134_BQ),
.I1(CLBLM_R_X7Y138_SLICE_X8Y138_CQ),
.I2(CLBLM_R_X5Y131_SLICE_X7Y131_BQ),
.I3(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I4(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y130_SLICE_X8Y130_CO5),
.O6(CLBLM_R_X7Y130_SLICE_X8Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaaf0f033cc)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_BLUT (
.I0(CLBLM_R_X7Y132_SLICE_X8Y132_DQ),
.I1(CLBLM_R_X7Y130_SLICE_X8Y130_BQ),
.I2(CLBLM_R_X5Y131_SLICE_X7Y131_CQ),
.I3(CLBLM_R_X7Y130_SLICE_X8Y130_DO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y133_SLICE_X6Y133_A5Q),
.O5(CLBLM_R_X7Y130_SLICE_X8Y130_BO5),
.O6(CLBLM_R_X7Y130_SLICE_X8Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaccaa0faaf0)
  ) CLBLM_R_X7Y130_SLICE_X8Y130_ALUT (
.I0(CLBLL_L_X4Y136_SLICE_X4Y136_A5Q),
.I1(CLBLM_L_X10Y135_SLICE_X12Y135_A5Q),
.I2(CLBLM_R_X7Y130_SLICE_X8Y130_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y130_SLICE_X8Y130_CO5),
.I5(CLBLM_R_X5Y133_SLICE_X6Y133_A5Q),
.O5(CLBLM_R_X7Y130_SLICE_X8Y130_AO5),
.O6(CLBLM_R_X7Y130_SLICE_X8Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X9Y130_AO6),
.Q(CLBLM_R_X7Y130_SLICE_X9Y130_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y130_SLICE_X9Y130_BO6),
.Q(CLBLM_R_X7Y130_SLICE_X9Y130_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y130_SLICE_X9Y130_DO5),
.O6(CLBLM_R_X7Y130_SLICE_X9Y130_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y130_SLICE_X9Y130_CO5),
.O6(CLBLM_R_X7Y130_SLICE_X9Y130_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff660000ff66)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_BLUT (
.I0(CLBLL_L_X4Y137_SLICE_X5Y137_C5Q),
.I1(CLBLM_R_X7Y130_SLICE_X9Y130_BQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y130_SLICE_X7Y130_DQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y131_SLICE_X8Y131_CQ),
.O5(CLBLM_R_X7Y130_SLICE_X9Y130_BO5),
.O6(CLBLM_R_X7Y130_SLICE_X9Y130_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff2ffd000f200d0)
  ) CLBLM_R_X7Y130_SLICE_X9Y130_ALUT (
.I0(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.I1(CLBLM_R_X7Y135_SLICE_X9Y135_C5Q),
.I2(CLBLM_R_X7Y130_SLICE_X9Y130_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y133_SLICE_X8Y133_AQ),
.I5(CLBLM_L_X10Y130_SLICE_X12Y130_C5Q),
.O5(CLBLM_R_X7Y130_SLICE_X9Y130_AO5),
.O6(CLBLM_R_X7Y130_SLICE_X9Y130_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X8Y131_BO6),
.Q(CLBLM_R_X7Y131_SLICE_X8Y131_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X8Y131_CO5),
.Q(CLBLM_R_X7Y131_SLICE_X8Y131_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X8Y131_AO6),
.Q(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X8Y131_CO6),
.Q(CLBLM_R_X7Y131_SLICE_X8Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X8Y131_DO6),
.Q(CLBLM_R_X7Y131_SLICE_X8Y131_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffa5550aafa0050)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(CLBLM_R_X7Y131_SLICE_X8Y131_DQ),
.I3(CLBLM_R_X13Y134_SLICE_X18Y134_AO6),
.I4(CLBLM_R_X7Y134_SLICE_X8Y134_A5Q),
.I5(CLBLM_R_X5Y142_SLICE_X6Y142_AQ),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_DO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefe5454f5a0f5a0)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y131_SLICE_X8Y131_CQ),
.I2(CLBLM_R_X7Y132_SLICE_X8Y132_D5Q),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(CLBLM_L_X8Y131_SLICE_X10Y131_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_CO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c5c0ca5555ffff)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_BLUT (
.I0(CLBLL_L_X4Y134_SLICE_X4Y134_CQ),
.I1(CLBLM_R_X7Y136_SLICE_X8Y136_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y130_SLICE_X6Y130_B5Q),
.I4(CLBLM_R_X7Y131_SLICE_X8Y131_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_BO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcced0021ccfc0030)
  ) CLBLM_R_X7Y131_SLICE_X8Y131_ALUT (
.I0(CLBLM_R_X7Y131_SLICE_X8Y131_BO5),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y131_SLICE_X8Y131_AQ),
.I3(CLBLM_R_X5Y130_SLICE_X6Y130_B5Q),
.I4(CLBLM_L_X8Y130_SLICE_X10Y130_AQ),
.I5(CLBLM_R_X5Y130_SLICE_X7Y130_BQ),
.O5(CLBLM_R_X7Y131_SLICE_X8Y131_AO5),
.O6(CLBLM_R_X7Y131_SLICE_X8Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X9Y131_DO5),
.Q(CLBLM_R_X7Y131_SLICE_X9Y131_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X9Y131_AO6),
.Q(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X9Y131_BO6),
.Q(CLBLM_R_X7Y131_SLICE_X9Y131_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X9Y131_CO6),
.Q(CLBLM_R_X7Y131_SLICE_X9Y131_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y131_SLICE_X9Y131_DO6),
.Q(CLBLM_R_X7Y131_SLICE_X9Y131_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88e4e4e4e4)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y140_SLICE_X13Y140_D5Q),
.I2(CLBLM_R_X5Y131_SLICE_X7Y131_D5Q),
.I3(CLBLL_L_X4Y137_SLICE_X5Y137_C5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_DO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33ee22dd11cc00)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_CLUT (
.I0(CLBLM_R_X7Y129_SLICE_X8Y129_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(1'b1),
.I3(CLBLM_R_X5Y130_SLICE_X7Y130_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(CLBLL_L_X4Y138_SLICE_X5Y138_D5Q),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_CO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaccffaaaac0f0)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_BLUT (
.I0(CLBLL_L_X4Y138_SLICE_X4Y138_BQ),
.I1(CLBLM_L_X10Y140_SLICE_X13Y140_D5Q),
.I2(CLBLL_L_X4Y129_SLICE_X4Y129_AQ),
.I3(CLBLM_R_X7Y131_SLICE_X9Y131_D5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y131_SLICE_X9Y131_BQ),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_BO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaff00aaaa0f0f)
  ) CLBLM_R_X7Y131_SLICE_X9Y131_ALUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_B5Q),
.I1(1'b1),
.I2(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I3(CLBLM_L_X8Y133_SLICE_X11Y133_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y133_SLICE_X6Y133_A5Q),
.O5(CLBLM_R_X7Y131_SLICE_X9Y131_AO5),
.O6(CLBLM_R_X7Y131_SLICE_X9Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X8Y132_DO5),
.Q(CLBLM_R_X7Y132_SLICE_X8Y132_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X8Y132_AO6),
.Q(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X8Y132_BO6),
.Q(CLBLM_R_X7Y132_SLICE_X8Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X8Y132_CO6),
.Q(CLBLM_R_X7Y132_SLICE_X8Y132_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X8Y132_DO6),
.Q(CLBLM_R_X7Y132_SLICE_X8Y132_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbb8888c0e2c0e2)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_DLUT (
.I0(CLBLM_R_X3Y131_SLICE_X2Y131_AQ),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y131_SLICE_X9Y131_BQ),
.I3(CLBLM_R_X7Y137_SLICE_X9Y137_D5Q),
.I4(CLBLM_R_X7Y132_SLICE_X9Y132_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_DO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hefef4545eaea4040)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y132_SLICE_X8Y132_CQ),
.I2(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.I3(1'b1),
.I4(CLBLM_L_X8Y133_SLICE_X10Y133_AQ),
.I5(CLBLM_R_X3Y132_SLICE_X2Y132_BQ),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_CO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0c5c0cac0)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_BLUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(CLBLL_L_X4Y132_SLICE_X4Y132_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y135_SLICE_X9Y135_B5Q),
.I4(CLBLM_R_X7Y133_SLICE_X8Y133_C5Q),
.I5(CLBLM_R_X7Y132_SLICE_X8Y132_BQ),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_BO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffe2f00000e2f0)
  ) CLBLM_R_X7Y132_SLICE_X8Y132_ALUT (
.I0(CLBLM_R_X7Y133_SLICE_X9Y133_B5Q),
.I1(CLBLM_R_X7Y135_SLICE_X9Y135_C5Q),
.I2(CLBLM_R_X7Y132_SLICE_X8Y132_AQ),
.I3(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_CQ),
.O5(CLBLM_R_X7Y132_SLICE_X8Y132_AO5),
.O6(CLBLM_R_X7Y132_SLICE_X8Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X9Y132_AO5),
.Q(CLBLM_R_X7Y132_SLICE_X9Y132_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X9Y132_DO5),
.Q(CLBLM_R_X7Y132_SLICE_X9Y132_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X9Y132_AO6),
.Q(CLBLM_R_X7Y132_SLICE_X9Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X9Y132_BO6),
.Q(CLBLM_R_X7Y132_SLICE_X9Y132_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X9Y132_CO6),
.Q(CLBLM_R_X7Y132_SLICE_X9Y132_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y132_SLICE_X9Y132_DO6),
.Q(CLBLM_R_X7Y132_SLICE_X9Y132_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaccf0ccf0cc)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_DLUT (
.I0(CLBLM_R_X7Y133_SLICE_X8Y133_C5Q),
.I1(CLBLL_L_X4Y134_SLICE_X4Y134_C5Q),
.I2(CLBLM_R_X7Y131_SLICE_X9Y131_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_DO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hddd888d8ddd888d8)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y133_SLICE_X9Y133_AQ),
.I2(CLBLM_R_X7Y132_SLICE_X9Y132_BQ),
.I3(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.I4(CLBLM_R_X7Y132_SLICE_X9Y132_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_CO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afafaca0acac)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_BLUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_D5Q),
.I1(CLBLM_R_X7Y132_SLICE_X9Y132_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y140_SLICE_X13Y140_D5Q),
.I4(CLBLM_R_X7Y131_SLICE_X9Y131_D5Q),
.I5(CLBLM_R_X7Y134_SLICE_X8Y134_BQ),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_BO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0afaff000ff0f)
  ) CLBLM_R_X7Y132_SLICE_X9Y132_ALUT (
.I0(CLBLM_L_X8Y133_SLICE_X11Y133_A5Q),
.I1(1'b1),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y133_SLICE_X6Y133_AQ),
.I4(CLBLM_R_X11Y142_SLICE_X14Y142_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y132_SLICE_X9Y132_AO5),
.O6(CLBLM_R_X7Y132_SLICE_X9Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X8Y133_AO5),
.Q(CLBLM_R_X7Y133_SLICE_X8Y133_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X8Y133_CO5),
.Q(CLBLM_R_X7Y133_SLICE_X8Y133_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X8Y133_DO5),
.Q(CLBLM_R_X7Y133_SLICE_X8Y133_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X8Y133_AO6),
.Q(CLBLM_R_X7Y133_SLICE_X8Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X8Y133_BO6),
.Q(CLBLM_R_X7Y133_SLICE_X8Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X8Y133_CO6),
.Q(CLBLM_R_X7Y133_SLICE_X8Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X8Y133_DO6),
.Q(CLBLM_R_X7Y133_SLICE_X8Y133_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0acacacac)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_DLUT (
.I0(CLBLM_R_X7Y132_SLICE_X9Y132_D5Q),
.I1(CLBLM_L_X12Y136_SLICE_X16Y136_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y132_SLICE_X7Y132_C5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y133_SLICE_X8Y133_DO5),
.O6(CLBLM_R_X7Y133_SLICE_X8Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaaccfff000f0)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_CLUT (
.I0(CLBLM_L_X8Y141_SLICE_X11Y141_AQ),
.I1(CLBLL_L_X4Y137_SLICE_X5Y137_C5Q),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y136_SLICE_X8Y136_DQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y133_SLICE_X8Y133_CO5),
.O6(CLBLM_R_X7Y133_SLICE_X8Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00fc000000fc)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y133_SLICE_X8Y133_BQ),
.I2(CLBLM_R_X7Y141_SLICE_X8Y141_AQ),
.I3(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y132_SLICE_X8Y132_DQ),
.O5(CLBLM_R_X7Y133_SLICE_X8Y133_BO5),
.O6(CLBLM_R_X7Y133_SLICE_X8Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0afa0afa0)
  ) CLBLM_R_X7Y133_SLICE_X8Y133_ALUT (
.I0(CLBLM_R_X7Y134_SLICE_X9Y134_DQ),
.I1(CLBLM_R_X7Y141_SLICE_X8Y141_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y133_SLICE_X4Y133_A5Q),
.I4(CLBLM_R_X5Y130_SLICE_X7Y130_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y133_SLICE_X8Y133_AO5),
.O6(CLBLM_R_X7Y133_SLICE_X8Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X9Y133_AO5),
.Q(CLBLM_R_X7Y133_SLICE_X9Y133_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X9Y133_BO5),
.Q(CLBLM_R_X7Y133_SLICE_X9Y133_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X9Y133_CO5),
.Q(CLBLM_R_X7Y133_SLICE_X9Y133_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X9Y133_DO5),
.Q(CLBLM_R_X7Y133_SLICE_X9Y133_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X9Y133_AO6),
.Q(CLBLM_R_X7Y133_SLICE_X9Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X9Y133_BO6),
.Q(CLBLM_R_X7Y133_SLICE_X9Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X9Y133_CO6),
.Q(CLBLM_R_X7Y133_SLICE_X9Y133_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y133_SLICE_X9Y133_DO6),
.Q(CLBLM_R_X7Y133_SLICE_X9Y133_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44d8d8d8d8)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X5Y133_SLICE_X7Y133_CQ),
.I2(CLBLM_L_X8Y136_SLICE_X11Y136_B5Q),
.I3(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y133_SLICE_X9Y133_DO5),
.O6(CLBLM_R_X7Y133_SLICE_X9Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00ff558888dddd)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y134_SLICE_X3Y134_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X7Y134_SLICE_X8Y134_BQ),
.I4(CLBLM_L_X10Y140_SLICE_X13Y140_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y133_SLICE_X9Y133_CO5),
.O6(CLBLM_R_X7Y133_SLICE_X9Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5cac5cafcfc0c0c)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_BLUT (
.I0(CLBLM_R_X5Y134_SLICE_X6Y134_CQ),
.I1(CLBLM_R_X3Y131_SLICE_X3Y131_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y135_SLICE_X10Y135_BQ),
.I4(CLBLL_L_X4Y131_SLICE_X5Y131_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y133_SLICE_X9Y133_BO5),
.O6(CLBLM_R_X7Y133_SLICE_X9Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0afaff101f101)
  ) CLBLM_R_X7Y133_SLICE_X9Y133_ALUT (
.I0(CLBLM_R_X5Y133_SLICE_X7Y133_DQ),
.I1(CLBLM_R_X7Y138_SLICE_X8Y138_AQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y135_SLICE_X10Y135_BQ),
.I4(CLBLM_L_X10Y140_SLICE_X13Y140_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y133_SLICE_X9Y133_AO5),
.O6(CLBLM_R_X7Y133_SLICE_X9Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X8Y134_AO5),
.Q(CLBLM_R_X7Y134_SLICE_X8Y134_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X8Y134_BO5),
.Q(CLBLM_R_X7Y134_SLICE_X8Y134_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X8Y134_CO5),
.Q(CLBLM_R_X7Y134_SLICE_X8Y134_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X8Y134_AO6),
.Q(CLBLM_R_X7Y134_SLICE_X8Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X8Y134_BO6),
.Q(CLBLM_R_X7Y134_SLICE_X8Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X8Y134_CO6),
.Q(CLBLM_R_X7Y134_SLICE_X8Y134_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3fff3fff0fff0fff)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y134_SLICE_X9Y134_BQ),
.I2(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I3(CLBLM_R_X7Y138_SLICE_X8Y138_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y134_SLICE_X8Y134_DO5),
.O6(CLBLM_R_X7Y134_SLICE_X8Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaaaaaa00cc)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_CLUT (
.I0(CLBLM_R_X7Y133_SLICE_X9Y133_D5Q),
.I1(CLBLL_L_X2Y138_SLICE_X1Y138_BO6),
.I2(CLBLL_L_X4Y135_SLICE_X4Y135_DQ),
.I3(CLBLM_R_X7Y140_SLICE_X9Y140_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y134_SLICE_X8Y134_CO5),
.O6(CLBLM_R_X7Y134_SLICE_X8Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfc0c0f505fa0a)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_BLUT (
.I0(CLBLM_R_X7Y136_SLICE_X8Y136_B5Q),
.I1(CLBLM_R_X5Y134_SLICE_X7Y134_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y134_SLICE_X9Y134_BQ),
.I4(CLBLM_R_X5Y134_SLICE_X6Y134_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y134_SLICE_X8Y134_BO5),
.O6(CLBLM_R_X7Y134_SLICE_X8Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f000ffcccc00ff)
  ) CLBLM_R_X7Y134_SLICE_X8Y134_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y135_SLICE_X4Y135_BQ),
.I2(CLBLM_L_X8Y136_SLICE_X10Y136_BQ),
.I3(CLBLM_L_X12Y136_SLICE_X16Y136_AQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y134_SLICE_X8Y134_AO5),
.O6(CLBLM_R_X7Y134_SLICE_X8Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X9Y134_AO6),
.Q(CLBLM_R_X7Y134_SLICE_X9Y134_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X9Y134_BO6),
.Q(CLBLM_R_X7Y134_SLICE_X9Y134_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X9Y134_CO6),
.Q(CLBLM_R_X7Y134_SLICE_X9Y134_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y134_SLICE_X9Y134_DO6),
.Q(CLBLM_R_X7Y134_SLICE_X9Y134_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaafa00550050)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(CLBLM_R_X7Y134_SLICE_X9Y134_DQ),
.I3(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.I4(CLBLL_L_X4Y134_SLICE_X4Y134_AQ),
.I5(CLBLM_R_X7Y134_SLICE_X9Y134_AQ),
.O5(CLBLM_R_X7Y134_SLICE_X9Y134_DO5),
.O6(CLBLM_R_X7Y134_SLICE_X9Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaca0acafafa0a0)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_CLUT (
.I0(CLBLM_R_X7Y138_SLICE_X8Y138_AQ),
.I1(CLBLM_R_X7Y134_SLICE_X9Y134_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_CQ),
.I4(CLBLM_R_X7Y138_SLICE_X9Y138_A5Q),
.I5(CLBLL_L_X4Y136_SLICE_X4Y136_D5Q),
.O5(CLBLM_R_X7Y134_SLICE_X9Y134_CO5),
.O6(CLBLM_R_X7Y134_SLICE_X9Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafc0a0cfaf30a03)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_BLUT (
.I0(CLBLM_L_X8Y134_SLICE_X11Y134_B5Q),
.I1(CLBLM_R_X7Y134_SLICE_X8Y134_DO5),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y133_SLICE_X6Y133_A5Q),
.I4(CLBLM_R_X7Y140_SLICE_X9Y140_D5Q),
.I5(CLBLM_R_X7Y134_SLICE_X9Y134_BQ),
.O5(CLBLM_R_X7Y134_SLICE_X9Y134_BO5),
.O6(CLBLM_R_X7Y134_SLICE_X9Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa3a3afa0a3a0)
  ) CLBLM_R_X7Y134_SLICE_X9Y134_ALUT (
.I0(CLBLM_R_X7Y133_SLICE_X8Y133_AQ),
.I1(CLBLL_L_X4Y135_SLICE_X4Y135_D5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y134_SLICE_X9Y134_AQ),
.I4(CLBLM_R_X5Y133_SLICE_X7Y133_AQ),
.I5(CLBLM_R_X7Y138_SLICE_X9Y138_CQ),
.O5(CLBLM_R_X7Y134_SLICE_X9Y134_AO5),
.O6(CLBLM_R_X7Y134_SLICE_X9Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X3Y135_SLICE_X3Y135_BQ),
.Q(CLBLM_R_X7Y135_SLICE_X8Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X7Y134_SLICE_X8Y134_B5Q),
.Q(CLBLM_R_X7Y135_SLICE_X8Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf444fffff444f444)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_DLUT (
.I0(CLBLM_L_X12Y134_SLICE_X17Y134_AO6),
.I1(CLBLM_R_X7Y132_SLICE_X8Y132_CQ),
.I2(CLBLM_R_X3Y135_SLICE_X2Y135_BQ),
.I3(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.I4(CLBLM_L_X10Y137_SLICE_X13Y137_BO6),
.I5(CLBLM_R_X5Y135_SLICE_X7Y135_BQ),
.O5(CLBLM_R_X7Y135_SLICE_X8Y135_DO5),
.O6(CLBLM_R_X7Y135_SLICE_X8Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f33bfbb0f00afaa)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_CLUT (
.I0(CLBLM_R_X3Y135_SLICE_X3Y135_AQ),
.I1(CLBLM_R_X11Y133_SLICE_X14Y133_CO5),
.I2(CLBLM_L_X10Y137_SLICE_X13Y137_BO6),
.I3(CLBLL_L_X4Y138_SLICE_X5Y138_A5Q),
.I4(CLBLM_L_X12Y135_SLICE_X16Y135_AO6),
.I5(CLBLM_R_X7Y135_SLICE_X9Y135_BQ),
.O5(CLBLM_R_X7Y135_SLICE_X8Y135_CO5),
.O6(CLBLM_R_X7Y135_SLICE_X8Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f3f5f0f77335500)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_BLUT (
.I0(CLBLM_L_X10Y137_SLICE_X13Y137_BO6),
.I1(CLBLM_L_X12Y135_SLICE_X16Y135_AO6),
.I2(CLBLM_R_X11Y133_SLICE_X14Y133_CO5),
.I3(CLBLL_L_X4Y132_SLICE_X5Y132_D5Q),
.I4(CLBLL_L_X4Y132_SLICE_X5Y132_AQ),
.I5(CLBLL_L_X4Y135_SLICE_X4Y135_BQ),
.O5(CLBLM_R_X7Y135_SLICE_X8Y135_BO5),
.O6(CLBLM_R_X7Y135_SLICE_X8Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X7Y135_SLICE_X8Y135_ALUT (
.I0(CLBLM_R_X7Y136_SLICE_X8Y136_DQ),
.I1(CLBLL_L_X4Y133_SLICE_X5Y133_DQ),
.I2(CLBLM_R_X7Y135_SLICE_X9Y135_A5Q),
.I3(CLBLL_L_X4Y135_SLICE_X4Y135_C5Q),
.I4(CLBLM_L_X8Y135_SLICE_X10Y135_DQ),
.I5(CLBLM_R_X7Y134_SLICE_X8Y134_B5Q),
.O5(CLBLM_R_X7Y135_SLICE_X8Y135_AO5),
.O6(CLBLM_R_X7Y135_SLICE_X8Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y135_SLICE_X9Y135_AO5),
.Q(CLBLM_R_X7Y135_SLICE_X9Y135_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y135_SLICE_X5Y135_DO5),
.Q(CLBLM_R_X7Y135_SLICE_X9Y135_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y135_SLICE_X9Y135_CO5),
.Q(CLBLM_R_X7Y135_SLICE_X9Y135_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y135_SLICE_X9Y135_DO5),
.Q(CLBLM_R_X7Y135_SLICE_X9Y135_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y135_SLICE_X9Y135_AO6),
.Q(CLBLM_R_X7Y135_SLICE_X9Y135_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y135_SLICE_X9Y135_BO6),
.Q(CLBLM_R_X7Y135_SLICE_X9Y135_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y135_SLICE_X9Y135_CO6),
.Q(CLBLM_R_X7Y135_SLICE_X9Y135_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y135_SLICE_X9Y135_DO6),
.Q(CLBLM_R_X7Y135_SLICE_X9Y135_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbee1144f5a0f5a0)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X10Y135_SLICE_X13Y135_AQ),
.I2(CLBLM_R_X5Y142_SLICE_X6Y142_B5Q),
.I3(CLBLL_L_X4Y137_SLICE_X5Y137_C5Q),
.I4(CLBLM_L_X8Y139_SLICE_X11Y139_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y135_SLICE_X9Y135_DO5),
.O6(CLBLM_R_X7Y135_SLICE_X9Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfc0cacacacac)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_CLUT (
.I0(CLBLM_R_X7Y130_SLICE_X9Y130_AQ),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y140_SLICE_X8Y140_C5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y135_SLICE_X9Y135_CO5),
.O6(CLBLM_R_X7Y135_SLICE_X9Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f00000ffcc)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y135_SLICE_X9Y135_BQ),
.I2(CLBLM_R_X3Y134_SLICE_X2Y134_AQ),
.I3(CLBLM_R_X7Y130_SLICE_X9Y130_AQ),
.I4(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X7Y135_SLICE_X9Y135_BO5),
.O6(CLBLM_R_X7Y135_SLICE_X9Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0a0af606f606)
  ) CLBLM_R_X7Y135_SLICE_X9Y135_ALUT (
.I0(CLBLL_L_X4Y138_SLICE_X5Y138_DQ),
.I1(CLBLM_L_X10Y140_SLICE_X12Y140_D5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y134_SLICE_X6Y134_A5Q),
.I4(CLBLM_R_X3Y135_SLICE_X2Y135_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y135_SLICE_X9Y135_AO5),
.O6(CLBLM_R_X7Y135_SLICE_X9Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X8Y136_AO5),
.Q(CLBLM_R_X7Y136_SLICE_X8Y136_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X8Y136_BO5),
.Q(CLBLM_R_X7Y136_SLICE_X8Y136_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X8Y136_CO5),
.Q(CLBLM_R_X7Y136_SLICE_X8Y136_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X8Y136_DO5),
.Q(CLBLM_R_X7Y136_SLICE_X8Y136_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X8Y136_AO6),
.Q(CLBLM_R_X7Y136_SLICE_X8Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X8Y136_BO6),
.Q(CLBLM_R_X7Y136_SLICE_X8Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X8Y136_CO6),
.Q(CLBLM_R_X7Y136_SLICE_X8Y136_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X8Y136_DO6),
.Q(CLBLM_R_X7Y136_SLICE_X8Y136_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5cac5cafcfc0c0c)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_DLUT (
.I0(CLBLM_R_X3Y135_SLICE_X3Y135_CQ),
.I1(CLBLM_L_X10Y141_SLICE_X12Y141_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y132_SLICE_X9Y132_A5Q),
.I4(CLBLM_R_X3Y135_SLICE_X2Y135_DQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y136_SLICE_X8Y136_DO5),
.O6(CLBLM_R_X7Y136_SLICE_X8Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacacaccfc0cfc0)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_CLUT (
.I0(CLBLM_R_X5Y140_SLICE_X7Y140_A5Q),
.I1(CLBLM_R_X7Y131_SLICE_X8Y131_A5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y131_SLICE_X12Y131_D5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y136_SLICE_X8Y136_CO5),
.O6(CLBLM_R_X7Y136_SLICE_X8Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a0f5a0dd88dd88)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I2(CLBLM_R_X3Y138_SLICE_X2Y138_AQ),
.I3(CLBLM_L_X12Y136_SLICE_X16Y136_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y136_SLICE_X8Y136_BO5),
.O6(CLBLM_R_X7Y136_SLICE_X8Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00f0f0f0aaaa)
  ) CLBLM_R_X7Y136_SLICE_X8Y136_ALUT (
.I0(CLBLM_R_X7Y130_SLICE_X9Y130_BQ),
.I1(CLBLM_R_X7Y135_SLICE_X9Y135_A5Q),
.I2(CLBLM_R_X7Y136_SLICE_X8Y136_AQ),
.I3(CLBLM_R_X7Y133_SLICE_X8Y133_DQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y136_SLICE_X8Y136_AO5),
.O6(CLBLM_R_X7Y136_SLICE_X8Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X9Y136_AO5),
.Q(CLBLM_R_X7Y136_SLICE_X9Y136_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X9Y136_DO5),
.Q(CLBLM_R_X7Y136_SLICE_X9Y136_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X9Y136_AO6),
.Q(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X9Y136_BO6),
.Q(CLBLM_R_X7Y136_SLICE_X9Y136_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X9Y136_CO6),
.Q(CLBLM_R_X7Y136_SLICE_X9Y136_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y136_SLICE_X9Y136_DO6),
.Q(CLBLM_R_X7Y136_SLICE_X9Y136_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf0aaf0aaf0)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_DLUT (
.I0(CLBLM_R_X7Y138_SLICE_X9Y138_AQ),
.I1(CLBLM_R_X5Y131_SLICE_X7Y131_AQ),
.I2(CLBLM_R_X5Y134_SLICE_X6Y134_DQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y136_SLICE_X9Y136_DO5),
.O6(CLBLM_R_X7Y136_SLICE_X9Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff002222ff008888)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_CLUT (
.I0(CLBLM_R_X5Y141_SLICE_X6Y141_AQ),
.I1(CLBLM_R_X7Y136_SLICE_X9Y136_CQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y136_SLICE_X7Y136_CQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X8Y136_SLICE_X10Y136_AO6),
.O5(CLBLM_R_X7Y136_SLICE_X9Y136_CO5),
.O6(CLBLM_R_X7Y136_SLICE_X9Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaee5044faee5044)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y136_SLICE_X9Y136_BQ),
.I2(CLBLM_R_X7Y134_SLICE_X9Y134_AQ),
.I3(CLBLM_R_X11Y131_SLICE_X14Y131_BO6),
.I4(CLBLM_R_X7Y136_SLICE_X9Y136_DQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y136_SLICE_X9Y136_BO5),
.O6(CLBLM_R_X7Y136_SLICE_X9Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0f5f5aa00ff55)
  ) CLBLM_R_X7Y136_SLICE_X9Y136_ALUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(1'b1),
.I2(CLBLM_L_X8Y136_SLICE_X10Y136_AQ),
.I3(CLBLM_R_X7Y136_SLICE_X9Y136_D5Q),
.I4(CLBLM_R_X11Y142_SLICE_X14Y142_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y136_SLICE_X9Y136_AO5),
.O6(CLBLM_R_X7Y136_SLICE_X9Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y137_SLICE_X8Y137_BO5),
.Q(CLBLM_R_X7Y137_SLICE_X8Y137_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y137_SLICE_X8Y137_CO5),
.Q(CLBLM_R_X7Y137_SLICE_X8Y137_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y137_SLICE_X8Y137_DO5),
.Q(CLBLM_R_X7Y137_SLICE_X8Y137_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y137_SLICE_X8Y137_AO6),
.Q(CLBLM_R_X7Y137_SLICE_X8Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y137_SLICE_X8Y137_BO6),
.Q(CLBLM_R_X7Y137_SLICE_X8Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y137_SLICE_X8Y137_CO6),
.Q(CLBLM_R_X7Y137_SLICE_X8Y137_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y137_SLICE_X8Y137_DO6),
.Q(CLBLM_R_X7Y137_SLICE_X8Y137_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc00ccf0fff000)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y136_SLICE_X7Y136_CQ),
.I2(CLBLM_R_X7Y138_SLICE_X8Y138_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y137_SLICE_X9Y137_DQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X8Y137_DO5),
.O6(CLBLM_R_X7Y137_SLICE_X8Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0ff00cccc)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y137_SLICE_X5Y137_AQ),
.I2(CLBLM_L_X12Y136_SLICE_X16Y136_A5Q),
.I3(CLBLM_L_X8Y135_SLICE_X10Y135_B5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X8Y137_CO5),
.O6(CLBLM_R_X7Y137_SLICE_X8Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0fcc0faaf0aaf0)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_BLUT (
.I0(CLBLM_R_X7Y140_SLICE_X8Y140_B5Q),
.I1(CLBLM_L_X8Y137_SLICE_X10Y137_CQ),
.I2(CLBLL_L_X4Y131_SLICE_X5Y131_B5Q),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X8Y137_BO5),
.O6(CLBLM_R_X7Y137_SLICE_X8Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaf0aa33aa30)
  ) CLBLM_R_X7Y137_SLICE_X8Y137_ALUT (
.I0(CLBLM_R_X7Y133_SLICE_X8Y133_DQ),
.I1(CLBLM_R_X7Y131_SLICE_X9Y131_D5Q),
.I2(CLBLM_R_X7Y137_SLICE_X8Y137_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y138_SLICE_X8Y138_B5Q),
.I5(CLBLM_L_X10Y140_SLICE_X13Y140_D5Q),
.O5(CLBLM_R_X7Y137_SLICE_X8Y137_AO5),
.O6(CLBLM_R_X7Y137_SLICE_X8Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y137_SLICE_X9Y137_DO5),
.Q(CLBLM_R_X7Y137_SLICE_X9Y137_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y137_SLICE_X9Y137_AO6),
.Q(CLBLM_R_X7Y137_SLICE_X9Y137_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y137_SLICE_X9Y137_BO6),
.Q(CLBLM_R_X7Y137_SLICE_X9Y137_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y137_SLICE_X9Y137_CO6),
.Q(CLBLM_R_X7Y137_SLICE_X9Y137_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y137_SLICE_X9Y137_DO6),
.Q(CLBLM_R_X7Y137_SLICE_X9Y137_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00ccaaf0ccf0cc)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_DLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_R_X7Y131_SLICE_X9Y131_CQ),
.I2(CLBLM_L_X8Y139_SLICE_X11Y139_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLL_L_X4Y138_SLICE_X4Y138_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X9Y137_DO5),
.O6(CLBLM_R_X7Y137_SLICE_X9Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff5fcf40f050c04)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_CLUT (
.I0(CLBLL_L_X4Y136_SLICE_X4Y136_D5Q),
.I1(CLBLM_R_X7Y137_SLICE_X9Y137_CQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_CQ),
.I4(CLBLM_R_X7Y135_SLICE_X9Y135_AQ),
.I5(CLBLM_R_X7Y143_SLICE_X8Y143_A5Q),
.O5(CLBLM_R_X7Y137_SLICE_X9Y137_CO5),
.O6(CLBLM_R_X7Y137_SLICE_X9Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfa0afc0cfa0a)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_BLUT (
.I0(CLBLM_R_X7Y137_SLICE_X9Y137_CQ),
.I1(CLBLM_R_X7Y137_SLICE_X9Y137_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y137_SLICE_X9Y137_D5Q),
.I4(CLBLM_L_X12Y132_SLICE_X16Y132_AO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y137_SLICE_X9Y137_BO5),
.O6(CLBLM_R_X7Y137_SLICE_X9Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaccffc0f0)
  ) CLBLM_R_X7Y137_SLICE_X9Y137_ALUT (
.I0(CLBLM_R_X7Y137_SLICE_X9Y137_CQ),
.I1(CLBLM_R_X5Y133_SLICE_X7Y133_AQ),
.I2(CLBLM_R_X7Y137_SLICE_X9Y137_AQ),
.I3(CLBLL_L_X4Y135_SLICE_X4Y135_D5Q),
.I4(CLBLM_R_X5Y135_SLICE_X6Y135_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X7Y137_SLICE_X9Y137_AO5),
.O6(CLBLM_R_X7Y137_SLICE_X9Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y138_SLICE_X8Y138_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y138_SLICE_X8Y138_BO5),
.Q(CLBLM_R_X7Y138_SLICE_X8Y138_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y138_SLICE_X8Y138_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y138_SLICE_X8Y138_DO5),
.Q(CLBLM_R_X7Y138_SLICE_X8Y138_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y138_SLICE_X8Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y138_SLICE_X8Y138_AO6),
.Q(CLBLM_R_X7Y138_SLICE_X8Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y138_SLICE_X8Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y138_SLICE_X8Y138_BO6),
.Q(CLBLM_R_X7Y138_SLICE_X8Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y138_SLICE_X8Y138_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y138_SLICE_X8Y138_CO6),
.Q(CLBLM_R_X7Y138_SLICE_X8Y138_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y138_SLICE_X8Y138_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y138_SLICE_X8Y138_DO6),
.Q(CLBLM_R_X7Y138_SLICE_X8Y138_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3a3acacfc0cfc0c)
  ) CLBLM_R_X7Y138_SLICE_X8Y138_DLUT (
.I0(CLBLM_R_X5Y136_SLICE_X7Y136_AQ),
.I1(CLBLM_R_X7Y130_SLICE_X9Y130_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y139_SLICE_X6Y139_AQ),
.I4(CLBLL_L_X4Y138_SLICE_X5Y138_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y138_SLICE_X8Y138_DO5),
.O6(CLBLM_R_X7Y138_SLICE_X8Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff0660000f066)
  ) CLBLM_R_X7Y138_SLICE_X8Y138_CLUT (
.I0(CLBLM_R_X7Y131_SLICE_X9Y131_AQ),
.I1(CLBLM_R_X7Y138_SLICE_X8Y138_CQ),
.I2(CLBLM_R_X7Y140_SLICE_X8Y140_CQ),
.I3(CLBLM_R_X5Y133_SLICE_X6Y133_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X10Y138_SLICE_X13Y138_BQ),
.O5(CLBLM_R_X7Y138_SLICE_X8Y138_CO5),
.O6(CLBLM_R_X7Y138_SLICE_X8Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf505fa0acacacaca)
  ) CLBLM_R_X7Y138_SLICE_X8Y138_BLUT (
.I0(CLBLM_R_X5Y140_SLICE_X6Y140_CQ),
.I1(CLBLM_R_X7Y135_SLICE_X8Y135_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X5Y139_SLICE_X7Y139_B5Q),
.I4(CLBLM_R_X3Y135_SLICE_X3Y135_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y138_SLICE_X8Y138_BO5),
.O6(CLBLM_R_X7Y138_SLICE_X8Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcfffc0f0c0f0c)
  ) CLBLM_R_X7Y138_SLICE_X8Y138_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y138_SLICE_X7Y138_BO6),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X7Y139_SLICE_X8Y139_BO6),
.I4(1'b1),
.I5(CLBLM_L_X8Y131_SLICE_X11Y131_CQ),
.O5(CLBLM_R_X7Y138_SLICE_X8Y138_AO5),
.O6(CLBLM_R_X7Y138_SLICE_X8Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y138_SLICE_X9Y138_AO5),
.Q(CLBLM_R_X7Y138_SLICE_X9Y138_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y138_SLICE_X9Y138_BO5),
.Q(CLBLM_R_X7Y138_SLICE_X9Y138_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y138_SLICE_X9Y138_CO5),
.Q(CLBLM_R_X7Y138_SLICE_X9Y138_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y138_SLICE_X9Y138_AO6),
.Q(CLBLM_R_X7Y138_SLICE_X9Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y138_SLICE_X9Y138_BO6),
.Q(CLBLM_R_X7Y138_SLICE_X9Y138_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y138_SLICE_X9Y138_CO6),
.Q(CLBLM_R_X7Y138_SLICE_X9Y138_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000001000)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_DLUT (
.I0(CLBLM_R_X5Y135_SLICE_X6Y135_CO5),
.I1(CLBLM_R_X11Y138_SLICE_X15Y138_CO6),
.I2(CLBLL_L_X4Y138_SLICE_X4Y138_BO5),
.I3(CLBLM_L_X12Y139_SLICE_X17Y139_AO6),
.I4(CLBLM_R_X5Y130_SLICE_X7Y130_DQ),
.I5(CLBLM_L_X8Y143_SLICE_X10Y143_BO6),
.O5(CLBLM_R_X7Y138_SLICE_X9Y138_DO5),
.O6(CLBLM_R_X7Y138_SLICE_X9Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaaaff00aaaa)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_CLUT (
.I0(CLBLM_R_X5Y134_SLICE_X6Y134_CQ),
.I1(CLBLM_R_X3Y138_SLICE_X2Y138_CQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y138_SLICE_X9Y138_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y138_SLICE_X9Y138_CO5),
.O6(CLBLM_R_X7Y138_SLICE_X9Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00aaaaccccffa5)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_BLUT (
.I0(CLBLM_R_X7Y138_SLICE_X9Y138_B5Q),
.I1(CLBLM_L_X10Y141_SLICE_X12Y141_AQ),
.I2(CLBLM_R_X5Y138_SLICE_X7Y138_CO6),
.I3(CLBLM_R_X5Y130_SLICE_X7Y130_DQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y138_SLICE_X9Y138_BO5),
.O6(CLBLM_R_X7Y138_SLICE_X9Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf055f0aaccffcc00)
  ) CLBLM_R_X7Y138_SLICE_X9Y138_ALUT (
.I0(CLBLM_R_X3Y140_SLICE_X3Y140_C5Q),
.I1(CLBLM_R_X3Y133_SLICE_X3Y133_B5Q),
.I2(CLBLM_L_X10Y139_SLICE_X13Y139_CQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y138_SLICE_X9Y138_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y138_SLICE_X9Y138_AO5),
.O6(CLBLM_R_X7Y138_SLICE_X9Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X8Y137_SLICE_X10Y137_B5Q),
.Q(CLBLM_R_X7Y139_SLICE_X8Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hacaaacaaacaaacaa)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_DLUT (
.I0(CLBLM_R_X7Y141_SLICE_X8Y141_AQ),
.I1(CLBLM_R_X5Y139_SLICE_X6Y139_CQ),
.I2(CLBLM_R_X7Y135_SLICE_X9Y135_C5Q),
.I3(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y139_SLICE_X8Y139_DO5),
.O6(CLBLM_R_X7Y139_SLICE_X8Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffafffa)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_CLUT (
.I0(CLBLM_R_X7Y138_SLICE_X9Y138_AQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y139_SLICE_X4Y139_A5Q),
.I3(CLBLM_L_X8Y137_SLICE_X10Y137_B5Q),
.I4(1'b1),
.I5(CLBLM_R_X7Y138_SLICE_X8Y138_BQ),
.O5(CLBLM_R_X7Y139_SLICE_X8Y139_CO5),
.O6(CLBLM_R_X7Y139_SLICE_X8Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffefffefffe)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_BLUT (
.I0(CLBLM_R_X5Y134_SLICE_X6Y134_DQ),
.I1(CLBLM_R_X5Y140_SLICE_X6Y140_CQ),
.I2(CLBLM_R_X3Y135_SLICE_X3Y135_DQ),
.I3(CLBLM_R_X5Y132_SLICE_X6Y132_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y139_SLICE_X8Y139_BO5),
.O6(CLBLM_R_X7Y139_SLICE_X8Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00010000fffcfffc)
  ) CLBLM_R_X7Y139_SLICE_X8Y139_ALUT (
.I0(CLBLL_L_X4Y138_SLICE_X4Y138_CO6),
.I1(CLBLM_R_X7Y140_SLICE_X9Y140_DQ),
.I2(CLBLM_R_X5Y138_SLICE_X6Y138_BQ),
.I3(CLBLM_R_X7Y135_SLICE_X9Y135_DQ),
.I4(CLBLM_R_X7Y135_SLICE_X8Y135_AO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y139_SLICE_X8Y139_AO5),
.O6(CLBLM_R_X7Y139_SLICE_X8Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y139_SLICE_X9Y139_AO6),
.Q(CLBLM_R_X7Y139_SLICE_X9Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y139_SLICE_X9Y139_BO6),
.Q(CLBLM_R_X7Y139_SLICE_X9Y139_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000400000004)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_DLUT (
.I0(CLBLM_R_X5Y140_SLICE_X6Y140_CQ),
.I1(CLBLM_R_X7Y138_SLICE_X9Y138_DO6),
.I2(CLBLL_L_X4Y138_SLICE_X4Y138_CO6),
.I3(CLBLM_R_X5Y141_SLICE_X7Y141_CO6),
.I4(CLBLM_L_X10Y141_SLICE_X13Y141_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y139_SLICE_X9Y139_DO5),
.O6(CLBLM_R_X7Y139_SLICE_X9Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffa)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_CLUT (
.I0(CLBLM_R_X5Y138_SLICE_X6Y138_BQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y134_SLICE_X8Y134_DO6),
.I3(CLBLM_R_X7Y140_SLICE_X9Y140_DQ),
.I4(CLBLM_R_X3Y133_SLICE_X3Y133_DO6),
.I5(CLBLM_R_X7Y135_SLICE_X9Y135_DQ),
.O5(CLBLM_R_X7Y139_SLICE_X9Y139_CO5),
.O6(CLBLM_R_X7Y139_SLICE_X9Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0f5f5e4e4)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y139_SLICE_X9Y139_BQ),
.I2(CLBLM_R_X7Y137_SLICE_X9Y137_AQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y140_SLICE_X10Y140_AQ),
.I5(CLBLM_L_X12Y132_SLICE_X16Y132_AO6),
.O5(CLBLM_R_X7Y139_SLICE_X9Y139_BO5),
.O6(CLBLM_R_X7Y139_SLICE_X9Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcccfc33300030)
  ) CLBLM_R_X7Y139_SLICE_X9Y139_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y139_SLICE_X9Y139_AQ),
.I3(CLBLM_R_X11Y131_SLICE_X14Y131_BO6),
.I4(CLBLM_R_X7Y137_SLICE_X9Y137_AQ),
.I5(CLBLM_R_X5Y139_SLICE_X7Y139_A5Q),
.O5(CLBLM_R_X7Y139_SLICE_X9Y139_AO5),
.O6(CLBLM_R_X7Y139_SLICE_X9Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y140_SLICE_X8Y140_BO5),
.Q(CLBLM_R_X7Y140_SLICE_X8Y140_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y140_SLICE_X8Y140_CO5),
.Q(CLBLM_R_X7Y140_SLICE_X8Y140_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y140_SLICE_X8Y140_DO5),
.Q(CLBLM_R_X7Y140_SLICE_X8Y140_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y140_SLICE_X8Y140_AO6),
.Q(CLBLM_R_X7Y140_SLICE_X8Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y140_SLICE_X8Y140_BO6),
.Q(CLBLM_R_X7Y140_SLICE_X8Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y140_SLICE_X8Y140_CO6),
.Q(CLBLM_R_X7Y140_SLICE_X8Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y140_SLICE_X8Y140_DO6),
.Q(CLBLM_R_X7Y140_SLICE_X8Y140_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafa0afa0fff00f00)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_DLUT (
.I0(CLBLL_L_X4Y140_SLICE_X5Y140_BQ),
.I1(1'b1),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_R_X11Y141_SLICE_X14Y141_AQ),
.I4(CLBLL_L_X4Y136_SLICE_X5Y136_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y140_SLICE_X8Y140_DO5),
.O6(CLBLM_R_X7Y140_SLICE_X8Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccaaffcc00cc)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_CLUT (
.I0(CLBLM_R_X7Y133_SLICE_X8Y133_D5Q),
.I1(CLBLM_R_X3Y139_SLICE_X2Y139_CQ),
.I2(1'b1),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_L_X10Y142_SLICE_X12Y142_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y140_SLICE_X8Y140_CO5),
.O6(CLBLM_R_X7Y140_SLICE_X8Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d8affa0550)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_BLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_L_X8Y140_SLICE_X10Y140_D5Q),
.I2(CLBLM_R_X3Y135_SLICE_X3Y135_BQ),
.I3(CLBLM_R_X5Y135_SLICE_X7Y135_BQ),
.I4(CLBLM_L_X8Y143_SLICE_X11Y143_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y140_SLICE_X8Y140_BO5),
.O6(CLBLM_R_X7Y140_SLICE_X8Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbbb00000bbb0)
  ) CLBLM_R_X7Y140_SLICE_X8Y140_ALUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_CQ),
.I1(CLBLL_L_X4Y136_SLICE_X4Y136_D5Q),
.I2(CLBLM_R_X7Y140_SLICE_X8Y140_AQ),
.I3(CLBLM_R_X5Y135_SLICE_X7Y135_D5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y141_SLICE_X9Y141_A5Q),
.O5(CLBLM_R_X7Y140_SLICE_X8Y140_AO5),
.O6(CLBLM_R_X7Y140_SLICE_X8Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_D5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y140_SLICE_X9Y140_DO5),
.Q(CLBLM_R_X7Y140_SLICE_X9Y140_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y140_SLICE_X9Y140_AO6),
.Q(CLBLM_R_X7Y140_SLICE_X9Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y140_SLICE_X9Y140_BO6),
.Q(CLBLM_R_X7Y140_SLICE_X9Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y140_SLICE_X9Y140_CO6),
.Q(CLBLM_R_X7Y140_SLICE_X9Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y140_SLICE_X9Y140_DO6),
.Q(CLBLM_R_X7Y140_SLICE_X9Y140_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff006666f0f0ff00)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_DLUT (
.I0(CLBLM_R_X7Y133_SLICE_X9Y133_AQ),
.I1(CLBLM_R_X5Y134_SLICE_X6Y134_DQ),
.I2(CLBLM_L_X10Y141_SLICE_X13Y141_CQ),
.I3(CLBLM_R_X7Y136_SLICE_X8Y136_D5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y140_SLICE_X9Y140_DO5),
.O6(CLBLM_R_X7Y140_SLICE_X9Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0f5e4e4a0e4)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_CLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X7Y140_SLICE_X9Y140_CQ),
.I2(CLBLM_L_X10Y131_SLICE_X12Y131_D5Q),
.I3(CLBLL_L_X4Y135_SLICE_X5Y135_CQ),
.I4(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.I5(CLBLM_R_X7Y138_SLICE_X8Y138_D5Q),
.O5(CLBLM_R_X7Y140_SLICE_X9Y140_CO5),
.O6(CLBLM_R_X7Y140_SLICE_X9Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f02222f0f00000)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_R_X7Y140_SLICE_X9Y140_BQ),
.I2(CLBLM_R_X7Y140_SLICE_X9Y140_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y134_SLICE_X8Y134_C5Q),
.O5(CLBLM_R_X7Y140_SLICE_X9Y140_BO5),
.O6(CLBLM_R_X7Y140_SLICE_X9Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccf5a0f0f0)
  ) CLBLM_R_X7Y140_SLICE_X9Y140_ALUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_C5Q),
.I1(CLBLM_R_X7Y138_SLICE_X8Y138_D5Q),
.I2(CLBLM_R_X7Y140_SLICE_X9Y140_AQ),
.I3(CLBLM_L_X8Y138_SLICE_X11Y138_C5Q),
.I4(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X7Y140_SLICE_X9Y140_AO5),
.O6(CLBLM_R_X7Y140_SLICE_X9Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X9Y142_DO6),
.Q(CLBLM_R_X7Y141_SLICE_X8Y141_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y141_SLICE_X8Y141_AO6),
.Q(CLBLM_R_X7Y141_SLICE_X8Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff733333ff333333)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_DLUT (
.I0(CLBLM_L_X8Y140_SLICE_X10Y140_DQ),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLM_R_X7Y141_SLICE_X8Y141_BO5),
.I5(CLBLL_L_X4Y139_SLICE_X4Y139_AQ),
.O5(CLBLM_R_X7Y141_SLICE_X8Y141_DO5),
.O6(CLBLM_R_X7Y141_SLICE_X8Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3737373733373737)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_CLUT (
.I0(CLBLL_L_X2Y138_SLICE_X1Y138_BO6),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(CLBLL_L_X4Y140_SLICE_X5Y140_BQ),
.I3(CLBLM_R_X7Y134_SLICE_X8Y134_C5Q),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_R_X7Y140_SLICE_X9Y140_BQ),
.O5(CLBLM_R_X7Y141_SLICE_X8Y141_CO5),
.O6(CLBLM_R_X7Y141_SLICE_X8Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0a0000003133)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLL_L_X4Y140_SLICE_X5Y140_BQ),
.I2(CLBLM_R_X7Y140_SLICE_X9Y140_BQ),
.I3(CLBLM_R_X7Y134_SLICE_X8Y134_C5Q),
.I4(CLBLL_L_X2Y138_SLICE_X1Y138_BO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y141_SLICE_X8Y141_BO5),
.O6(CLBLM_R_X7Y141_SLICE_X8Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd31fc30ec20fc30)
  ) CLBLM_R_X7Y141_SLICE_X8Y141_ALUT (
.I0(CLBLM_R_X7Y135_SLICE_X9Y135_C5Q),
.I1(LIOB33_X0Y61_IOB_X0Y62_I),
.I2(CLBLM_R_X7Y141_SLICE_X8Y141_AQ),
.I3(CLBLM_R_X5Y142_SLICE_X6Y142_CQ),
.I4(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.I5(CLBLM_R_X5Y139_SLICE_X6Y139_CQ),
.O5(CLBLM_R_X7Y141_SLICE_X8Y141_AO5),
.O6(CLBLM_R_X7Y141_SLICE_X8Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y141_SLICE_X9Y141_AO5),
.Q(CLBLM_R_X7Y141_SLICE_X9Y141_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y141_SLICE_X9Y141_AO6),
.Q(CLBLM_R_X7Y141_SLICE_X9Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y141_SLICE_X9Y141_DO5),
.O6(CLBLM_R_X7Y141_SLICE_X9Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y141_SLICE_X9Y141_CO5),
.O6(CLBLM_R_X7Y141_SLICE_X9Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf070f070f070f070)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_R_X7Y134_SLICE_X8Y134_C5Q),
.I2(CLBLM_R_X3Y135_SLICE_X2Y135_AQ),
.I3(CLBLM_R_X7Y140_SLICE_X9Y140_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y141_SLICE_X9Y141_BO5),
.O6(CLBLM_R_X7Y141_SLICE_X9Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00f0aaf0aa)
  ) CLBLM_R_X7Y141_SLICE_X9Y141_ALUT (
.I0(CLBLM_L_X10Y130_SLICE_X12Y130_B5Q),
.I1(1'b1),
.I2(CLBLM_L_X10Y133_SLICE_X12Y133_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y135_SLICE_X9Y135_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y141_SLICE_X9Y141_AO5),
.O6(CLBLM_R_X7Y141_SLICE_X9Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y142_SLICE_X8Y142_DO5),
.O6(CLBLM_R_X7Y142_SLICE_X8Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y142_SLICE_X8Y142_CO5),
.O6(CLBLM_R_X7Y142_SLICE_X8Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y142_SLICE_X8Y142_BO5),
.O6(CLBLM_R_X7Y142_SLICE_X8Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y142_SLICE_X8Y142_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y142_SLICE_X8Y142_AO5),
.O6(CLBLM_R_X7Y142_SLICE_X8Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X9Y142_AO6),
.Q(CLBLM_R_X7Y142_SLICE_X9Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X9Y142_BO6),
.Q(CLBLM_R_X7Y142_SLICE_X9Y142_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y142_SLICE_X9Y142_CO6),
.Q(CLBLM_R_X7Y142_SLICE_X9Y142_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4e4f0000000)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_DLUT (
.I0(LIOB33_X0Y61_IOB_X0Y62_I),
.I1(CLBLM_R_X3Y140_SLICE_X3Y140_CQ),
.I2(CLBLM_R_X7Y142_SLICE_X9Y142_BQ),
.I3(CLBLM_R_X7Y142_SLICE_X9Y142_AQ),
.I4(CLBLM_L_X8Y142_SLICE_X10Y142_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y142_SLICE_X9Y142_DO5),
.O6(CLBLM_R_X7Y142_SLICE_X9Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa003caaaa00cc)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_CLUT (
.I0(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I1(CLBLM_R_X7Y142_SLICE_X9Y142_CQ),
.I2(CLBLM_L_X8Y141_SLICE_X11Y141_AQ),
.I3(CLBLM_R_X5Y140_SLICE_X7Y140_A5Q),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X10Y134_SLICE_X12Y134_AQ),
.O5(CLBLM_R_X7Y142_SLICE_X9Y142_CO5),
.O6(CLBLM_R_X7Y142_SLICE_X9Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafafa3aca3ac)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_BLUT (
.I0(CLBLL_L_X4Y138_SLICE_X5Y138_DQ),
.I1(CLBLM_R_X7Y142_SLICE_X9Y142_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X8Y142_SLICE_X10Y142_CO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y140_SLICE_X7Y140_A5Q),
.O5(CLBLM_R_X7Y142_SLICE_X9Y142_BO5),
.O6(CLBLM_R_X7Y142_SLICE_X9Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ffffff007878)
  ) CLBLM_R_X7Y142_SLICE_X9Y142_ALUT (
.I0(CLBLM_L_X8Y142_SLICE_X10Y142_CO6),
.I1(CLBLM_R_X7Y142_SLICE_X9Y142_BQ),
.I2(CLBLM_R_X7Y142_SLICE_X9Y142_AQ),
.I3(CLBLL_L_X4Y133_SLICE_X4Y133_BQ),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X5Y140_SLICE_X7Y140_A5Q),
.O5(CLBLM_R_X7Y142_SLICE_X9Y142_AO5),
.O6(CLBLM_R_X7Y142_SLICE_X9Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X8Y143_BO6),
.Q(CLBLM_R_X7Y143_SLICE_X8Y143_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X8Y143_AO6),
.Q(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y143_SLICE_X8Y143_DO5),
.O6(CLBLM_R_X7Y143_SLICE_X8Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y143_SLICE_X8Y143_CO5),
.O6(CLBLM_R_X7Y143_SLICE_X8Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0afc0c00ff00ff)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_BLUT (
.I0(CLBLM_R_X7Y143_SLICE_X9Y143_BO6),
.I1(CLBLM_R_X7Y143_SLICE_X9Y143_DO6),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLL_L_X4Y141_SLICE_X4Y141_AQ),
.I4(CLBLM_R_X7Y143_SLICE_X8Y143_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y143_SLICE_X8Y143_BO5),
.O6(CLBLM_R_X7Y143_SLICE_X8Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haacfaac0aac0aac0)
  ) CLBLM_R_X7Y143_SLICE_X8Y143_ALUT (
.I0(CLBLM_R_X7Y138_SLICE_X8Y138_B5Q),
.I1(CLBLM_R_X7Y143_SLICE_X9Y143_BO6),
.I2(CLBLM_R_X7Y143_SLICE_X8Y143_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X7Y143_SLICE_X8Y143_A5Q),
.I5(CLBLM_R_X7Y143_SLICE_X9Y143_DO6),
.O5(CLBLM_R_X7Y143_SLICE_X8Y143_AO5),
.O6(CLBLM_R_X7Y143_SLICE_X8Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y143_SLICE_X9Y143_AO6),
.Q(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000400000)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_DLUT (
.I0(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.I1(CLBLM_R_X7Y133_SLICE_X8Y133_A5Q),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_BO5),
.I4(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I5(CLBLM_L_X8Y141_SLICE_X11Y141_BQ),
.O5(CLBLM_R_X7Y143_SLICE_X9Y143_DO5),
.O6(CLBLM_R_X7Y143_SLICE_X9Y143_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccffff0040ffff)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_CLUT (
.I0(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.I1(CLBLM_R_X7Y133_SLICE_X8Y133_A5Q),
.I2(CLBLM_L_X8Y141_SLICE_X10Y141_AQ),
.I3(CLBLM_L_X8Y143_SLICE_X10Y143_BO5),
.I4(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I5(CLBLM_L_X8Y141_SLICE_X11Y141_BQ),
.O5(CLBLM_R_X7Y143_SLICE_X9Y143_CO5),
.O6(CLBLM_R_X7Y143_SLICE_X9Y143_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33f3f3f3f3f3)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y133_SLICE_X8Y133_A5Q),
.I2(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.I3(CLBLM_L_X8Y141_SLICE_X11Y141_BQ),
.I4(CLBLM_L_X8Y143_SLICE_X10Y143_BO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y143_SLICE_X9Y143_BO5),
.O6(CLBLM_R_X7Y143_SLICE_X9Y143_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0505ccccffff)
  ) CLBLM_R_X7Y143_SLICE_X9Y143_ALUT (
.I0(CLBLM_L_X8Y143_SLICE_X10Y143_CO6),
.I1(CLBLM_L_X8Y132_SLICE_X10Y132_BQ),
.I2(CLBLM_R_X7Y143_SLICE_X9Y143_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_R_X7Y143_SLICE_X9Y143_CO6),
.O5(CLBLM_R_X7Y143_SLICE_X9Y143_AO5),
.O6(CLBLM_R_X7Y143_SLICE_X9Y143_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000080)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_DLUT (
.I0(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I1(CLBLM_L_X10Y132_SLICE_X13Y132_AQ),
.I2(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I3(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I5(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_DO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000100000000)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_CLUT (
.I0(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I2(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I3(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I4(CLBLM_R_X11Y140_SLICE_X14Y140_BO6),
.I5(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_CO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffbf)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_BLUT (
.I0(CLBLM_R_X11Y140_SLICE_X14Y140_BO6),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I2(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I3(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I4(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I5(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_BO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffefffffffdfffff)
  ) CLBLM_R_X11Y131_SLICE_X14Y131_ALUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I1(CLBLM_L_X12Y131_SLICE_X16Y131_AO6),
.I2(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I3(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I4(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y131_SLICE_X14Y131_AO5),
.O6(CLBLM_R_X11Y131_SLICE_X14Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_DO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_CO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_BO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffefffff)
  ) CLBLM_R_X11Y131_SLICE_X15Y131_ALUT (
.I0(CLBLM_L_X8Y134_SLICE_X10Y134_A5Q),
.I1(CLBLM_R_X7Y137_SLICE_X8Y137_CQ),
.I2(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I3(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.I4(CLBLL_L_X4Y136_SLICE_X5Y136_D5Q),
.I5(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.O5(CLBLM_R_X11Y131_SLICE_X15Y131_AO5),
.O6(CLBLM_R_X11Y131_SLICE_X15Y131_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y132_SLICE_X14Y132_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X10Y133_SLICE_X12Y133_AQ),
.Q(CLBLM_R_X11Y132_SLICE_X14Y132_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000004000000)
  ) CLBLM_R_X11Y132_SLICE_X14Y132_DLUT (
.I0(CLBLM_L_X12Y131_SLICE_X16Y131_AO6),
.I1(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I2(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I3(CLBLM_L_X10Y140_SLICE_X13Y140_BQ),
.I4(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.O5(CLBLM_R_X11Y132_SLICE_X14Y132_DO5),
.O6(CLBLM_R_X11Y132_SLICE_X14Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffdfddffffcfcc)
  ) CLBLM_R_X11Y132_SLICE_X14Y132_CLUT (
.I0(CLBLM_R_X11Y134_SLICE_X14Y134_AO6),
.I1(CLBLM_L_X10Y132_SLICE_X13Y132_DO6),
.I2(CLBLM_R_X11Y132_SLICE_X15Y132_BO6),
.I3(CLBLM_R_X5Y126_SLICE_X6Y126_A5Q),
.I4(CLBLM_R_X11Y132_SLICE_X14Y132_DO6),
.I5(CLBLM_R_X7Y133_SLICE_X9Y133_CQ),
.O5(CLBLM_R_X11Y132_SLICE_X14Y132_CO5),
.O6(CLBLM_R_X11Y132_SLICE_X14Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3337ffff0005)
  ) CLBLM_R_X11Y132_SLICE_X14Y132_BLUT (
.I0(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I1(CLBLM_R_X11Y132_SLICE_X15Y132_BO6),
.I2(CLBLM_L_X12Y136_SLICE_X17Y136_BO6),
.I3(CLBLM_R_X11Y142_SLICE_X14Y142_AQ),
.I4(CLBLM_R_X11Y132_SLICE_X14Y132_AO6),
.I5(CLBLL_L_X4Y130_SLICE_X4Y130_B5Q),
.O5(CLBLM_R_X11Y132_SLICE_X14Y132_BO5),
.O6(CLBLM_R_X11Y132_SLICE_X14Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000a0088880a00)
  ) CLBLM_R_X11Y132_SLICE_X14Y132_ALUT (
.I0(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_A5Q),
.I2(CLBLM_R_X11Y131_SLICE_X15Y131_AO6),
.I3(CLBLM_L_X8Y132_SLICE_X10Y132_AQ),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I5(CLBLM_L_X12Y132_SLICE_X16Y132_BO6),
.O5(CLBLM_R_X11Y132_SLICE_X14Y132_AO5),
.O6(CLBLM_R_X11Y132_SLICE_X14Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5000303050000000)
  ) CLBLM_R_X11Y132_SLICE_X15Y132_DLUT (
.I0(CLBLM_R_X11Y132_SLICE_X15Y132_AO6),
.I1(CLBLM_R_X11Y131_SLICE_X15Y131_AO6),
.I2(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I3(CLBLL_L_X4Y133_SLICE_X4Y133_D5Q),
.I4(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I5(CLBLM_R_X3Y137_SLICE_X3Y137_C5Q),
.O5(CLBLM_R_X11Y132_SLICE_X15Y132_DO5),
.O6(CLBLM_R_X11Y132_SLICE_X15Y132_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5073ffff5050)
  ) CLBLM_R_X11Y132_SLICE_X15Y132_CLUT (
.I0(CLBLM_R_X11Y134_SLICE_X14Y134_AO6),
.I1(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I2(CLBLM_R_X7Y132_SLICE_X9Y132_DQ),
.I3(CLBLM_L_X12Y136_SLICE_X17Y136_BO6),
.I4(CLBLM_R_X11Y132_SLICE_X15Y132_DO6),
.I5(CLBLL_L_X4Y134_SLICE_X4Y134_C5Q),
.O5(CLBLM_R_X11Y132_SLICE_X15Y132_CO5),
.O6(CLBLM_R_X11Y132_SLICE_X15Y132_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffefffffffff)
  ) CLBLM_R_X11Y132_SLICE_X15Y132_BLUT (
.I0(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.I1(CLBLM_L_X12Y140_SLICE_X16Y140_AO5),
.I2(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I3(CLBLM_L_X8Y134_SLICE_X10Y134_A5Q),
.I4(CLBLM_R_X7Y137_SLICE_X8Y137_CQ),
.I5(CLBLL_L_X4Y136_SLICE_X5Y136_D5Q),
.O5(CLBLM_R_X11Y132_SLICE_X15Y132_BO5),
.O6(CLBLM_R_X11Y132_SLICE_X15Y132_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffdfffffffef)
  ) CLBLM_R_X11Y132_SLICE_X15Y132_ALUT (
.I0(CLBLL_L_X4Y136_SLICE_X5Y136_D5Q),
.I1(CLBLM_R_X7Y137_SLICE_X8Y137_CQ),
.I2(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I3(CLBLM_L_X8Y134_SLICE_X10Y134_A5Q),
.I4(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y132_SLICE_X15Y132_AO5),
.O6(CLBLM_R_X11Y132_SLICE_X15Y132_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y133_SLICE_X14Y133_AO6),
.Q(CLBLM_R_X11Y133_SLICE_X14Y133_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y133_SLICE_X14Y133_BO6),
.Q(CLBLM_R_X11Y133_SLICE_X14Y133_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0035003000050000)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_DLUT (
.I0(CLBLM_L_X12Y132_SLICE_X16Y132_BO6),
.I1(CLBLM_R_X11Y133_SLICE_X15Y133_AO6),
.I2(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I4(CLBLM_R_X5Y133_SLICE_X7Y133_B5Q),
.I5(CLBLM_L_X10Y140_SLICE_X12Y140_D5Q),
.O5(CLBLM_R_X11Y133_SLICE_X14Y133_DO5),
.O6(CLBLM_R_X11Y133_SLICE_X14Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h01000000ffffbfff)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_CLUT (
.I0(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I1(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I2(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I4(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y133_SLICE_X14Y133_CO5),
.O6(CLBLM_R_X11Y133_SLICE_X14Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hacacacacafafa0a0)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_BLUT (
.I0(CLBLM_R_X7Y134_SLICE_X9Y134_CQ),
.I1(CLBLM_R_X11Y133_SLICE_X14Y133_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(1'b1),
.I4(CLBLM_L_X8Y137_SLICE_X10Y137_AQ),
.I5(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.O5(CLBLM_R_X11Y133_SLICE_X14Y133_BO5),
.O6(CLBLM_R_X11Y133_SLICE_X14Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfff0cccc00f0)
  ) CLBLM_R_X11Y133_SLICE_X14Y133_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y133_SLICE_X3Y133_AQ),
.I2(CLBLM_R_X11Y133_SLICE_X14Y133_AQ),
.I3(CLBLM_R_X11Y131_SLICE_X14Y131_BO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLM_L_X10Y133_SLICE_X13Y133_AQ),
.O5(CLBLM_R_X11Y133_SLICE_X14Y133_AO5),
.O6(CLBLM_R_X11Y133_SLICE_X14Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfdfcfcf5f5f0f0)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_DLUT (
.I0(CLBLM_L_X12Y134_SLICE_X17Y134_AO6),
.I1(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.I2(CLBLM_R_X11Y133_SLICE_X14Y133_DO6),
.I3(1'b1),
.I4(CLBLM_R_X7Y134_SLICE_X9Y134_DQ),
.I5(CLBLM_R_X3Y133_SLICE_X3Y133_AQ),
.O5(CLBLM_R_X11Y133_SLICE_X15Y133_DO5),
.O6(CLBLM_R_X11Y133_SLICE_X15Y133_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fcfafef00ccaaee)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_CLUT (
.I0(CLBLM_R_X3Y137_SLICE_X3Y137_C5Q),
.I1(CLBLL_L_X4Y134_SLICE_X4Y134_C5Q),
.I2(CLBLM_R_X11Y132_SLICE_X15Y132_BO6),
.I3(CLBLM_L_X12Y135_SLICE_X17Y135_DO6),
.I4(CLBLM_R_X11Y131_SLICE_X14Y131_AO6),
.I5(CLBLL_L_X4Y133_SLICE_X4Y133_D5Q),
.O5(CLBLM_R_X11Y133_SLICE_X15Y133_CO5),
.O6(CLBLM_R_X11Y133_SLICE_X15Y133_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffcfeffffccee)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_BLUT (
.I0(CLBLM_R_X7Y134_SLICE_X9Y134_DQ),
.I1(CLBLM_R_X11Y133_SLICE_X14Y133_DO6),
.I2(CLBLM_R_X3Y133_SLICE_X3Y133_AQ),
.I3(CLBLM_L_X12Y134_SLICE_X17Y134_AO6),
.I4(CLBLM_L_X10Y137_SLICE_X13Y137_DO6),
.I5(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.O5(CLBLM_R_X11Y133_SLICE_X15Y133_BO5),
.O6(CLBLM_R_X11Y133_SLICE_X15Y133_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffeffffff)
  ) CLBLM_R_X11Y133_SLICE_X15Y133_ALUT (
.I0(CLBLM_L_X8Y134_SLICE_X10Y134_A5Q),
.I1(CLBLM_R_X7Y137_SLICE_X8Y137_CQ),
.I2(CLBLL_L_X4Y136_SLICE_X5Y136_D5Q),
.I3(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I4(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I5(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.O5(CLBLM_R_X11Y133_SLICE_X15Y133_AO5),
.O6(CLBLM_R_X11Y133_SLICE_X15Y133_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff73ff73ff50ff50)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_DLUT (
.I0(CLBLM_L_X12Y134_SLICE_X17Y134_AO6),
.I1(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.I2(CLBLM_L_X8Y133_SLICE_X10Y133_C5Q),
.I3(CLBLM_R_X11Y134_SLICE_X14Y134_AO5),
.I4(1'b1),
.I5(CLBLM_L_X8Y134_SLICE_X11Y134_AQ),
.O5(CLBLM_R_X11Y134_SLICE_X14Y134_DO5),
.O6(CLBLM_R_X11Y134_SLICE_X14Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffc)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y134_SLICE_X12Y134_CO6),
.I2(CLBLM_R_X11Y134_SLICE_X15Y134_BO6),
.I3(CLBLM_L_X10Y139_SLICE_X12Y139_BO6),
.I4(CLBLM_R_X11Y134_SLICE_X14Y134_DO6),
.I5(CLBLM_R_X7Y135_SLICE_X8Y135_BO6),
.O5(CLBLM_R_X11Y134_SLICE_X14Y134_CO5),
.O6(CLBLM_R_X11Y134_SLICE_X14Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffcfccefee)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_BLUT (
.I0(CLBLM_L_X8Y133_SLICE_X10Y133_C5Q),
.I1(CLBLM_R_X7Y135_SLICE_X8Y135_BO6),
.I2(CLBLM_R_X11Y131_SLICE_X14Y131_CO6),
.I3(CLBLM_L_X8Y134_SLICE_X11Y134_AQ),
.I4(CLBLM_L_X12Y134_SLICE_X17Y134_AO6),
.I5(CLBLM_R_X11Y134_SLICE_X14Y134_AO5),
.O5(CLBLM_R_X11Y134_SLICE_X14Y134_BO5),
.O6(CLBLM_R_X11Y134_SLICE_X14Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5f5f00000d08)
  ) CLBLM_R_X11Y134_SLICE_X14Y134_ALUT (
.I0(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I1(CLBLM_L_X10Y140_SLICE_X13Y140_DQ),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I3(CLBLM_L_X10Y134_SLICE_X13Y134_A5Q),
.I4(CLBLM_L_X12Y132_SLICE_X16Y132_BO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y134_SLICE_X14Y134_AO5),
.O6(CLBLM_R_X11Y134_SLICE_X14Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3010200030102000)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_DLUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I1(CLBLM_R_X11Y136_SLICE_X14Y136_CO6),
.I2(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I3(CLBLM_R_X5Y136_SLICE_X6Y136_AQ),
.I4(CLBLM_L_X10Y136_SLICE_X13Y136_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y134_SLICE_X15Y134_DO5),
.O6(CLBLM_R_X11Y134_SLICE_X15Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ffaaffccffee)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_CLUT (
.I0(CLBLM_R_X5Y132_SLICE_X7Y132_AQ),
.I1(CLBLM_L_X10Y134_SLICE_X13Y134_AQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y140_SLICE_X14Y140_BO6),
.I4(CLBLM_R_X11Y133_SLICE_X14Y133_CO6),
.I5(CLBLM_L_X12Y134_SLICE_X16Y134_AO6),
.O5(CLBLM_R_X11Y134_SLICE_X15Y134_CO5),
.O6(CLBLM_R_X11Y134_SLICE_X15Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfffbfbfafffafa)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_BLUT (
.I0(CLBLM_R_X11Y134_SLICE_X15Y134_DO6),
.I1(CLBLM_L_X12Y134_SLICE_X16Y134_AO6),
.I2(CLBLM_R_X11Y140_SLICE_X14Y140_BO6),
.I3(CLBLM_R_X11Y133_SLICE_X14Y133_CO6),
.I4(CLBLM_R_X5Y132_SLICE_X7Y132_AQ),
.I5(CLBLM_L_X10Y134_SLICE_X13Y134_AQ),
.O5(CLBLM_R_X11Y134_SLICE_X15Y134_BO5),
.O6(CLBLM_R_X11Y134_SLICE_X15Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000080)
  ) CLBLM_R_X11Y134_SLICE_X15Y134_ALUT (
.I0(LIOB33_X0Y51_IOB_X0Y52_I),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I2(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I3(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I4(CLBLM_L_X12Y135_SLICE_X17Y135_AO6),
.I5(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.O5(CLBLM_R_X11Y134_SLICE_X15Y134_AO5),
.O6(CLBLM_R_X11Y134_SLICE_X15Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff3bff3bff0aff0a)
  ) CLBLM_R_X11Y135_SLICE_X14Y135_DLUT (
.I0(CLBLM_L_X8Y137_SLICE_X11Y137_DQ),
.I1(CLBLM_R_X11Y133_SLICE_X14Y133_CO5),
.I2(CLBLM_L_X8Y136_SLICE_X11Y136_CO5),
.I3(CLBLM_L_X8Y136_SLICE_X10Y136_CO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y133_SLICE_X8Y133_BQ),
.O5(CLBLM_R_X11Y135_SLICE_X14Y135_DO5),
.O6(CLBLM_R_X11Y135_SLICE_X14Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffa)
  ) CLBLM_R_X11Y135_SLICE_X14Y135_CLUT (
.I0(CLBLM_L_X10Y135_SLICE_X12Y135_CO5),
.I1(1'b1),
.I2(CLBLM_R_X7Y135_SLICE_X8Y135_DO6),
.I3(CLBLM_L_X10Y134_SLICE_X13Y134_CO6),
.I4(CLBLM_R_X11Y135_SLICE_X14Y135_DO6),
.I5(CLBLM_L_X10Y135_SLICE_X13Y135_DO6),
.O5(CLBLM_R_X11Y135_SLICE_X14Y135_CO5),
.O6(CLBLM_R_X11Y135_SLICE_X14Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffbabaffba)
  ) CLBLM_R_X11Y135_SLICE_X14Y135_BLUT (
.I0(CLBLM_R_X7Y135_SLICE_X8Y135_DO6),
.I1(CLBLM_L_X8Y136_SLICE_X11Y136_CO5),
.I2(CLBLM_L_X8Y137_SLICE_X11Y137_DQ),
.I3(CLBLM_R_X7Y133_SLICE_X8Y133_BQ),
.I4(CLBLM_R_X11Y133_SLICE_X14Y133_CO5),
.I5(CLBLM_L_X8Y136_SLICE_X10Y136_CO6),
.O5(CLBLM_R_X11Y135_SLICE_X14Y135_BO5),
.O6(CLBLM_R_X11Y135_SLICE_X14Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffcfff4)
  ) CLBLM_R_X11Y135_SLICE_X14Y135_ALUT (
.I0(CLBLM_L_X12Y137_SLICE_X17Y137_CO6),
.I1(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I2(CLBLM_L_X10Y135_SLICE_X13Y135_BO6),
.I3(CLBLM_R_X11Y135_SLICE_X14Y135_BO6),
.I4(CLBLM_L_X10Y133_SLICE_X13Y133_DO6),
.I5(CLBLM_L_X10Y134_SLICE_X13Y134_CO6),
.O5(CLBLM_R_X11Y135_SLICE_X14Y135_AO5),
.O6(CLBLM_R_X11Y135_SLICE_X14Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55550000ff55ff00)
  ) CLBLM_R_X11Y135_SLICE_X15Y135_DLUT (
.I0(CLBLM_L_X12Y135_SLICE_X16Y135_AO6),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X8Y137_SLICE_X10Y137_BQ),
.I4(CLBLM_R_X3Y140_SLICE_X3Y140_C5Q),
.I5(CLBLM_L_X8Y136_SLICE_X11Y136_CO5),
.O5(CLBLM_R_X11Y135_SLICE_X15Y135_DO5),
.O6(CLBLM_R_X11Y135_SLICE_X15Y135_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffc)
  ) CLBLM_R_X11Y135_SLICE_X15Y135_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y135_SLICE_X13Y135_AO6),
.I2(CLBLM_L_X10Y134_SLICE_X13Y134_DO6),
.I3(CLBLM_R_X11Y133_SLICE_X15Y133_DO6),
.I4(CLBLM_R_X11Y135_SLICE_X15Y135_DO6),
.I5(CLBLM_L_X10Y137_SLICE_X13Y137_DO6),
.O5(CLBLM_R_X11Y135_SLICE_X15Y135_CO5),
.O6(CLBLM_R_X11Y135_SLICE_X15Y135_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffcfcffffecfc)
  ) CLBLM_R_X11Y135_SLICE_X15Y135_BLUT (
.I0(CLBLM_R_X11Y136_SLICE_X14Y136_DO6),
.I1(CLBLM_R_X11Y133_SLICE_X15Y133_BO6),
.I2(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I3(CLBLM_L_X12Y137_SLICE_X16Y137_BO6),
.I4(CLBLM_L_X12Y135_SLICE_X16Y135_BO6),
.I5(CLBLM_L_X10Y131_SLICE_X13Y131_DO6),
.O5(CLBLM_R_X11Y135_SLICE_X15Y135_BO5),
.O6(CLBLM_R_X11Y135_SLICE_X15Y135_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff2fff2fffffff2)
  ) CLBLM_R_X11Y135_SLICE_X15Y135_ALUT (
.I0(CLBLM_L_X10Y136_SLICE_X13Y136_AQ),
.I1(CLBLM_L_X12Y136_SLICE_X17Y136_AO6),
.I2(CLBLM_L_X10Y134_SLICE_X12Y134_CO6),
.I3(CLBLM_R_X11Y134_SLICE_X15Y134_CO6),
.I4(CLBLM_R_X5Y136_SLICE_X6Y136_AQ),
.I5(CLBLM_R_X11Y136_SLICE_X15Y136_AO5),
.O5(CLBLM_R_X11Y135_SLICE_X15Y135_AO5),
.O6(CLBLM_R_X11Y135_SLICE_X15Y135_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y136_SLICE_X14Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y136_SLICE_X14Y136_AO6),
.Q(CLBLM_R_X11Y136_SLICE_X14Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h303030ff30303030)
  ) CLBLM_R_X11Y136_SLICE_X14Y136_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y134_SLICE_X14Y134_AO6),
.I2(CLBLM_R_X7Y133_SLICE_X9Y133_CQ),
.I3(CLBLM_L_X12Y136_SLICE_X17Y136_BO6),
.I4(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I5(CLBLM_L_X10Y140_SLICE_X13Y140_BQ),
.O5(CLBLM_R_X11Y136_SLICE_X14Y136_DO5),
.O6(CLBLM_R_X11Y136_SLICE_X14Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffeffff)
  ) CLBLM_R_X11Y136_SLICE_X14Y136_CLUT (
.I0(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I1(CLBLM_R_X7Y137_SLICE_X8Y137_CQ),
.I2(CLBLL_L_X4Y136_SLICE_X5Y136_D5Q),
.I3(CLBLM_L_X8Y134_SLICE_X10Y134_A5Q),
.I4(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I5(CLBLM_L_X10Y135_SLICE_X12Y135_AQ),
.O5(CLBLM_R_X11Y136_SLICE_X14Y136_CO5),
.O6(CLBLM_R_X11Y136_SLICE_X14Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000022223000)
  ) CLBLM_R_X11Y136_SLICE_X14Y136_BLUT (
.I0(CLBLM_R_X11Y140_SLICE_X15Y140_BQ),
.I1(CLBLM_L_X12Y131_SLICE_X16Y131_AO6),
.I2(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I3(CLBLL_L_X4Y140_SLICE_X4Y140_AQ),
.I4(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I5(CLBLM_L_X12Y140_SLICE_X16Y140_AO5),
.O5(CLBLM_R_X11Y136_SLICE_X14Y136_BO5),
.O6(CLBLM_R_X11Y136_SLICE_X14Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaff00f0f0)
  ) CLBLM_R_X11Y136_SLICE_X14Y136_ALUT (
.I0(CLBLM_R_X7Y138_SLICE_X8Y138_CQ),
.I1(1'b1),
.I2(CLBLM_R_X11Y136_SLICE_X14Y136_AQ),
.I3(CLBLM_L_X10Y136_SLICE_X12Y136_AQ),
.I4(CLBLM_R_X13Y134_SLICE_X18Y134_AO6),
.I5(LIOB33_X0Y61_IOB_X0Y62_I),
.O5(CLBLM_R_X11Y136_SLICE_X14Y136_AO5),
.O6(CLBLM_R_X11Y136_SLICE_X14Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y136_SLICE_X15Y136_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X11Y136_SLICE_X14Y136_AQ),
.Q(CLBLM_R_X11Y136_SLICE_X15Y136_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcdcfcdc0323f3d3)
  ) CLBLM_R_X11Y136_SLICE_X15Y136_DLUT (
.I0(CLBLM_R_X11Y138_SLICE_X15Y138_AO6),
.I1(CLBLM_R_X11Y134_SLICE_X14Y134_CO6),
.I2(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I3(CLBLM_L_X10Y136_SLICE_X13Y136_DO6),
.I4(CLBLM_L_X12Y137_SLICE_X16Y137_DO6),
.I5(CLBLM_R_X11Y135_SLICE_X15Y135_CO6),
.O5(CLBLM_R_X11Y136_SLICE_X15Y136_DO5),
.O6(CLBLM_R_X11Y136_SLICE_X15Y136_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000020)
  ) CLBLM_R_X11Y136_SLICE_X15Y136_CLUT (
.I0(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I1(CLBLM_R_X11Y140_SLICE_X14Y140_BO6),
.I2(CLBLL_L_X4Y137_SLICE_X4Y137_AQ),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I4(CLBLM_R_X11Y132_SLICE_X15Y132_AO6),
.I5(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.O5(CLBLM_R_X11Y136_SLICE_X15Y136_CO5),
.O6(CLBLM_R_X11Y136_SLICE_X15Y136_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000070003)
  ) CLBLM_R_X11Y136_SLICE_X15Y136_BLUT (
.I0(CLBLM_L_X10Y136_SLICE_X13Y136_DO6),
.I1(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I2(CLBLM_R_X11Y135_SLICE_X15Y135_AO6),
.I3(CLBLM_R_X11Y134_SLICE_X14Y134_BO6),
.I4(CLBLM_R_X11Y138_SLICE_X15Y138_AO6),
.I5(CLBLM_L_X10Y139_SLICE_X12Y139_BO6),
.O5(CLBLM_R_X11Y136_SLICE_X15Y136_BO5),
.O6(CLBLM_R_X11Y136_SLICE_X15Y136_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffefdffffff)
  ) CLBLM_R_X11Y136_SLICE_X15Y136_ALUT (
.I0(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I1(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I2(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I3(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I4(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y136_SLICE_X15Y136_AO5),
.O6(CLBLM_R_X11Y136_SLICE_X15Y136_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9669966969966996)
  ) CLBLM_R_X11Y137_SLICE_X14Y137_DLUT (
.I0(CLBLM_R_X11Y141_SLICE_X14Y141_AQ),
.I1(CLBLL_L_X4Y134_SLICE_X4Y134_C5Q),
.I2(CLBLM_L_X10Y140_SLICE_X13Y140_BQ),
.I3(CLBLM_L_X12Y136_SLICE_X16Y136_A5Q),
.I4(1'b1),
.I5(CLBLM_L_X10Y136_SLICE_X13Y136_CO6),
.O5(CLBLM_R_X11Y137_SLICE_X14Y137_DO5),
.O6(CLBLM_R_X11Y137_SLICE_X14Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X11Y137_SLICE_X14Y137_CLUT (
.I0(CLBLM_L_X10Y134_SLICE_X13Y134_BO6),
.I1(CLBLM_R_X11Y137_SLICE_X15Y137_CO6),
.I2(CLBLM_R_X11Y137_SLICE_X15Y137_DO6),
.I3(CLBLM_R_X11Y137_SLICE_X15Y137_BO6),
.I4(CLBLM_L_X8Y138_SLICE_X11Y138_DO6),
.I5(CLBLM_R_X11Y137_SLICE_X14Y137_BO6),
.O5(CLBLM_R_X11Y137_SLICE_X14Y137_CO5),
.O6(CLBLM_R_X11Y137_SLICE_X14Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000004)
  ) CLBLM_R_X11Y137_SLICE_X14Y137_BLUT (
.I0(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I1(CLBLM_R_X7Y136_SLICE_X8Y136_AQ),
.I2(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I3(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I4(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.O5(CLBLM_R_X11Y137_SLICE_X14Y137_BO5),
.O6(CLBLM_R_X11Y137_SLICE_X14Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000030f0307)
  ) CLBLM_R_X11Y137_SLICE_X14Y137_ALUT (
.I0(CLBLM_R_X11Y138_SLICE_X15Y138_CO6),
.I1(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I2(CLBLM_L_X8Y133_SLICE_X10Y133_DO6),
.I3(CLBLM_R_X11Y132_SLICE_X14Y132_BO6),
.I4(CLBLM_L_X12Y133_SLICE_X17Y133_AO6),
.I5(CLBLM_R_X11Y137_SLICE_X14Y137_CO6),
.O5(CLBLM_R_X11Y137_SLICE_X14Y137_AO5),
.O6(CLBLM_R_X11Y137_SLICE_X14Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000020000)
  ) CLBLM_R_X11Y137_SLICE_X15Y137_DLUT (
.I0(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I1(CLBLM_R_X11Y140_SLICE_X14Y140_BO6),
.I2(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I3(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I4(CLBLM_L_X10Y131_SLICE_X13Y131_AQ),
.I5(CLBLM_L_X10Y137_SLICE_X12Y137_AO6),
.O5(CLBLM_R_X11Y137_SLICE_X15Y137_DO5),
.O6(CLBLM_R_X11Y137_SLICE_X15Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff04ff00ff00)
  ) CLBLM_R_X11Y137_SLICE_X15Y137_CLUT (
.I0(CLBLM_L_X12Y139_SLICE_X16Y139_AO6),
.I1(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I2(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I3(CLBLM_R_X11Y140_SLICE_X14Y140_BO6),
.I4(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I5(CLBLL_L_X4Y139_SLICE_X4Y139_CQ),
.O5(CLBLM_R_X11Y137_SLICE_X15Y137_CO5),
.O6(CLBLM_R_X11Y137_SLICE_X15Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000008)
  ) CLBLM_R_X11Y137_SLICE_X15Y137_BLUT (
.I0(CLBLM_L_X10Y131_SLICE_X12Y131_AQ),
.I1(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I2(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I3(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I4(CLBLM_L_X12Y138_SLICE_X16Y138_AO6),
.I5(CLBLM_R_X11Y140_SLICE_X14Y140_BO6),
.O5(CLBLM_R_X11Y137_SLICE_X15Y137_BO5),
.O6(CLBLM_R_X11Y137_SLICE_X15Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffafffefafafefe)
  ) CLBLM_R_X11Y137_SLICE_X15Y137_ALUT (
.I0(CLBLM_L_X12Y137_SLICE_X17Y137_AO5),
.I1(CLBLM_R_X7Y135_SLICE_X8Y135_BQ),
.I2(CLBLM_R_X11Y134_SLICE_X15Y134_AO6),
.I3(CLBLM_R_X13Y134_SLICE_X18Y134_AO6),
.I4(CLBLM_R_X13Y137_SLICE_X18Y137_AO6),
.I5(CLBLL_L_X4Y131_SLICE_X4Y131_CQ),
.O5(CLBLM_R_X11Y137_SLICE_X15Y137_AO5),
.O6(CLBLM_R_X11Y137_SLICE_X15Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y138_SLICE_X14Y138_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X10Y138_SLICE_X13Y138_AQ),
.Q(CLBLM_R_X11Y138_SLICE_X14Y138_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffefffe)
  ) CLBLM_R_X11Y138_SLICE_X14Y138_DLUT (
.I0(CLBLM_L_X10Y137_SLICE_X12Y137_DO6),
.I1(CLBLM_R_X7Y135_SLICE_X8Y135_CO6),
.I2(CLBLM_L_X10Y137_SLICE_X13Y137_CO6),
.I3(CLBLM_L_X10Y138_SLICE_X12Y138_DO6),
.I4(1'b1),
.I5(CLBLM_R_X11Y138_SLICE_X14Y138_BO6),
.O5(CLBLM_R_X11Y138_SLICE_X14Y138_DO5),
.O6(CLBLM_R_X11Y138_SLICE_X14Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcceeffffcceeccee)
  ) CLBLM_R_X11Y138_SLICE_X14Y138_CLUT (
.I0(CLBLM_L_X10Y134_SLICE_X12Y134_BQ),
.I1(CLBLM_R_X11Y139_SLICE_X14Y139_BO6),
.I2(1'b1),
.I3(CLBLM_L_X8Y136_SLICE_X11Y136_CO5),
.I4(CLBLM_L_X12Y134_SLICE_X17Y134_AO6),
.I5(CLBLM_L_X10Y138_SLICE_X13Y138_AQ),
.O5(CLBLM_R_X11Y138_SLICE_X14Y138_CO5),
.O6(CLBLM_R_X11Y138_SLICE_X14Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0031000000200000)
  ) CLBLM_R_X11Y138_SLICE_X14Y138_BLUT (
.I0(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I1(CLBLM_L_X12Y139_SLICE_X16Y139_AO6),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_BQ),
.I3(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I4(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I5(CLBLM_L_X10Y139_SLICE_X13Y139_CQ),
.O5(CLBLM_R_X11Y138_SLICE_X14Y138_BO5),
.O6(CLBLM_R_X11Y138_SLICE_X14Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff30ffba)
  ) CLBLM_R_X11Y138_SLICE_X14Y138_ALUT (
.I0(CLBLM_L_X10Y139_SLICE_X13Y139_CQ),
.I1(CLBLM_L_X12Y134_SLICE_X17Y134_AO5),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_BQ),
.I3(CLBLM_L_X10Y137_SLICE_X13Y137_CO6),
.I4(CLBLM_L_X12Y134_SLICE_X17Y134_AO6),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_DO6),
.O5(CLBLM_R_X11Y138_SLICE_X14Y138_AO5),
.O6(CLBLM_R_X11Y138_SLICE_X14Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f050f055a50d2d8)
  ) CLBLM_R_X11Y138_SLICE_X15Y138_DLUT (
.I0(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I1(CLBLM_L_X12Y137_SLICE_X17Y137_CO6),
.I2(CLBLM_R_X11Y138_SLICE_X14Y138_DO6),
.I3(CLBLM_L_X12Y138_SLICE_X17Y138_BO6),
.I4(CLBLM_L_X10Y133_SLICE_X13Y133_DO6),
.I5(CLBLM_R_X11Y135_SLICE_X14Y135_CO6),
.O5(CLBLM_R_X11Y138_SLICE_X15Y138_DO5),
.O6(CLBLM_R_X11Y138_SLICE_X15Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffcfffd)
  ) CLBLM_R_X11Y138_SLICE_X15Y138_CLUT (
.I0(CLBLM_L_X12Y138_SLICE_X17Y138_AO6),
.I1(CLBLM_L_X12Y138_SLICE_X16Y138_AO5),
.I2(CLBLM_R_X11Y139_SLICE_X15Y139_AO6),
.I3(CLBLM_R_X11Y136_SLICE_X15Y136_CO6),
.I4(CLBLM_R_X13Y134_SLICE_X18Y134_AO6),
.I5(CLBLM_R_X11Y138_SLICE_X15Y138_BO6),
.O5(CLBLM_R_X11Y138_SLICE_X15Y138_CO5),
.O6(CLBLM_R_X11Y138_SLICE_X15Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0300575503000300)
  ) CLBLM_R_X11Y138_SLICE_X15Y138_BLUT (
.I0(CLBLM_L_X12Y136_SLICE_X17Y136_AO5),
.I1(CLBLM_L_X12Y135_SLICE_X17Y135_CO6),
.I2(CLBLM_L_X12Y138_SLICE_X16Y138_AO6),
.I3(RIOB33_X105Y145_IOB_X1Y145_I),
.I4(CLBLM_L_X12Y131_SLICE_X16Y131_AO6),
.I5(CLBLM_L_X10Y138_SLICE_X12Y138_BQ),
.O5(CLBLM_R_X11Y138_SLICE_X15Y138_BO5),
.O6(CLBLM_R_X11Y138_SLICE_X15Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff11ff00ff01ff00)
  ) CLBLM_R_X11Y138_SLICE_X15Y138_ALUT (
.I0(CLBLM_R_X11Y140_SLICE_X15Y140_DO6),
.I1(CLBLM_L_X12Y139_SLICE_X16Y139_BO6),
.I2(CLBLM_L_X10Y136_SLICE_X12Y136_BQ),
.I3(CLBLM_L_X12Y133_SLICE_X17Y133_AO6),
.I4(CLBLM_L_X12Y135_SLICE_X17Y135_BO6),
.I5(CLBLM_L_X12Y137_SLICE_X17Y137_BO6),
.O5(CLBLM_R_X11Y138_SLICE_X15Y138_AO5),
.O6(CLBLM_R_X11Y138_SLICE_X15Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y139_SLICE_X14Y139_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X11Y140_SLICE_X14Y140_CQ),
.Q(CLBLM_R_X11Y139_SLICE_X14Y139_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2222222f22222222)
  ) CLBLM_R_X11Y139_SLICE_X14Y139_DLUT (
.I0(CLBLM_L_X12Y135_SLICE_X17Y135_BO6),
.I1(CLBLM_L_X12Y139_SLICE_X16Y139_DO6),
.I2(CLBLM_L_X12Y134_SLICE_X17Y134_AO5),
.I3(CLBLL_L_X4Y130_SLICE_X5Y130_DO5),
.I4(CLBLM_L_X8Y139_SLICE_X10Y139_BO6),
.I5(CLBLM_R_X3Y139_SLICE_X3Y139_BO6),
.O5(CLBLM_R_X11Y139_SLICE_X14Y139_DO5),
.O6(CLBLM_R_X11Y139_SLICE_X14Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000003330323)
  ) CLBLM_R_X11Y139_SLICE_X14Y139_CLUT (
.I0(CLBLM_L_X12Y133_SLICE_X17Y133_AO6),
.I1(CLBLM_R_X11Y138_SLICE_X14Y138_CO6),
.I2(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I3(CLBLM_L_X10Y133_SLICE_X13Y133_BO6),
.I4(CLBLM_R_X11Y139_SLICE_X14Y139_DO6),
.I5(CLBLM_L_X10Y139_SLICE_X13Y139_DO6),
.O5(CLBLM_R_X11Y139_SLICE_X14Y139_CO5),
.O6(CLBLM_R_X11Y139_SLICE_X14Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000540000000400)
  ) CLBLM_R_X11Y139_SLICE_X14Y139_BLUT (
.I0(CLBLM_L_X12Y140_SLICE_X16Y140_AO5),
.I1(CLBLM_L_X10Y131_SLICE_X12Y131_BQ),
.I2(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I3(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I4(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I5(CLBLM_R_X7Y140_SLICE_X8Y140_DQ),
.O5(CLBLM_R_X11Y139_SLICE_X14Y139_BO5),
.O6(CLBLM_R_X11Y139_SLICE_X14Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a5a5a5f5f57575)
  ) CLBLM_R_X11Y139_SLICE_X14Y139_ALUT (
.I0(CLBLM_R_X11Y137_SLICE_X14Y137_DO6),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(CLBLM_R_X11Y140_SLICE_X15Y140_B5Q),
.I3(1'b1),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y139_SLICE_X14Y139_AO5),
.O6(CLBLM_R_X11Y139_SLICE_X14Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3322ffff3332ffff)
  ) CLBLM_R_X11Y139_SLICE_X15Y139_DLUT (
.I0(CLBLM_L_X12Y133_SLICE_X17Y133_AO6),
.I1(CLBLM_L_X10Y133_SLICE_X13Y133_BO6),
.I2(CLBLM_R_X3Y139_SLICE_X3Y139_BO6),
.I3(CLBLM_L_X12Y139_SLICE_X16Y139_CO6),
.I4(CLBLM_L_X12Y131_SLICE_X16Y131_BO6),
.I5(CLBLM_L_X8Y139_SLICE_X10Y139_CO6),
.O5(CLBLM_R_X11Y139_SLICE_X15Y139_DO5),
.O6(CLBLM_R_X11Y139_SLICE_X15Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he11e1ee1f00f0ff0)
  ) CLBLM_R_X11Y139_SLICE_X15Y139_CLUT (
.I0(CLBLM_R_X11Y138_SLICE_X14Y138_CO6),
.I1(CLBLM_L_X10Y139_SLICE_X13Y139_DO6),
.I2(CLBLM_L_X12Y136_SLICE_X17Y136_CO6),
.I3(CLBLM_R_X11Y137_SLICE_X14Y137_AO6),
.I4(CLBLM_L_X12Y134_SLICE_X17Y134_DO6),
.I5(CLBLM_R_X11Y139_SLICE_X15Y139_DO6),
.O5(CLBLM_R_X11Y139_SLICE_X15Y139_CO5),
.O6(CLBLM_R_X11Y139_SLICE_X15Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699f0f09966f0f0)
  ) CLBLM_R_X11Y139_SLICE_X15Y139_BLUT (
.I0(CLBLM_R_X7Y139_SLICE_X9Y139_DO6),
.I1(CLBLM_R_X11Y138_SLICE_X15Y138_DO6),
.I2(CLBLM_R_X11Y139_SLICE_X14Y139_AO6),
.I3(CLBLM_R_X11Y136_SLICE_X15Y136_DO6),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(CLBLM_R_X11Y139_SLICE_X15Y139_CO6),
.O5(CLBLM_R_X11Y139_SLICE_X15Y139_BO5),
.O6(CLBLM_R_X11Y139_SLICE_X15Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000000d0008)
  ) CLBLM_R_X11Y139_SLICE_X15Y139_ALUT (
.I0(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I1(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.I2(CLBLM_L_X12Y135_SLICE_X17Y135_AO6),
.I3(CLBLM_L_X10Y137_SLICE_X12Y137_AO6),
.I4(CLBLM_R_X11Y139_SLICE_X14Y139_AQ),
.I5(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.O5(CLBLM_R_X11Y139_SLICE_X15Y139_AO5),
.O6(CLBLM_R_X11Y139_SLICE_X15Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y140_SLICE_X14Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X10Y137_SLICE_X12Y137_AQ),
.Q(CLBLM_R_X11Y140_SLICE_X14Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y140_SLICE_X14Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLL_L_X4Y136_SLICE_X4Y136_BQ),
.Q(CLBLM_R_X11Y140_SLICE_X14Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y140_SLICE_X14Y140_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_R_X5Y140_SLICE_X7Y140_CQ),
.Q(CLBLM_R_X11Y140_SLICE_X14Y140_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y140_SLICE_X14Y140_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(LIOB33_X0Y61_IOB_X0Y62_I),
.D(CLBLM_L_X8Y138_SLICE_X10Y138_A5Q),
.Q(CLBLM_R_X11Y140_SLICE_X14Y140_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y140_SLICE_X14Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y140_SLICE_X14Y140_DO5),
.O6(CLBLM_R_X11Y140_SLICE_X14Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y140_SLICE_X14Y140_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y140_SLICE_X14Y140_CO5),
.O6(CLBLM_R_X11Y140_SLICE_X14Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffefffffefefefe)
  ) CLBLM_R_X11Y140_SLICE_X14Y140_BLUT (
.I0(RIOB33_X105Y129_IOB_X1Y130_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y129_IOB_X1Y129_I),
.I3(CLBLM_L_X10Y138_SLICE_X13Y138_BQ),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y140_SLICE_X14Y140_BO5),
.O6(CLBLM_R_X11Y140_SLICE_X14Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0afaf3333ffff)
  ) CLBLM_R_X11Y140_SLICE_X14Y140_ALUT (
.I0(CLBLM_L_X8Y137_SLICE_X11Y137_DQ),
.I1(CLBLM_L_X10Y139_SLICE_X13Y139_A5Q),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(1'b1),
.I4(CLBLM_R_X11Y139_SLICE_X14Y139_CO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y140_SLICE_X14Y140_AO5),
.O6(CLBLM_R_X11Y140_SLICE_X14Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y140_SLICE_X15Y140_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y140_SLICE_X15Y140_BO5),
.Q(CLBLM_R_X11Y140_SLICE_X15Y140_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y140_SLICE_X15Y140_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y140_SLICE_X15Y140_AO6),
.Q(CLBLM_R_X11Y140_SLICE_X15Y140_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y140_SLICE_X15Y140_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y140_SLICE_X15Y140_BO6),
.Q(CLBLM_R_X11Y140_SLICE_X15Y140_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf2fff2fff2f2f2f2)
  ) CLBLM_R_X11Y140_SLICE_X15Y140_DLUT (
.I0(CLBLM_R_X11Y140_SLICE_X14Y140_AQ),
.I1(CLBLM_R_X13Y137_SLICE_X18Y137_AO6),
.I2(CLBLM_L_X12Y140_SLICE_X16Y140_AO6),
.I3(CLBLM_L_X12Y136_SLICE_X17Y136_BO6),
.I4(1'b1),
.I5(CLBLM_L_X10Y133_SLICE_X12Y133_BQ),
.O5(CLBLM_R_X11Y140_SLICE_X15Y140_DO5),
.O6(CLBLM_R_X11Y140_SLICE_X15Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffffeac0eac0)
  ) CLBLM_R_X11Y140_SLICE_X15Y140_CLUT (
.I0(CLBLM_R_X11Y139_SLICE_X14Y139_AQ),
.I1(CLBLM_R_X7Y135_SLICE_X8Y135_BQ),
.I2(CLBLM_L_X8Y140_SLICE_X10Y140_CQ),
.I3(RIOB33_X105Y145_IOB_X1Y145_I),
.I4(CLBLM_R_X7Y133_SLICE_X8Y133_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y140_SLICE_X15Y140_CO5),
.O6(CLBLM_R_X11Y140_SLICE_X15Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff000f0f0ccf0cc)
  ) CLBLM_R_X11Y140_SLICE_X15Y140_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y139_SLICE_X15Y139_BO6),
.I2(CLBLL_L_X4Y130_SLICE_X5Y130_BQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X11Y140_SLICE_X15Y140_BO5),
.O6(CLBLM_R_X11Y140_SLICE_X15Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccf0ccf0ccfa)
  ) CLBLM_R_X11Y140_SLICE_X15Y140_ALUT (
.I0(CLBLM_R_X11Y139_SLICE_X14Y139_AO6),
.I1(CLBLM_R_X7Y133_SLICE_X9Y133_B5Q),
.I2(CLBLM_R_X11Y140_SLICE_X15Y140_AQ),
.I3(LIOB33_X0Y61_IOB_X0Y62_I),
.I4(CLBLM_R_X11Y140_SLICE_X14Y140_BO5),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X11Y140_SLICE_X15Y140_AO5),
.O6(CLBLM_R_X11Y140_SLICE_X15Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y141_SLICE_X14Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y140_SLICE_X14Y140_AO6),
.Q(CLBLM_R_X11Y141_SLICE_X14Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y141_SLICE_X14Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y141_SLICE_X14Y141_DO5),
.O6(CLBLM_R_X11Y141_SLICE_X14Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y141_SLICE_X14Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y141_SLICE_X14Y141_CO5),
.O6(CLBLM_R_X11Y141_SLICE_X14Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y141_SLICE_X14Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y141_SLICE_X14Y141_BO5),
.O6(CLBLM_R_X11Y141_SLICE_X14Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y141_SLICE_X14Y141_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y141_SLICE_X14Y141_AO5),
.O6(CLBLM_R_X11Y141_SLICE_X14Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y141_SLICE_X15Y141_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y141_SLICE_X15Y141_AO6),
.Q(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y141_SLICE_X15Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y141_SLICE_X15Y141_DO5),
.O6(CLBLM_R_X11Y141_SLICE_X15Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y141_SLICE_X15Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y141_SLICE_X15Y141_CO5),
.O6(CLBLM_R_X11Y141_SLICE_X15Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y141_SLICE_X15Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y141_SLICE_X15Y141_BO5),
.O6(CLBLM_R_X11Y141_SLICE_X15Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcfcfc5c0c5c0)
  ) CLBLM_R_X11Y141_SLICE_X15Y141_ALUT (
.I0(CLBLM_R_X11Y140_SLICE_X14Y140_BO5),
.I1(CLBLM_R_X11Y140_SLICE_X14Y140_BQ),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y138_SLICE_X13Y138_BQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y141_SLICE_X15Y141_AQ),
.O5(CLBLM_R_X11Y141_SLICE_X15Y141_AO5),
.O6(CLBLM_R_X11Y141_SLICE_X15Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y142_SLICE_X14Y142_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y142_SLICE_X14Y142_AO5),
.Q(CLBLM_R_X11Y142_SLICE_X14Y142_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y142_SLICE_X14Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y142_SLICE_X14Y142_DO5),
.O6(CLBLM_R_X11Y142_SLICE_X14Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y142_SLICE_X14Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y142_SLICE_X14Y142_CO5),
.O6(CLBLM_R_X11Y142_SLICE_X14Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y142_SLICE_X14Y142_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y142_SLICE_X14Y142_BO5),
.O6(CLBLM_R_X11Y142_SLICE_X14Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33fff3f30303)
  ) CLBLM_R_X11Y142_SLICE_X14Y142_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y137_SLICE_X14Y137_AO6),
.I2(LIOB33_X0Y61_IOB_X0Y62_I),
.I3(CLBLM_L_X10Y139_SLICE_X13Y139_A5Q),
.I4(CLBLM_R_X5Y143_SLICE_X7Y143_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y142_SLICE_X14Y142_AO5),
.O6(CLBLM_R_X11Y142_SLICE_X14Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y142_SLICE_X15Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y142_SLICE_X15Y142_DO5),
.O6(CLBLM_R_X11Y142_SLICE_X15Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y142_SLICE_X15Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y142_SLICE_X15Y142_CO5),
.O6(CLBLM_R_X11Y142_SLICE_X15Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y142_SLICE_X15Y142_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y142_SLICE_X15Y142_BO5),
.O6(CLBLM_R_X11Y142_SLICE_X15Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haabbaabb0fff0fff)
  ) CLBLM_R_X11Y142_SLICE_X15Y142_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(CLBLL_L_X4Y138_SLICE_X4Y138_AQ),
.I2(CLBLM_R_X11Y136_SLICE_X15Y136_BO6),
.I3(CLBLM_L_X10Y139_SLICE_X13Y139_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y142_SLICE_X15Y142_AO5),
.O6(CLBLM_R_X11Y142_SLICE_X15Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf2fff2f2f2fff2f2)
  ) CLBLM_R_X13Y134_SLICE_X18Y134_DLUT (
.I0(LIOB33_X0Y51_IOB_X0Y51_I),
.I1(CLBLM_R_X13Y138_SLICE_X18Y138_BO6),
.I2(CLBLM_R_X13Y137_SLICE_X18Y137_BO5),
.I3(CLBLM_L_X12Y136_SLICE_X17Y136_BO6),
.I4(CLBLM_R_X7Y131_SLICE_X8Y131_DQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y134_SLICE_X18Y134_DO5),
.O6(CLBLM_R_X13Y134_SLICE_X18Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000002000)
  ) CLBLM_R_X13Y134_SLICE_X18Y134_CLUT (
.I0(LIOB33_X0Y51_IOB_X0Y51_I),
.I1(CLBLM_L_X12Y135_SLICE_X17Y135_AO6),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I3(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I4(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I5(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.O5(CLBLM_R_X13Y134_SLICE_X18Y134_CO5),
.O6(CLBLM_R_X13Y134_SLICE_X18Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000055115011)
  ) CLBLM_R_X13Y134_SLICE_X18Y134_BLUT (
.I0(CLBLM_R_X13Y137_SLICE_X18Y137_BO5),
.I1(CLBLM_R_X7Y131_SLICE_X8Y131_DQ),
.I2(CLBLM_R_X13Y138_SLICE_X18Y138_AO5),
.I3(CLBLM_L_X12Y136_SLICE_X17Y136_BO6),
.I4(CLBLM_R_X13Y134_SLICE_X18Y134_AO6),
.I5(CLBLM_R_X13Y134_SLICE_X18Y134_CO6),
.O5(CLBLM_R_X13Y134_SLICE_X18Y134_BO5),
.O6(CLBLM_R_X13Y134_SLICE_X18Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000400)
  ) CLBLM_R_X13Y134_SLICE_X18Y134_ALUT (
.I0(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I1(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I3(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I4(CLBLM_L_X12Y131_SLICE_X16Y131_AO6),
.I5(CLBLM_R_X11Y140_SLICE_X14Y140_BO6),
.O5(CLBLM_R_X13Y134_SLICE_X18Y134_AO5),
.O6(CLBLM_R_X13Y134_SLICE_X18Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y134_SLICE_X19Y134_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y134_SLICE_X19Y134_DO5),
.O6(CLBLM_R_X13Y134_SLICE_X19Y134_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y134_SLICE_X19Y134_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y134_SLICE_X19Y134_CO5),
.O6(CLBLM_R_X13Y134_SLICE_X19Y134_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y134_SLICE_X19Y134_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y134_SLICE_X19Y134_BO5),
.O6(CLBLM_R_X13Y134_SLICE_X19Y134_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y134_SLICE_X19Y134_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y134_SLICE_X19Y134_AO5),
.O6(CLBLM_R_X13Y134_SLICE_X19Y134_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000000a000a)
  ) CLBLM_R_X13Y137_SLICE_X18Y137_DLUT (
.I0(RIOB33_X105Y143_IOB_X1Y144_I),
.I1(1'b1),
.I2(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I3(CLBLM_L_X12Y135_SLICE_X17Y135_CO6),
.I4(1'b1),
.I5(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.O5(CLBLM_R_X13Y137_SLICE_X18Y137_DO5),
.O6(CLBLM_R_X13Y137_SLICE_X18Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heaeaeaeac0c0c0c0)
  ) CLBLM_R_X13Y137_SLICE_X18Y137_CLUT (
.I0(CLBLM_R_X11Y136_SLICE_X15Y136_AQ),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(CLBLM_L_X10Y137_SLICE_X12Y137_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLM_R_X13Y137_SLICE_X18Y137_CO5),
.O6(CLBLM_R_X13Y137_SLICE_X18Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffddffdd20222000)
  ) CLBLM_R_X13Y137_SLICE_X18Y137_BLUT (
.I0(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I1(CLBLM_L_X12Y135_SLICE_X17Y135_CO6),
.I2(CLBLM_L_X8Y136_SLICE_X10Y136_AQ),
.I3(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I4(RIOB33_X105Y135_IOB_X1Y135_I),
.I5(1'b1),
.O5(CLBLM_R_X13Y137_SLICE_X18Y137_BO5),
.O6(CLBLM_R_X13Y137_SLICE_X18Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff5fff5f00a80008)
  ) CLBLM_R_X13Y137_SLICE_X18Y137_ALUT (
.I0(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I1(RIOB33_X105Y135_IOB_X1Y136_I),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I3(CLBLM_L_X12Y135_SLICE_X17Y135_CO6),
.I4(CLBLM_R_X11Y136_SLICE_X15Y136_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y137_SLICE_X18Y137_AO5),
.O6(CLBLM_R_X13Y137_SLICE_X18Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y137_SLICE_X19Y137_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y137_SLICE_X19Y137_DO5),
.O6(CLBLM_R_X13Y137_SLICE_X19Y137_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y137_SLICE_X19Y137_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y137_SLICE_X19Y137_CO5),
.O6(CLBLM_R_X13Y137_SLICE_X19Y137_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y137_SLICE_X19Y137_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y137_SLICE_X19Y137_BO5),
.O6(CLBLM_R_X13Y137_SLICE_X19Y137_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y137_SLICE_X19Y137_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y137_SLICE_X19Y137_AO5),
.O6(CLBLM_R_X13Y137_SLICE_X19Y137_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y138_SLICE_X18Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y138_SLICE_X18Y138_DO5),
.O6(CLBLM_R_X13Y138_SLICE_X18Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff88ff8888888888)
  ) CLBLM_R_X13Y138_SLICE_X18Y138_CLUT (
.I0(CLBLM_L_X8Y136_SLICE_X10Y136_AQ),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(1'b1),
.I3(RIOB33_X105Y137_IOB_X1Y138_I),
.I4(1'b1),
.I5(CLBLM_L_X8Y139_SLICE_X10Y139_AQ),
.O5(CLBLM_R_X13Y138_SLICE_X18Y138_CO5),
.O6(CLBLM_R_X13Y138_SLICE_X18Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffefffffefefffff)
  ) CLBLM_R_X13Y138_SLICE_X18Y138_BLUT (
.I0(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I1(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I2(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I3(CLBLM_L_X12Y135_SLICE_X17Y135_AO6),
.I4(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y138_SLICE_X18Y138_BO5),
.O6(CLBLM_R_X13Y138_SLICE_X18Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffdff0004030f)
  ) CLBLM_R_X13Y138_SLICE_X18Y138_ALUT (
.I0(CLBLM_R_X5Y136_SLICE_X6Y136_B5Q),
.I1(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.I2(CLBLM_L_X12Y135_SLICE_X17Y135_AO6),
.I3(CLBLM_R_X7Y136_SLICE_X9Y136_AQ),
.I4(CLBLM_R_X3Y136_SLICE_X3Y136_BQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y138_SLICE_X18Y138_AO5),
.O6(CLBLM_R_X13Y138_SLICE_X18Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y138_SLICE_X19Y138_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y138_SLICE_X19Y138_DO5),
.O6(CLBLM_R_X13Y138_SLICE_X19Y138_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y138_SLICE_X19Y138_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y138_SLICE_X19Y138_CO5),
.O6(CLBLM_R_X13Y138_SLICE_X19Y138_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y138_SLICE_X19Y138_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y138_SLICE_X19Y138_BO5),
.O6(CLBLM_R_X13Y138_SLICE_X19Y138_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y138_SLICE_X19Y138_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y138_SLICE_X19Y138_AO5),
.O6(CLBLM_R_X13Y138_SLICE_X19Y138_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X162Y178_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X162Y178_DO5),
.O6(CLBLM_R_X103Y178_SLICE_X162Y178_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X162Y178_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X162Y178_CO5),
.O6(CLBLM_R_X103Y178_SLICE_X162Y178_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X162Y178_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X162Y178_BO5),
.O6(CLBLM_R_X103Y178_SLICE_X162Y178_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X162Y178_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X162Y178_AO5),
.O6(CLBLM_R_X103Y178_SLICE_X162Y178_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X163Y178_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X163Y178_DO5),
.O6(CLBLM_R_X103Y178_SLICE_X163Y178_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X163Y178_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X163Y178_CO5),
.O6(CLBLM_R_X103Y178_SLICE_X163Y178_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y178_SLICE_X163Y178_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y178_SLICE_X163Y178_BO5),
.O6(CLBLM_R_X103Y178_SLICE_X163Y178_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccff00ff00)
  ) CLBLM_R_X103Y178_SLICE_X163Y178_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y125_IOB_X1Y125_I),
.I2(1'b1),
.I3(RIOB33_X105Y125_IOB_X1Y126_I),
.I4(1'b1),
.I5(RIOB33_X105Y127_IOB_X1Y127_I),
.O5(CLBLM_R_X103Y178_SLICE_X163Y178_AO5),
.O6(CLBLM_R_X103Y178_SLICE_X163Y178_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(LIOB33_X0Y77_IOB_X0Y78_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y51_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y51_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y51_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y52_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y52_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y53_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y53_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y53_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y54_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y54_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y55_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y55_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y56_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y56_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y57_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y57_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y57_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y58_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y58_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y59_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y59_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y60_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y60_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y61_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y61_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y62_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y62_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y63_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y63_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y63_IOB_X0Y64_OBUF (
.I(CLBLL_L_X2Y134_SLICE_X1Y134_AO5),
.O(LIOB33_X0Y63_IOB_X0Y64_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y65_IOB_X0Y65_OBUF (
.I(CLBLL_L_X2Y133_SLICE_X1Y133_BO6),
.O(LIOB33_X0Y65_IOB_X0Y65_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y65_IOB_X0Y66_OBUF (
.I(CLBLM_L_X8Y140_SLICE_X10Y140_DQ),
.O(LIOB33_X0Y65_IOB_X0Y66_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y78_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y78_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y78_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y101_OBUF (
.I(CLBLM_R_X3Y136_SLICE_X2Y136_BQ),
.O(LIOB33_X0Y101_IOB_X0Y101_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y102_OBUF (
.I(CLBLM_R_X5Y129_SLICE_X7Y129_BQ),
.O(LIOB33_X0Y101_IOB_X0Y102_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y103_OBUF (
.I(CLBLM_L_X10Y134_SLICE_X12Y134_B5Q),
.O(LIOB33_X0Y103_IOB_X0Y103_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y104_OBUF (
.I(CLBLM_R_X5Y130_SLICE_X7Y130_D5Q),
.O(LIOB33_X0Y103_IOB_X0Y104_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y105_OBUF (
.I(CLBLL_L_X4Y137_SLICE_X5Y137_B5Q),
.O(LIOB33_X0Y105_IOB_X0Y105_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y106_OBUF (
.I(CLBLL_L_X4Y132_SLICE_X5Y132_BQ),
.O(LIOB33_X0Y105_IOB_X0Y106_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y107_OBUF (
.I(CLBLM_R_X5Y133_SLICE_X7Y133_CQ),
.O(LIOB33_X0Y107_IOB_X0Y107_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y108_OBUF (
.I(CLBLM_R_X5Y130_SLICE_X6Y130_BQ),
.O(LIOB33_X0Y107_IOB_X0Y108_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y109_OBUF (
.I(CLBLL_L_X4Y130_SLICE_X4Y130_BQ),
.O(LIOB33_X0Y109_IOB_X0Y109_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y110_OBUF (
.I(CLBLM_R_X5Y133_SLICE_X7Y133_BQ),
.O(LIOB33_X0Y109_IOB_X0Y110_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y111_OBUF (
.I(CLBLL_L_X4Y131_SLICE_X4Y131_D5Q),
.O(LIOB33_X0Y111_IOB_X0Y111_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y112_OBUF (
.I(CLBLL_L_X4Y132_SLICE_X5Y132_A5Q),
.O(LIOB33_X0Y111_IOB_X0Y112_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y113_OBUF (
.I(CLBLL_L_X4Y130_SLICE_X4Y130_DQ),
.O(LIOB33_X0Y113_IOB_X0Y113_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y114_OBUF (
.I(CLBLM_R_X3Y141_SLICE_X2Y141_BQ),
.O(LIOB33_X0Y113_IOB_X0Y114_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y115_OBUF (
.I(CLBLM_R_X5Y138_SLICE_X6Y138_B5Q),
.O(LIOB33_X0Y115_IOB_X0Y115_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y116_OBUF (
.I(CLBLM_L_X10Y131_SLICE_X12Y131_D5Q),
.O(LIOB33_X0Y115_IOB_X0Y116_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y117_OBUF (
.I(CLBLM_L_X10Y130_SLICE_X12Y130_B5Q),
.O(LIOB33_X0Y117_IOB_X0Y117_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y118_OBUF (
.I(CLBLM_R_X5Y130_SLICE_X7Y130_CQ),
.O(LIOB33_X0Y117_IOB_X0Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUF (
.I(CLBLM_R_X3Y132_SLICE_X3Y132_BQ),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUF (
.I(CLBLM_R_X5Y138_SLICE_X7Y138_AQ),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUF (
.I(CLBLM_R_X7Y135_SLICE_X9Y135_C5Q),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUF (
.I(CLBLL_L_X4Y136_SLICE_X4Y136_CQ),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUF (
.I(CLBLM_R_X3Y132_SLICE_X3Y132_BQ),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(CLBLM_L_X8Y140_SLICE_X10Y140_DQ),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y125_OBUF (
.I(CLBLM_L_X8Y138_SLICE_X10Y138_CQ),
.O(LIOB33_X0Y125_IOB_X0Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y126_OBUF (
.I(CLBLM_R_X5Y133_SLICE_X7Y133_AQ),
.O(LIOB33_X0Y125_IOB_X0Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y127_OBUF (
.I(CLBLM_L_X10Y140_SLICE_X13Y140_D5Q),
.O(LIOB33_X0Y127_IOB_X0Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y128_OBUF (
.I(CLBLM_L_X10Y130_SLICE_X12Y130_CQ),
.O(LIOB33_X0Y127_IOB_X0Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y129_OBUF (
.I(CLBLM_R_X3Y132_SLICE_X3Y132_BQ),
.O(LIOB33_X0Y129_IOB_X0Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y130_OBUF (
.I(CLBLM_R_X3Y132_SLICE_X3Y132_AQ),
.O(LIOB33_X0Y129_IOB_X0Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y131_OBUF (
.I(CLBLL_L_X2Y75_SLICE_X0Y75_AO6),
.O(LIOB33_X0Y131_IOB_X0Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y132_OBUF (
.I(CLBLM_R_X3Y131_SLICE_X2Y131_AO6),
.O(LIOB33_X0Y131_IOB_X0Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y133_OBUF (
.I(CLBLL_L_X4Y133_SLICE_X4Y133_BO5),
.O(LIOB33_X0Y133_IOB_X0Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y134_OBUF (
.I(CLBLM_R_X3Y132_SLICE_X3Y132_AQ),
.O(LIOB33_X0Y133_IOB_X0Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y135_OBUF (
.I(CLBLM_R_X3Y132_SLICE_X3Y132_AQ),
.O(LIOB33_X0Y135_IOB_X0Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUF (
.I(CLBLM_L_X8Y141_SLICE_X11Y141_BQ),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUF (
.I(CLBLM_R_X7Y137_SLICE_X9Y137_D5Q),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUF (
.I(CLBLM_R_X3Y139_SLICE_X3Y139_A5Q),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUF (
.I(CLBLM_R_X3Y139_SLICE_X2Y139_C5Q),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUF (
.I(CLBLM_R_X3Y137_SLICE_X3Y137_D5Q),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y141_OBUF (
.I(CLBLL_L_X4Y134_SLICE_X5Y134_DQ),
.O(LIOB33_X0Y141_IOB_X0Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y142_OBUF (
.I(CLBLM_R_X3Y132_SLICE_X3Y132_BQ),
.O(LIOB33_X0Y141_IOB_X0Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y143_IOB_X0Y143_OBUF (
.I(CLBLL_L_X4Y138_SLICE_X4Y138_AO5),
.O(LIOB33_X0Y143_IOB_X0Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y145_OBUF (
.I(CLBLM_R_X3Y137_SLICE_X2Y137_DO6),
.O(LIOB33_X0Y145_IOB_X0Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y146_OBUF (
.I(CLBLM_R_X3Y141_SLICE_X3Y141_BO6),
.O(LIOB33_X0Y145_IOB_X0Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y147_OBUF (
.I(CLBLL_L_X4Y139_SLICE_X5Y139_DO5),
.O(LIOB33_X0Y147_IOB_X0Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y148_OBUF (
.I(CLBLL_L_X4Y141_SLICE_X5Y141_DO6),
.O(LIOB33_X0Y147_IOB_X0Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y151_OBUF (
.I(CLBLM_R_X3Y132_SLICE_X3Y132_BQ),
.O(LIOB33_X0Y151_IOB_X0Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y152_OBUF (
.I(CLBLM_R_X5Y133_SLICE_X7Y133_A5Q),
.O(LIOB33_X0Y151_IOB_X0Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y153_OBUF (
.I(CLBLM_L_X10Y140_SLICE_X12Y140_AQ),
.O(LIOB33_X0Y153_IOB_X0Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y154_OBUF (
.I(CLBLM_L_X10Y137_SLICE_X13Y137_AQ),
.O(LIOB33_X0Y153_IOB_X0Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y155_OBUF (
.I(CLBLM_L_X8Y135_SLICE_X11Y135_AQ),
.O(LIOB33_X0Y155_IOB_X0Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y156_OBUF (
.I(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.O(LIOB33_X0Y155_IOB_X0Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y157_OBUF (
.I(CLBLM_R_X3Y140_SLICE_X3Y140_AQ),
.O(LIOB33_X0Y157_IOB_X0Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y158_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_I),
.O(LIOB33_X0Y157_IOB_X0Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y159_OBUF (
.I(CLBLM_R_X3Y132_SLICE_X3Y132_BQ),
.O(LIOB33_X0Y159_IOB_X0Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y160_OBUF (
.I(CLBLM_R_X3Y134_SLICE_X2Y134_AQ),
.O(LIOB33_X0Y159_IOB_X0Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y161_OBUF (
.I(CLBLM_R_X5Y140_SLICE_X6Y140_A5Q),
.O(LIOB33_X0Y161_IOB_X0Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y162_OBUF (
.I(CLBLL_L_X4Y142_SLICE_X5Y142_CO5),
.O(LIOB33_X0Y161_IOB_X0Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y163_OBUF (
.I(CLBLM_R_X5Y140_SLICE_X6Y140_BO5),
.O(LIOB33_X0Y163_IOB_X0Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y164_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_I),
.O(LIOB33_X0Y163_IOB_X0Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y165_OBUF (
.I(LIOB33_X0Y57_IOB_X0Y57_I),
.O(LIOB33_X0Y165_IOB_X0Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y166_OBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O(LIOB33_X0Y165_IOB_X0Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y167_OBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_I),
.O(LIOB33_X0Y167_IOB_X0Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y168_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_I),
.O(LIOB33_X0Y167_IOB_X0Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y169_OBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_I),
.O(LIOB33_X0Y169_IOB_X0Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y170_OBUF (
.I(RIOB33_X105Y117_IOB_X1Y118_I),
.O(LIOB33_X0Y169_IOB_X0Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y171_OBUF (
.I(RIOB33_X105Y119_IOB_X1Y119_I),
.O(LIOB33_X0Y171_IOB_X0Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y172_OBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_I),
.O(LIOB33_X0Y171_IOB_X0Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y173_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_I),
.O(LIOB33_X0Y173_IOB_X0Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y174_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_I),
.O(LIOB33_X0Y173_IOB_X0Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y175_OBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_I),
.O(LIOB33_X0Y175_IOB_X0Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y176_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_I),
.O(LIOB33_X0Y175_IOB_X0Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y177_OBUF (
.I(RIOB33_X105Y123_IOB_X1Y124_I),
.O(LIOB33_X0Y177_IOB_X0Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y178_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_I),
.O(LIOB33_X0Y177_IOB_X0Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y179_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_I),
.O(LIOB33_X0Y179_IOB_X0Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y180_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_I),
.O(LIOB33_X0Y179_IOB_X0Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y181_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_I),
.O(LIOB33_X0Y181_IOB_X0Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y182_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_I),
.O(LIOB33_X0Y181_IOB_X0Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y183_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_I),
.O(LIOB33_X0Y183_IOB_X0Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y184_OBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_I),
.O(LIOB33_X0Y183_IOB_X0Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y185_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_I),
.O(LIOB33_X0Y185_IOB_X0Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y186_OBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_I),
.O(LIOB33_X0Y185_IOB_X0Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y187_OBUF (
.I(CLBLM_R_X3Y135_SLICE_X2Y135_AQ),
.O(LIOB33_X0Y187_IOB_X0Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y188_OBUF (
.I(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.O(LIOB33_X0Y187_IOB_X0Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y189_OBUF (
.I(CLBLM_R_X5Y139_SLICE_X6Y139_BQ),
.O(LIOB33_X0Y189_IOB_X0Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y190_OBUF (
.I(CLBLM_R_X7Y143_SLICE_X8Y143_BO5),
.O(LIOB33_X0Y189_IOB_X0Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y191_OBUF (
.I(CLBLM_R_X3Y133_SLICE_X3Y133_CO6),
.O(LIOB33_X0Y191_IOB_X0Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y192_OBUF (
.I(CLBLM_R_X3Y141_SLICE_X2Y141_AO5),
.O(LIOB33_X0Y191_IOB_X0Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y193_OBUF (
.I(CLBLL_L_X4Y142_SLICE_X4Y142_BO6),
.O(LIOB33_X0Y193_IOB_X0Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y194_OBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_I),
.O(LIOB33_X0Y193_IOB_X0Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y195_OBUF (
.I(CLBLL_L_X4Y140_SLICE_X4Y140_DO6),
.O(LIOB33_X0Y195_IOB_X0Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y196_OBUF (
.I(CLBLL_L_X4Y143_SLICE_X4Y143_AO6),
.O(LIOB33_X0Y195_IOB_X0Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y197_OBUF (
.I(CLBLM_R_X3Y141_SLICE_X2Y141_BO6),
.O(LIOB33_X0Y197_IOB_X0Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y198_OBUF (
.I(1'b1),
.O(LIOB33_X0Y197_IOB_X0Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y50_IOB_X0Y50_IBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_IPAD),
.O(LIOB33_SING_X0Y50_IOB_X0Y50_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y100_IOB_X0Y100_OBUF (
.I(CLBLM_R_X3Y136_SLICE_X2Y136_A5Q),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_I),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y150_IOB_X0Y150_OBUF (
.I(CLBLM_R_X3Y134_SLICE_X2Y134_AO5),
.O(LIOB33_SING_X0Y150_IOB_X0Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y199_IOB_X0Y199_OBUF (
.I(1'b1),
.O(LIOB33_SING_X0Y199_IOB_X0Y199_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y101_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y102_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y103_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y104_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y105_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y105_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y106_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y107_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y108_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y109_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y110_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y111_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y112_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y113_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y114_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y115_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y116_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y117_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y118_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y118_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y119_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y119_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y120_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y121_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y122_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y123_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y124_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y124_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y125_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y126_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y127_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y128_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y129_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y129_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y130_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y130_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y131_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y131_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y131_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y132_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y132_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y133_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y133_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y134_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y134_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y135_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y135_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y135_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y136_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y136_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y136_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y137_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y137_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y137_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y138_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y138_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y138_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y139_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y139_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y139_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y140_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y140_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y140_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y141_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y141_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y141_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y142_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y142_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y142_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y143_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y143_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y143_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y144_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y144_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y144_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y145_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y145_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y145_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y146_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y146_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y146_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y147_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y147_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y147_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y148_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y148_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y151_OBUF (
.I(1'b1),
.O(RIOB33_X105Y151_IOB_X1Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y152_OBUF (
.I(1'b1),
.O(RIOB33_X105Y151_IOB_X1Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y153_OBUF (
.I(1'b1),
.O(RIOB33_X105Y153_IOB_X1Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y154_OBUF (
.I(1'b1),
.O(RIOB33_X105Y153_IOB_X1Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y155_OBUF (
.I(1'b1),
.O(RIOB33_X105Y155_IOB_X1Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y156_OBUF (
.I(1'b1),
.O(RIOB33_X105Y155_IOB_X1Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y157_OBUF (
.I(1'b1),
.O(RIOB33_X105Y157_IOB_X1Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y158_OBUF (
.I(1'b1),
.O(RIOB33_X105Y157_IOB_X1Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y159_OBUF (
.I(1'b1),
.O(RIOB33_X105Y159_IOB_X1Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y160_OBUF (
.I(1'b1),
.O(RIOB33_X105Y159_IOB_X1Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y161_OBUF (
.I(CLBLM_R_X3Y141_SLICE_X3Y141_AO5),
.O(RIOB33_X105Y161_IOB_X1Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y162_OBUF (
.I(CLBLM_R_X7Y140_SLICE_X9Y140_D5Q),
.O(RIOB33_X105Y161_IOB_X1Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y163_OBUF (
.I(CLBLM_R_X7Y136_SLICE_X8Y136_D5Q),
.O(RIOB33_X105Y163_IOB_X1Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y164_OBUF (
.I(CLBLM_L_X10Y141_SLICE_X12Y141_BQ),
.O(RIOB33_X105Y163_IOB_X1Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y165_OBUF (
.I(CLBLM_R_X11Y142_SLICE_X15Y142_AO6),
.O(RIOB33_X105Y165_IOB_X1Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y166_OBUF (
.I(CLBLM_L_X10Y140_SLICE_X12Y140_AQ),
.O(RIOB33_X105Y165_IOB_X1Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y167_OBUF (
.I(CLBLM_L_X10Y137_SLICE_X13Y137_AQ),
.O(RIOB33_X105Y167_IOB_X1Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y168_OBUF (
.I(CLBLM_L_X8Y135_SLICE_X11Y135_AQ),
.O(RIOB33_X105Y167_IOB_X1Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y169_OBUF (
.I(CLBLL_L_X4Y142_SLICE_X5Y142_AQ),
.O(RIOB33_X105Y169_IOB_X1Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y170_OBUF (
.I(CLBLM_R_X3Y140_SLICE_X3Y140_AQ),
.O(RIOB33_X105Y169_IOB_X1Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y171_OBUF (
.I(CLBLM_R_X7Y141_SLICE_X9Y141_BO6),
.O(RIOB33_X105Y171_IOB_X1Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y172_OBUF (
.I(CLBLM_R_X3Y134_SLICE_X2Y134_AQ),
.O(RIOB33_X105Y171_IOB_X1Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y173_OBUF (
.I(CLBLM_R_X5Y140_SLICE_X6Y140_A5Q),
.O(RIOB33_X105Y173_IOB_X1Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y174_OBUF (
.I(CLBLM_R_X5Y140_SLICE_X6Y140_BO5),
.O(RIOB33_X105Y173_IOB_X1Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y175_OBUF (
.I(CLBLL_L_X4Y142_SLICE_X5Y142_CO5),
.O(RIOB33_X105Y175_IOB_X1Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y176_OBUF (
.I(CLBLM_R_X3Y138_SLICE_X3Y138_DO6),
.O(RIOB33_X105Y175_IOB_X1Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y177_OBUF (
.I(CLBLM_L_X8Y140_SLICE_X11Y140_BQ),
.O(RIOB33_X105Y177_IOB_X1Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y178_OBUF (
.I(CLBLM_R_X5Y138_SLICE_X6Y138_AQ),
.O(RIOB33_X105Y177_IOB_X1Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y179_OBUF (
.I(CLBLM_R_X5Y139_SLICE_X6Y139_BQ),
.O(RIOB33_X105Y179_IOB_X1Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y180_OBUF (
.I(CLBLM_R_X3Y135_SLICE_X2Y135_AQ),
.O(RIOB33_X105Y179_IOB_X1Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y181_OBUF (
.I(CLBLM_R_X7Y143_SLICE_X8Y143_BO5),
.O(RIOB33_X105Y181_IOB_X1Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y182_OBUF (
.I(CLBLL_L_X4Y141_SLICE_X5Y141_BO5),
.O(RIOB33_X105Y181_IOB_X1Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y183_OBUF (
.I(1'b0),
.O(RIOB33_X105Y183_IOB_X1Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y184_OBUF (
.I(CLBLL_L_X4Y143_SLICE_X4Y143_AO6),
.O(RIOB33_X105Y183_IOB_X1Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y185_OBUF (
.I(CLBLM_R_X7Y141_SLICE_X8Y141_CO6),
.O(RIOB33_X105Y185_IOB_X1Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y186_OBUF (
.I(CLBLM_R_X7Y141_SLICE_X8Y141_DO6),
.O(RIOB33_X105Y185_IOB_X1Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y187_OBUF (
.I(CLBLM_R_X103Y178_SLICE_X163Y178_AO6),
.O(RIOB33_X105Y187_IOB_X1Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y188_OBUF (
.I(CLBLL_L_X4Y141_SLICE_X5Y141_BO5),
.O(RIOB33_X105Y187_IOB_X1Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y189_OBUF (
.I(CLBLM_R_X103Y178_SLICE_X163Y178_AO6),
.O(RIOB33_X105Y189_IOB_X1Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y190_OBUF (
.I(CLBLM_R_X11Y142_SLICE_X15Y142_AO5),
.O(RIOB33_X105Y189_IOB_X1Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y191_OBUF (
.I(CLBLM_L_X12Y142_SLICE_X16Y142_BO5),
.O(RIOB33_X105Y191_IOB_X1Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y192_OBUF (
.I(CLBLM_L_X12Y142_SLICE_X16Y142_AO6),
.O(RIOB33_X105Y191_IOB_X1Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y193_OBUF (
.I(CLBLM_R_X11Y142_SLICE_X14Y142_AO6),
.O(RIOB33_X105Y193_IOB_X1Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y194_OBUF (
.I(CLBLM_L_X12Y142_SLICE_X16Y142_BO6),
.O(RIOB33_X105Y193_IOB_X1Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y195_OBUF (
.I(CLBLM_L_X12Y143_SLICE_X16Y143_AO6),
.O(RIOB33_X105Y195_IOB_X1Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y196_OBUF (
.I(CLBLM_L_X12Y142_SLICE_X16Y142_AO5),
.O(RIOB33_X105Y195_IOB_X1Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y197_OBUF (
.I(CLBLM_R_X11Y140_SLICE_X14Y140_AO5),
.O(RIOB33_X105Y197_IOB_X1Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y198_OBUF (
.I(CLBLM_L_X12Y143_SLICE_X16Y143_AO5),
.O(RIOB33_X105Y197_IOB_X1Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y100_IOB_X1Y100_IBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_IPAD),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y149_IOB_X1Y149_IBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_IPAD),
.O(RIOB33_SING_X105Y149_IOB_X1Y149_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y150_IOB_X1Y150_OBUF (
.I(1'b1),
.O(RIOB33_SING_X105Y150_IOB_X1Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y199_IOB_X1Y199_OBUF (
.I(CLBLM_L_X8Y138_SLICE_X10Y138_B5Q),
.O(RIOB33_SING_X105Y199_IOB_X1Y199_OPAD)
  );
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A = CLBLL_L_X2Y75_SLICE_X0Y75_AO6;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B = CLBLL_L_X2Y75_SLICE_X0Y75_BO6;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C = CLBLL_L_X2Y75_SLICE_X0Y75_CO6;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D = CLBLL_L_X2Y75_SLICE_X0Y75_DO6;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A = CLBLL_L_X2Y75_SLICE_X1Y75_AO6;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B = CLBLL_L_X2Y75_SLICE_X1Y75_BO6;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C = CLBLL_L_X2Y75_SLICE_X1Y75_CO6;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D = CLBLL_L_X2Y75_SLICE_X1Y75_DO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A = CLBLL_L_X2Y133_SLICE_X0Y133_AO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B = CLBLL_L_X2Y133_SLICE_X0Y133_BO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C = CLBLL_L_X2Y133_SLICE_X0Y133_CO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D = CLBLL_L_X2Y133_SLICE_X0Y133_DO6;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A = CLBLL_L_X2Y133_SLICE_X1Y133_AO6;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B = CLBLL_L_X2Y133_SLICE_X1Y133_BO6;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C = CLBLL_L_X2Y133_SLICE_X1Y133_CO6;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D = CLBLL_L_X2Y133_SLICE_X1Y133_DO6;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_A = CLBLL_L_X2Y134_SLICE_X0Y134_AO6;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_B = CLBLL_L_X2Y134_SLICE_X0Y134_BO6;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_C = CLBLL_L_X2Y134_SLICE_X0Y134_CO6;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_D = CLBLL_L_X2Y134_SLICE_X0Y134_DO6;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_A = CLBLL_L_X2Y134_SLICE_X1Y134_AO6;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_B = CLBLL_L_X2Y134_SLICE_X1Y134_BO6;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_C = CLBLL_L_X2Y134_SLICE_X1Y134_CO6;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_D = CLBLL_L_X2Y134_SLICE_X1Y134_DO6;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_AMUX = CLBLL_L_X2Y134_SLICE_X1Y134_AO5;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A = CLBLL_L_X2Y138_SLICE_X0Y138_AO6;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B = CLBLL_L_X2Y138_SLICE_X0Y138_BO6;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C = CLBLL_L_X2Y138_SLICE_X0Y138_CO6;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D = CLBLL_L_X2Y138_SLICE_X0Y138_DO6;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A = CLBLL_L_X2Y138_SLICE_X1Y138_AO6;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B = CLBLL_L_X2Y138_SLICE_X1Y138_BO6;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C = CLBLL_L_X2Y138_SLICE_X1Y138_CO6;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D = CLBLL_L_X2Y138_SLICE_X1Y138_DO6;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_AMUX = CLBLL_L_X2Y138_SLICE_X1Y138_AO5;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A = CLBLL_L_X4Y129_SLICE_X4Y129_AO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B = CLBLL_L_X4Y129_SLICE_X4Y129_BO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C = CLBLL_L_X4Y129_SLICE_X4Y129_CO6;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D = CLBLL_L_X4Y129_SLICE_X4Y129_DO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A = CLBLL_L_X4Y129_SLICE_X5Y129_AO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B = CLBLL_L_X4Y129_SLICE_X5Y129_BO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C = CLBLL_L_X4Y129_SLICE_X5Y129_CO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D = CLBLL_L_X4Y129_SLICE_X5Y129_DO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A = CLBLL_L_X4Y130_SLICE_X4Y130_AO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B = CLBLL_L_X4Y130_SLICE_X4Y130_BO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C = CLBLL_L_X4Y130_SLICE_X4Y130_CO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D = CLBLL_L_X4Y130_SLICE_X4Y130_DO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_BMUX = CLBLL_L_X4Y130_SLICE_X4Y130_B5Q;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_CMUX = CLBLL_L_X4Y130_SLICE_X4Y130_CO5;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_DMUX = CLBLL_L_X4Y130_SLICE_X4Y130_D5Q;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A = CLBLL_L_X4Y130_SLICE_X5Y130_AO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B = CLBLL_L_X4Y130_SLICE_X5Y130_BO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C = CLBLL_L_X4Y130_SLICE_X5Y130_CO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D = CLBLL_L_X4Y130_SLICE_X5Y130_DO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_AMUX = CLBLL_L_X4Y130_SLICE_X5Y130_A5Q;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_BMUX = CLBLL_L_X4Y130_SLICE_X5Y130_B5Q;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_CMUX = CLBLL_L_X4Y130_SLICE_X5Y130_CO5;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_DMUX = CLBLL_L_X4Y130_SLICE_X5Y130_DO5;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A = CLBLL_L_X4Y131_SLICE_X4Y131_AO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B = CLBLL_L_X4Y131_SLICE_X4Y131_BO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C = CLBLL_L_X4Y131_SLICE_X4Y131_CO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D = CLBLL_L_X4Y131_SLICE_X4Y131_DO6;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_DMUX = CLBLL_L_X4Y131_SLICE_X4Y131_D5Q;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A = CLBLL_L_X4Y131_SLICE_X5Y131_AO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B = CLBLL_L_X4Y131_SLICE_X5Y131_BO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C = CLBLL_L_X4Y131_SLICE_X5Y131_CO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D = CLBLL_L_X4Y131_SLICE_X5Y131_DO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_BMUX = CLBLL_L_X4Y131_SLICE_X5Y131_B5Q;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A = CLBLL_L_X4Y132_SLICE_X4Y132_AO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B = CLBLL_L_X4Y132_SLICE_X4Y132_BO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C = CLBLL_L_X4Y132_SLICE_X4Y132_CO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D = CLBLL_L_X4Y132_SLICE_X4Y132_DO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A = CLBLL_L_X4Y132_SLICE_X5Y132_AO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B = CLBLL_L_X4Y132_SLICE_X5Y132_BO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C = CLBLL_L_X4Y132_SLICE_X5Y132_CO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D = CLBLL_L_X4Y132_SLICE_X5Y132_DO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_AMUX = CLBLL_L_X4Y132_SLICE_X5Y132_A5Q;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_CMUX = CLBLL_L_X4Y132_SLICE_X5Y132_C5Q;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_DMUX = CLBLL_L_X4Y132_SLICE_X5Y132_D5Q;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A = CLBLL_L_X4Y133_SLICE_X4Y133_AO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B = CLBLL_L_X4Y133_SLICE_X4Y133_BO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C = CLBLL_L_X4Y133_SLICE_X4Y133_CO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D = CLBLL_L_X4Y133_SLICE_X4Y133_DO6;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_AMUX = CLBLL_L_X4Y133_SLICE_X4Y133_A5Q;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_BMUX = CLBLL_L_X4Y133_SLICE_X4Y133_BO5;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_CMUX = CLBLL_L_X4Y133_SLICE_X4Y133_C5Q;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_DMUX = CLBLL_L_X4Y133_SLICE_X4Y133_D5Q;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A = CLBLL_L_X4Y133_SLICE_X5Y133_AO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B = CLBLL_L_X4Y133_SLICE_X5Y133_BO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C = CLBLL_L_X4Y133_SLICE_X5Y133_CO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D = CLBLL_L_X4Y133_SLICE_X5Y133_DO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_BMUX = CLBLL_L_X4Y133_SLICE_X5Y133_B5Q;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_CMUX = CLBLL_L_X4Y133_SLICE_X5Y133_C5Q;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_DMUX = CLBLL_L_X4Y133_SLICE_X5Y133_D5Q;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A = CLBLL_L_X4Y134_SLICE_X4Y134_AO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B = CLBLL_L_X4Y134_SLICE_X4Y134_BO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C = CLBLL_L_X4Y134_SLICE_X4Y134_CO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D = CLBLL_L_X4Y134_SLICE_X4Y134_DO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_AMUX = CLBLL_L_X4Y134_SLICE_X4Y134_A5Q;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_CMUX = CLBLL_L_X4Y134_SLICE_X4Y134_C5Q;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_DMUX = CLBLL_L_X4Y134_SLICE_X4Y134_D5Q;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A = CLBLL_L_X4Y134_SLICE_X5Y134_AO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B = CLBLL_L_X4Y134_SLICE_X5Y134_BO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C = CLBLL_L_X4Y134_SLICE_X5Y134_CO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D = CLBLL_L_X4Y134_SLICE_X5Y134_DO6;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_DMUX = CLBLL_L_X4Y134_SLICE_X5Y134_D5Q;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A = CLBLL_L_X4Y135_SLICE_X4Y135_AO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B = CLBLL_L_X4Y135_SLICE_X4Y135_BO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C = CLBLL_L_X4Y135_SLICE_X4Y135_CO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D = CLBLL_L_X4Y135_SLICE_X4Y135_DO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_CMUX = CLBLL_L_X4Y135_SLICE_X4Y135_C5Q;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_DMUX = CLBLL_L_X4Y135_SLICE_X4Y135_D5Q;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A = CLBLL_L_X4Y135_SLICE_X5Y135_AO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B = CLBLL_L_X4Y135_SLICE_X5Y135_BO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C = CLBLL_L_X4Y135_SLICE_X5Y135_CO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D = CLBLL_L_X4Y135_SLICE_X5Y135_DO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_CMUX = CLBLL_L_X4Y135_SLICE_X5Y135_C5Q;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_DMUX = CLBLL_L_X4Y135_SLICE_X5Y135_DO5;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A = CLBLL_L_X4Y136_SLICE_X4Y136_AO6;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B = CLBLL_L_X4Y136_SLICE_X4Y136_BO6;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C = CLBLL_L_X4Y136_SLICE_X4Y136_CO6;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D = CLBLL_L_X4Y136_SLICE_X4Y136_DO6;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_AMUX = CLBLL_L_X4Y136_SLICE_X4Y136_A5Q;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_BMUX = CLBLL_L_X4Y136_SLICE_X4Y136_B5Q;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_DMUX = CLBLL_L_X4Y136_SLICE_X4Y136_D5Q;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A = CLBLL_L_X4Y136_SLICE_X5Y136_AO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B = CLBLL_L_X4Y136_SLICE_X5Y136_BO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C = CLBLL_L_X4Y136_SLICE_X5Y136_CO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D = CLBLL_L_X4Y136_SLICE_X5Y136_DO6;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_DMUX = CLBLL_L_X4Y136_SLICE_X5Y136_D5Q;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A = CLBLL_L_X4Y137_SLICE_X4Y137_AO6;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B = CLBLL_L_X4Y137_SLICE_X4Y137_BO6;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C = CLBLL_L_X4Y137_SLICE_X4Y137_CO6;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D = CLBLL_L_X4Y137_SLICE_X4Y137_DO6;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_CMUX = CLBLL_L_X4Y137_SLICE_X4Y137_C5Q;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_DMUX = CLBLL_L_X4Y137_SLICE_X4Y137_DO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A = CLBLL_L_X4Y137_SLICE_X5Y137_AO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B = CLBLL_L_X4Y137_SLICE_X5Y137_BO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C = CLBLL_L_X4Y137_SLICE_X5Y137_CO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D = CLBLL_L_X4Y137_SLICE_X5Y137_DO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_AMUX = CLBLL_L_X4Y137_SLICE_X5Y137_A5Q;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_BMUX = CLBLL_L_X4Y137_SLICE_X5Y137_B5Q;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_CMUX = CLBLL_L_X4Y137_SLICE_X5Y137_C5Q;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_DMUX = CLBLL_L_X4Y137_SLICE_X5Y137_D5Q;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A = CLBLL_L_X4Y138_SLICE_X4Y138_AO6;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B = CLBLL_L_X4Y138_SLICE_X4Y138_BO6;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C = CLBLL_L_X4Y138_SLICE_X4Y138_CO6;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D = CLBLL_L_X4Y138_SLICE_X4Y138_DO6;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_AMUX = CLBLL_L_X4Y138_SLICE_X4Y138_AO5;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_BMUX = CLBLL_L_X4Y138_SLICE_X4Y138_BO5;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A = CLBLL_L_X4Y138_SLICE_X5Y138_AO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B = CLBLL_L_X4Y138_SLICE_X5Y138_BO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C = CLBLL_L_X4Y138_SLICE_X5Y138_CO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D = CLBLL_L_X4Y138_SLICE_X5Y138_DO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_AMUX = CLBLL_L_X4Y138_SLICE_X5Y138_A5Q;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_BMUX = CLBLL_L_X4Y138_SLICE_X5Y138_B5Q;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_CMUX = CLBLL_L_X4Y138_SLICE_X5Y138_C5Q;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_DMUX = CLBLL_L_X4Y138_SLICE_X5Y138_D5Q;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A = CLBLL_L_X4Y139_SLICE_X4Y139_AO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B = CLBLL_L_X4Y139_SLICE_X4Y139_BO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C = CLBLL_L_X4Y139_SLICE_X4Y139_CO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D = CLBLL_L_X4Y139_SLICE_X4Y139_DO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_AMUX = CLBLL_L_X4Y139_SLICE_X4Y139_A5Q;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A = CLBLL_L_X4Y139_SLICE_X5Y139_AO6;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B = CLBLL_L_X4Y139_SLICE_X5Y139_BO6;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C = CLBLL_L_X4Y139_SLICE_X5Y139_CO6;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D = CLBLL_L_X4Y139_SLICE_X5Y139_DO6;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_CMUX = CLBLL_L_X4Y139_SLICE_X5Y139_C5Q;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_DMUX = CLBLL_L_X4Y139_SLICE_X5Y139_DO5;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A = CLBLL_L_X4Y140_SLICE_X4Y140_AO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B = CLBLL_L_X4Y140_SLICE_X4Y140_BO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C = CLBLL_L_X4Y140_SLICE_X4Y140_CO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D = CLBLL_L_X4Y140_SLICE_X4Y140_DO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_AMUX = CLBLL_L_X4Y140_SLICE_X4Y140_AO5;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_BMUX = CLBLL_L_X4Y140_SLICE_X4Y140_BO5;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_CMUX = CLBLL_L_X4Y140_SLICE_X4Y140_CO5;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_DMUX = CLBLL_L_X4Y140_SLICE_X4Y140_DO5;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A = CLBLL_L_X4Y140_SLICE_X5Y140_AO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B = CLBLL_L_X4Y140_SLICE_X5Y140_BO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C = CLBLL_L_X4Y140_SLICE_X5Y140_CO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D = CLBLL_L_X4Y140_SLICE_X5Y140_DO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_CMUX = CLBLL_L_X4Y140_SLICE_X5Y140_C5Q;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A = CLBLL_L_X4Y141_SLICE_X4Y141_AO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B = CLBLL_L_X4Y141_SLICE_X4Y141_BO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C = CLBLL_L_X4Y141_SLICE_X4Y141_CO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D = CLBLL_L_X4Y141_SLICE_X4Y141_DO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A = CLBLL_L_X4Y141_SLICE_X5Y141_AO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B = CLBLL_L_X4Y141_SLICE_X5Y141_BO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C = CLBLL_L_X4Y141_SLICE_X5Y141_CO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D = CLBLL_L_X4Y141_SLICE_X5Y141_DO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_BMUX = CLBLL_L_X4Y141_SLICE_X5Y141_BO5;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A = CLBLL_L_X4Y142_SLICE_X4Y142_AO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B = CLBLL_L_X4Y142_SLICE_X4Y142_BO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C = CLBLL_L_X4Y142_SLICE_X4Y142_CO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D = CLBLL_L_X4Y142_SLICE_X4Y142_DO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_AMUX = CLBLL_L_X4Y142_SLICE_X4Y142_A5Q;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_BMUX = CLBLL_L_X4Y142_SLICE_X4Y142_BO5;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A = CLBLL_L_X4Y142_SLICE_X5Y142_AO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B = CLBLL_L_X4Y142_SLICE_X5Y142_BO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C = CLBLL_L_X4Y142_SLICE_X5Y142_CO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D = CLBLL_L_X4Y142_SLICE_X5Y142_DO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_AMUX = CLBLL_L_X4Y142_SLICE_X5Y142_A5Q;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_CMUX = CLBLL_L_X4Y142_SLICE_X5Y142_CO5;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A = CLBLL_L_X4Y143_SLICE_X4Y143_AO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B = CLBLL_L_X4Y143_SLICE_X4Y143_BO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C = CLBLL_L_X4Y143_SLICE_X4Y143_CO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D = CLBLL_L_X4Y143_SLICE_X4Y143_DO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A = CLBLL_L_X4Y143_SLICE_X5Y143_AO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B = CLBLL_L_X4Y143_SLICE_X5Y143_BO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C = CLBLL_L_X4Y143_SLICE_X5Y143_CO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D = CLBLL_L_X4Y143_SLICE_X5Y143_DO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_BMUX = CLBLL_L_X4Y143_SLICE_X5Y143_BO5;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A = CLBLM_L_X8Y130_SLICE_X10Y130_AO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B = CLBLM_L_X8Y130_SLICE_X10Y130_BO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C = CLBLM_L_X8Y130_SLICE_X10Y130_CO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D = CLBLM_L_X8Y130_SLICE_X10Y130_DO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A = CLBLM_L_X8Y130_SLICE_X11Y130_AO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B = CLBLM_L_X8Y130_SLICE_X11Y130_BO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C = CLBLM_L_X8Y130_SLICE_X11Y130_CO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D = CLBLM_L_X8Y130_SLICE_X11Y130_DO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A = CLBLM_L_X8Y131_SLICE_X10Y131_AO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B = CLBLM_L_X8Y131_SLICE_X10Y131_BO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C = CLBLM_L_X8Y131_SLICE_X10Y131_CO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D = CLBLM_L_X8Y131_SLICE_X10Y131_DO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A = CLBLM_L_X8Y131_SLICE_X11Y131_AO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B = CLBLM_L_X8Y131_SLICE_X11Y131_BO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C = CLBLM_L_X8Y131_SLICE_X11Y131_CO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D = CLBLM_L_X8Y131_SLICE_X11Y131_DO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_CMUX = CLBLM_L_X8Y131_SLICE_X11Y131_C5Q;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_DMUX = CLBLM_L_X8Y131_SLICE_X11Y131_D5Q;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A = CLBLM_L_X8Y132_SLICE_X10Y132_AO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B = CLBLM_L_X8Y132_SLICE_X10Y132_BO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C = CLBLM_L_X8Y132_SLICE_X10Y132_CO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D = CLBLM_L_X8Y132_SLICE_X10Y132_DO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_AMUX = CLBLM_L_X8Y132_SLICE_X10Y132_A5Q;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_BMUX = CLBLM_L_X8Y132_SLICE_X10Y132_B5Q;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A = CLBLM_L_X8Y132_SLICE_X11Y132_AO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B = CLBLM_L_X8Y132_SLICE_X11Y132_BO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C = CLBLM_L_X8Y132_SLICE_X11Y132_CO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D = CLBLM_L_X8Y132_SLICE_X11Y132_DO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_AMUX = CLBLM_L_X8Y132_SLICE_X11Y132_AO5;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_DMUX = CLBLM_L_X8Y132_SLICE_X11Y132_DO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A = CLBLM_L_X8Y133_SLICE_X10Y133_AO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B = CLBLM_L_X8Y133_SLICE_X10Y133_BO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C = CLBLM_L_X8Y133_SLICE_X10Y133_CO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D = CLBLM_L_X8Y133_SLICE_X10Y133_DO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_CMUX = CLBLM_L_X8Y133_SLICE_X10Y133_C5Q;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A = CLBLM_L_X8Y133_SLICE_X11Y133_AO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B = CLBLM_L_X8Y133_SLICE_X11Y133_BO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C = CLBLM_L_X8Y133_SLICE_X11Y133_CO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D = CLBLM_L_X8Y133_SLICE_X11Y133_DO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_AMUX = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_BMUX = CLBLM_L_X8Y133_SLICE_X11Y133_B5Q;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_CMUX = CLBLM_L_X8Y133_SLICE_X11Y133_CO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A = CLBLM_L_X8Y134_SLICE_X10Y134_AO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B = CLBLM_L_X8Y134_SLICE_X10Y134_BO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C = CLBLM_L_X8Y134_SLICE_X10Y134_CO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D = CLBLM_L_X8Y134_SLICE_X10Y134_DO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_AMUX = CLBLM_L_X8Y134_SLICE_X10Y134_A5Q;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_DMUX = CLBLM_L_X8Y134_SLICE_X10Y134_DO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A = CLBLM_L_X8Y134_SLICE_X11Y134_AO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B = CLBLM_L_X8Y134_SLICE_X11Y134_BO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C = CLBLM_L_X8Y134_SLICE_X11Y134_CO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D = CLBLM_L_X8Y134_SLICE_X11Y134_DO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_BMUX = CLBLM_L_X8Y134_SLICE_X11Y134_B5Q;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A = CLBLM_L_X8Y135_SLICE_X10Y135_AO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B = CLBLM_L_X8Y135_SLICE_X10Y135_BO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C = CLBLM_L_X8Y135_SLICE_X10Y135_CO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D = CLBLM_L_X8Y135_SLICE_X10Y135_DO6;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_BMUX = CLBLM_L_X8Y135_SLICE_X10Y135_B5Q;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_CMUX = CLBLM_L_X8Y135_SLICE_X10Y135_C5Q;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_DMUX = CLBLM_L_X8Y135_SLICE_X10Y135_D5Q;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A = CLBLM_L_X8Y135_SLICE_X11Y135_AO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B = CLBLM_L_X8Y135_SLICE_X11Y135_BO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C = CLBLM_L_X8Y135_SLICE_X11Y135_CO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D = CLBLM_L_X8Y135_SLICE_X11Y135_DO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A = CLBLM_L_X8Y136_SLICE_X10Y136_AO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B = CLBLM_L_X8Y136_SLICE_X10Y136_BO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C = CLBLM_L_X8Y136_SLICE_X10Y136_CO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D = CLBLM_L_X8Y136_SLICE_X10Y136_DO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_AMUX = CLBLM_L_X8Y136_SLICE_X10Y136_AO5;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A = CLBLM_L_X8Y136_SLICE_X11Y136_AO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B = CLBLM_L_X8Y136_SLICE_X11Y136_BO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C = CLBLM_L_X8Y136_SLICE_X11Y136_CO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D = CLBLM_L_X8Y136_SLICE_X11Y136_DO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_BMUX = CLBLM_L_X8Y136_SLICE_X11Y136_B5Q;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_CMUX = CLBLM_L_X8Y136_SLICE_X11Y136_CO5;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A = CLBLM_L_X8Y137_SLICE_X10Y137_AO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B = CLBLM_L_X8Y137_SLICE_X10Y137_BO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C = CLBLM_L_X8Y137_SLICE_X10Y137_CO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D = CLBLM_L_X8Y137_SLICE_X10Y137_DO6;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_BMUX = CLBLM_L_X8Y137_SLICE_X10Y137_B5Q;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_CMUX = CLBLM_L_X8Y137_SLICE_X10Y137_C5Q;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_DMUX = CLBLM_L_X8Y137_SLICE_X10Y137_D5Q;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A = CLBLM_L_X8Y137_SLICE_X11Y137_AO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B = CLBLM_L_X8Y137_SLICE_X11Y137_BO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C = CLBLM_L_X8Y137_SLICE_X11Y137_CO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D = CLBLM_L_X8Y137_SLICE_X11Y137_DO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_DMUX = CLBLM_L_X8Y137_SLICE_X11Y137_D5Q;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A = CLBLM_L_X8Y138_SLICE_X10Y138_AO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B = CLBLM_L_X8Y138_SLICE_X10Y138_BO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C = CLBLM_L_X8Y138_SLICE_X10Y138_CO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D = CLBLM_L_X8Y138_SLICE_X10Y138_DO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_AMUX = CLBLM_L_X8Y138_SLICE_X10Y138_A5Q;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_BMUX = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_CMUX = CLBLM_L_X8Y138_SLICE_X10Y138_C5Q;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_DMUX = CLBLM_L_X8Y138_SLICE_X10Y138_D5Q;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A = CLBLM_L_X8Y138_SLICE_X11Y138_AO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B = CLBLM_L_X8Y138_SLICE_X11Y138_BO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C = CLBLM_L_X8Y138_SLICE_X11Y138_CO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D = CLBLM_L_X8Y138_SLICE_X11Y138_DO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_BMUX = CLBLM_L_X8Y138_SLICE_X11Y138_B5Q;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_CMUX = CLBLM_L_X8Y138_SLICE_X11Y138_C5Q;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A = CLBLM_L_X8Y139_SLICE_X10Y139_AO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B = CLBLM_L_X8Y139_SLICE_X10Y139_BO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C = CLBLM_L_X8Y139_SLICE_X10Y139_CO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D = CLBLM_L_X8Y139_SLICE_X10Y139_DO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_BMUX = CLBLM_L_X8Y139_SLICE_X10Y139_BO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A = CLBLM_L_X8Y139_SLICE_X11Y139_AO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B = CLBLM_L_X8Y139_SLICE_X11Y139_BO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C = CLBLM_L_X8Y139_SLICE_X11Y139_CO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D = CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_CMUX = CLBLM_L_X8Y139_SLICE_X11Y139_C5Q;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A = CLBLM_L_X8Y140_SLICE_X10Y140_AO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B = CLBLM_L_X8Y140_SLICE_X10Y140_BO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C = CLBLM_L_X8Y140_SLICE_X10Y140_CO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D = CLBLM_L_X8Y140_SLICE_X10Y140_DO6;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_CMUX = CLBLM_L_X8Y140_SLICE_X10Y140_C5Q;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_DMUX = CLBLM_L_X8Y140_SLICE_X10Y140_D5Q;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A = CLBLM_L_X8Y140_SLICE_X11Y140_AO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B = CLBLM_L_X8Y140_SLICE_X11Y140_BO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C = CLBLM_L_X8Y140_SLICE_X11Y140_CO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D = CLBLM_L_X8Y140_SLICE_X11Y140_DO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_BMUX = CLBLM_L_X8Y140_SLICE_X11Y140_B5Q;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A = CLBLM_L_X8Y141_SLICE_X10Y141_AO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B = CLBLM_L_X8Y141_SLICE_X10Y141_BO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C = CLBLM_L_X8Y141_SLICE_X10Y141_CO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_CMUX = CLBLM_L_X8Y141_SLICE_X10Y141_CO5;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A = CLBLM_L_X8Y141_SLICE_X11Y141_AO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B = CLBLM_L_X8Y141_SLICE_X11Y141_BO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C = CLBLM_L_X8Y141_SLICE_X11Y141_CO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_AMUX = CLBLM_L_X8Y141_SLICE_X11Y141_AO5;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_CMUX = CLBLM_L_X8Y141_SLICE_X11Y141_CO5;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A = CLBLM_L_X8Y142_SLICE_X10Y142_AO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B = CLBLM_L_X8Y142_SLICE_X10Y142_BO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C = CLBLM_L_X8Y142_SLICE_X10Y142_CO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D = CLBLM_L_X8Y142_SLICE_X10Y142_DO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_AMUX = CLBLM_L_X8Y142_SLICE_X10Y142_A5Q;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_BMUX = CLBLM_L_X8Y142_SLICE_X10Y142_BO5;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_CMUX = CLBLM_L_X8Y142_SLICE_X10Y142_CO5;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A = CLBLM_L_X8Y142_SLICE_X11Y142_AO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B = CLBLM_L_X8Y142_SLICE_X11Y142_BO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C = CLBLM_L_X8Y142_SLICE_X11Y142_CO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D = CLBLM_L_X8Y142_SLICE_X11Y142_DO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_CMUX = CLBLM_L_X8Y142_SLICE_X11Y142_CO5;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A = CLBLM_L_X8Y143_SLICE_X10Y143_AO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B = CLBLM_L_X8Y143_SLICE_X10Y143_BO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C = CLBLM_L_X8Y143_SLICE_X10Y143_CO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D = CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_BMUX = CLBLM_L_X8Y143_SLICE_X10Y143_BO5;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A = CLBLM_L_X8Y143_SLICE_X11Y143_AO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B = CLBLM_L_X8Y143_SLICE_X11Y143_BO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C = CLBLM_L_X8Y143_SLICE_X11Y143_CO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D = CLBLM_L_X8Y143_SLICE_X11Y143_DO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A = CLBLM_L_X8Y144_SLICE_X10Y144_AO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B = CLBLM_L_X8Y144_SLICE_X10Y144_BO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C = CLBLM_L_X8Y144_SLICE_X10Y144_CO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D = CLBLM_L_X8Y144_SLICE_X10Y144_DO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A = CLBLM_L_X8Y144_SLICE_X11Y144_AO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B = CLBLM_L_X8Y144_SLICE_X11Y144_BO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C = CLBLM_L_X8Y144_SLICE_X11Y144_CO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D = CLBLM_L_X8Y144_SLICE_X11Y144_DO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A = CLBLM_L_X10Y130_SLICE_X12Y130_AO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B = CLBLM_L_X10Y130_SLICE_X12Y130_BO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C = CLBLM_L_X10Y130_SLICE_X12Y130_CO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D = CLBLM_L_X10Y130_SLICE_X12Y130_DO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_BMUX = CLBLM_L_X10Y130_SLICE_X12Y130_B5Q;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_CMUX = CLBLM_L_X10Y130_SLICE_X12Y130_C5Q;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A = CLBLM_L_X10Y130_SLICE_X13Y130_AO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B = CLBLM_L_X10Y130_SLICE_X13Y130_BO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C = CLBLM_L_X10Y130_SLICE_X13Y130_CO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D = CLBLM_L_X10Y130_SLICE_X13Y130_DO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A = CLBLM_L_X10Y131_SLICE_X12Y131_AO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B = CLBLM_L_X10Y131_SLICE_X12Y131_BO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C = CLBLM_L_X10Y131_SLICE_X12Y131_CO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D = CLBLM_L_X10Y131_SLICE_X12Y131_DO6;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_CMUX = CLBLM_L_X10Y131_SLICE_X12Y131_C5Q;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_DMUX = CLBLM_L_X10Y131_SLICE_X12Y131_D5Q;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A = CLBLM_L_X10Y131_SLICE_X13Y131_AO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B = CLBLM_L_X10Y131_SLICE_X13Y131_BO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C = CLBLM_L_X10Y131_SLICE_X13Y131_CO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D = CLBLM_L_X10Y131_SLICE_X13Y131_DO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A = CLBLM_L_X10Y132_SLICE_X12Y132_AO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B = CLBLM_L_X10Y132_SLICE_X12Y132_BO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C = CLBLM_L_X10Y132_SLICE_X12Y132_CO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D = CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_CMUX = CLBLM_L_X10Y132_SLICE_X12Y132_C5Q;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A = CLBLM_L_X10Y132_SLICE_X13Y132_AO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B = CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C = CLBLM_L_X10Y132_SLICE_X13Y132_CO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D = CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A = CLBLM_L_X10Y133_SLICE_X12Y133_AO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B = CLBLM_L_X10Y133_SLICE_X12Y133_BO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C = CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D = CLBLM_L_X10Y133_SLICE_X12Y133_DO6;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_AMUX = CLBLM_L_X10Y133_SLICE_X12Y133_A5Q;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A = CLBLM_L_X10Y133_SLICE_X13Y133_AO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B = CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C = CLBLM_L_X10Y133_SLICE_X13Y133_CO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A = CLBLM_L_X10Y134_SLICE_X12Y134_AO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B = CLBLM_L_X10Y134_SLICE_X12Y134_BO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C = CLBLM_L_X10Y134_SLICE_X12Y134_CO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D = CLBLM_L_X10Y134_SLICE_X12Y134_DO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_AMUX = CLBLM_L_X10Y134_SLICE_X12Y134_A5Q;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_BMUX = CLBLM_L_X10Y134_SLICE_X12Y134_B5Q;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A = CLBLM_L_X10Y134_SLICE_X13Y134_AO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B = CLBLM_L_X10Y134_SLICE_X13Y134_BO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C = CLBLM_L_X10Y134_SLICE_X13Y134_CO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D = CLBLM_L_X10Y134_SLICE_X13Y134_DO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_AMUX = CLBLM_L_X10Y134_SLICE_X13Y134_A5Q;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A = CLBLM_L_X10Y135_SLICE_X12Y135_AO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B = CLBLM_L_X10Y135_SLICE_X12Y135_BO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C = CLBLM_L_X10Y135_SLICE_X12Y135_CO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_AMUX = CLBLM_L_X10Y135_SLICE_X12Y135_A5Q;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_BMUX = CLBLM_L_X10Y135_SLICE_X12Y135_B5Q;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_CMUX = CLBLM_L_X10Y135_SLICE_X12Y135_CO5;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A = CLBLM_L_X10Y135_SLICE_X13Y135_AO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B = CLBLM_L_X10Y135_SLICE_X13Y135_BO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C = CLBLM_L_X10Y135_SLICE_X13Y135_CO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D = CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A = CLBLM_L_X10Y136_SLICE_X12Y136_AO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B = CLBLM_L_X10Y136_SLICE_X12Y136_BO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C = CLBLM_L_X10Y136_SLICE_X12Y136_CO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D = CLBLM_L_X10Y136_SLICE_X12Y136_DO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_CMUX = CLBLM_L_X10Y136_SLICE_X12Y136_C5Q;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A = CLBLM_L_X10Y136_SLICE_X13Y136_AO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B = CLBLM_L_X10Y136_SLICE_X13Y136_BO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C = CLBLM_L_X10Y136_SLICE_X13Y136_CO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D = CLBLM_L_X10Y136_SLICE_X13Y136_DO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_CMUX = CLBLM_L_X10Y136_SLICE_X13Y136_CO5;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_DMUX = CLBLM_L_X10Y136_SLICE_X13Y136_DO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A = CLBLM_L_X10Y137_SLICE_X12Y137_AO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B = CLBLM_L_X10Y137_SLICE_X12Y137_BO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C = CLBLM_L_X10Y137_SLICE_X12Y137_CO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D = CLBLM_L_X10Y137_SLICE_X12Y137_DO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_AMUX = CLBLM_L_X10Y137_SLICE_X12Y137_AO5;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A = CLBLM_L_X10Y137_SLICE_X13Y137_AO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B = CLBLM_L_X10Y137_SLICE_X13Y137_BO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C = CLBLM_L_X10Y137_SLICE_X13Y137_CO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D = CLBLM_L_X10Y137_SLICE_X13Y137_DO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_AMUX = CLBLM_L_X10Y137_SLICE_X13Y137_A5Q;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_BMUX = CLBLM_L_X10Y137_SLICE_X13Y137_BO5;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A = CLBLM_L_X10Y138_SLICE_X12Y138_AO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B = CLBLM_L_X10Y138_SLICE_X12Y138_BO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C = CLBLM_L_X10Y138_SLICE_X12Y138_CO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D = CLBLM_L_X10Y138_SLICE_X12Y138_DO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A = CLBLM_L_X10Y138_SLICE_X13Y138_AO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B = CLBLM_L_X10Y138_SLICE_X13Y138_BO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C = CLBLM_L_X10Y138_SLICE_X13Y138_CO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D = CLBLM_L_X10Y138_SLICE_X13Y138_DO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A = CLBLM_L_X10Y139_SLICE_X12Y139_AO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B = CLBLM_L_X10Y139_SLICE_X12Y139_BO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C = CLBLM_L_X10Y139_SLICE_X12Y139_CO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D = CLBLM_L_X10Y139_SLICE_X12Y139_DO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_AMUX = CLBLM_L_X10Y139_SLICE_X12Y139_AO5;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A = CLBLM_L_X10Y139_SLICE_X13Y139_AO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B = CLBLM_L_X10Y139_SLICE_X13Y139_BO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C = CLBLM_L_X10Y139_SLICE_X13Y139_CO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D = CLBLM_L_X10Y139_SLICE_X13Y139_DO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_AMUX = CLBLM_L_X10Y139_SLICE_X13Y139_A5Q;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A = CLBLM_L_X10Y140_SLICE_X12Y140_AO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B = CLBLM_L_X10Y140_SLICE_X12Y140_BO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C = CLBLM_L_X10Y140_SLICE_X12Y140_CO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D = CLBLM_L_X10Y140_SLICE_X12Y140_DO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_DMUX = CLBLM_L_X10Y140_SLICE_X12Y140_D5Q;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A = CLBLM_L_X10Y140_SLICE_X13Y140_AO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B = CLBLM_L_X10Y140_SLICE_X13Y140_BO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C = CLBLM_L_X10Y140_SLICE_X13Y140_CO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D = CLBLM_L_X10Y140_SLICE_X13Y140_DO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_BMUX = CLBLM_L_X10Y140_SLICE_X13Y140_B5Q;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_CMUX = CLBLM_L_X10Y140_SLICE_X13Y140_C5Q;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_DMUX = CLBLM_L_X10Y140_SLICE_X13Y140_D5Q;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A = CLBLM_L_X10Y141_SLICE_X12Y141_AO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B = CLBLM_L_X10Y141_SLICE_X12Y141_BO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C = CLBLM_L_X10Y141_SLICE_X12Y141_CO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D = CLBLM_L_X10Y141_SLICE_X12Y141_DO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_CMUX = CLBLM_L_X10Y141_SLICE_X12Y141_C5Q;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_DMUX = CLBLM_L_X10Y141_SLICE_X12Y141_DO5;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A = CLBLM_L_X10Y141_SLICE_X13Y141_AO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B = CLBLM_L_X10Y141_SLICE_X13Y141_BO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C = CLBLM_L_X10Y141_SLICE_X13Y141_CO6;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D = CLBLM_L_X10Y141_SLICE_X13Y141_DO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A = CLBLM_L_X10Y142_SLICE_X12Y142_AO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B = CLBLM_L_X10Y142_SLICE_X12Y142_BO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C = CLBLM_L_X10Y142_SLICE_X12Y142_CO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D = CLBLM_L_X10Y142_SLICE_X12Y142_DO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_BMUX = CLBLM_L_X10Y142_SLICE_X12Y142_BO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A = CLBLM_L_X10Y142_SLICE_X13Y142_AO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B = CLBLM_L_X10Y142_SLICE_X13Y142_BO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C = CLBLM_L_X10Y142_SLICE_X13Y142_CO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D = CLBLM_L_X10Y142_SLICE_X13Y142_DO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A = CLBLM_L_X12Y131_SLICE_X16Y131_AO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C = CLBLM_L_X12Y131_SLICE_X16Y131_CO6;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D = CLBLM_L_X12Y131_SLICE_X16Y131_DO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A = CLBLM_L_X12Y131_SLICE_X17Y131_AO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B = CLBLM_L_X12Y131_SLICE_X17Y131_BO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C = CLBLM_L_X12Y131_SLICE_X17Y131_CO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D = CLBLM_L_X12Y131_SLICE_X17Y131_DO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A = CLBLM_L_X12Y132_SLICE_X16Y132_AO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B = CLBLM_L_X12Y132_SLICE_X16Y132_BO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C = CLBLM_L_X12Y132_SLICE_X16Y132_CO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D = CLBLM_L_X12Y132_SLICE_X16Y132_DO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A = CLBLM_L_X12Y132_SLICE_X17Y132_AO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B = CLBLM_L_X12Y132_SLICE_X17Y132_BO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C = CLBLM_L_X12Y132_SLICE_X17Y132_CO6;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D = CLBLM_L_X12Y132_SLICE_X17Y132_DO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A = CLBLM_L_X12Y133_SLICE_X16Y133_AO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B = CLBLM_L_X12Y133_SLICE_X16Y133_BO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C = CLBLM_L_X12Y133_SLICE_X16Y133_CO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D = CLBLM_L_X12Y133_SLICE_X16Y133_DO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A = CLBLM_L_X12Y133_SLICE_X17Y133_AO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B = CLBLM_L_X12Y133_SLICE_X17Y133_BO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C = CLBLM_L_X12Y133_SLICE_X17Y133_CO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D = CLBLM_L_X12Y133_SLICE_X17Y133_DO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_DMUX = CLBLM_L_X12Y133_SLICE_X17Y133_DO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A = CLBLM_L_X12Y134_SLICE_X16Y134_AO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B = CLBLM_L_X12Y134_SLICE_X16Y134_BO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C = CLBLM_L_X12Y134_SLICE_X16Y134_CO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D = CLBLM_L_X12Y134_SLICE_X16Y134_DO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_AMUX = CLBLM_L_X12Y134_SLICE_X16Y134_AO5;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_DMUX = CLBLM_L_X12Y134_SLICE_X16Y134_DO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A = CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B = CLBLM_L_X12Y134_SLICE_X17Y134_BO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C = CLBLM_L_X12Y134_SLICE_X17Y134_CO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D = CLBLM_L_X12Y134_SLICE_X17Y134_DO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_AMUX = CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_CMUX = CLBLM_L_X12Y134_SLICE_X17Y134_CO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A = CLBLM_L_X12Y135_SLICE_X16Y135_AO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B = CLBLM_L_X12Y135_SLICE_X16Y135_BO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C = CLBLM_L_X12Y135_SLICE_X16Y135_CO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D = CLBLM_L_X12Y135_SLICE_X16Y135_DO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_AMUX = CLBLM_L_X12Y135_SLICE_X16Y135_AO5;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_DMUX = CLBLM_L_X12Y135_SLICE_X16Y135_DO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A = CLBLM_L_X12Y135_SLICE_X17Y135_AO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B = CLBLM_L_X12Y135_SLICE_X17Y135_BO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C = CLBLM_L_X12Y135_SLICE_X17Y135_CO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D = CLBLM_L_X12Y135_SLICE_X17Y135_DO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_AMUX = CLBLM_L_X12Y135_SLICE_X17Y135_AO5;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_A = CLBLM_L_X12Y136_SLICE_X16Y136_AO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_B = CLBLM_L_X12Y136_SLICE_X16Y136_BO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_C = CLBLM_L_X12Y136_SLICE_X16Y136_CO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_D = CLBLM_L_X12Y136_SLICE_X16Y136_DO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_AMUX = CLBLM_L_X12Y136_SLICE_X16Y136_A5Q;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_A = CLBLM_L_X12Y136_SLICE_X17Y136_AO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_B = CLBLM_L_X12Y136_SLICE_X17Y136_BO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_C = CLBLM_L_X12Y136_SLICE_X17Y136_CO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_D = CLBLM_L_X12Y136_SLICE_X17Y136_DO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_AMUX = CLBLM_L_X12Y136_SLICE_X17Y136_AO5;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_BMUX = CLBLM_L_X12Y136_SLICE_X17Y136_BO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_CMUX = CLBLM_L_X12Y136_SLICE_X17Y136_CO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A = CLBLM_L_X12Y137_SLICE_X16Y137_AO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B = CLBLM_L_X12Y137_SLICE_X16Y137_BO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C = CLBLM_L_X12Y137_SLICE_X16Y137_CO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D = CLBLM_L_X12Y137_SLICE_X16Y137_DO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A = CLBLM_L_X12Y137_SLICE_X17Y137_AO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B = CLBLM_L_X12Y137_SLICE_X17Y137_BO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C = CLBLM_L_X12Y137_SLICE_X17Y137_CO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D = CLBLM_L_X12Y137_SLICE_X17Y137_DO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_AMUX = CLBLM_L_X12Y137_SLICE_X17Y137_AO5;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_A = CLBLM_L_X12Y138_SLICE_X16Y138_AO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_B = CLBLM_L_X12Y138_SLICE_X16Y138_BO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_C = CLBLM_L_X12Y138_SLICE_X16Y138_CO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_D = CLBLM_L_X12Y138_SLICE_X16Y138_DO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_AMUX = CLBLM_L_X12Y138_SLICE_X16Y138_AO5;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_A = CLBLM_L_X12Y138_SLICE_X17Y138_AO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_B = CLBLM_L_X12Y138_SLICE_X17Y138_BO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_C = CLBLM_L_X12Y138_SLICE_X17Y138_CO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_D = CLBLM_L_X12Y138_SLICE_X17Y138_DO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_BMUX = CLBLM_L_X12Y138_SLICE_X17Y138_BO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_CMUX = CLBLM_L_X12Y138_SLICE_X17Y138_CO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A = CLBLM_L_X12Y139_SLICE_X16Y139_AO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B = CLBLM_L_X12Y139_SLICE_X16Y139_BO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C = CLBLM_L_X12Y139_SLICE_X16Y139_CO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D = CLBLM_L_X12Y139_SLICE_X16Y139_DO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_AMUX = CLBLM_L_X12Y139_SLICE_X16Y139_AO5;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A = CLBLM_L_X12Y139_SLICE_X17Y139_AO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B = CLBLM_L_X12Y139_SLICE_X17Y139_BO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C = CLBLM_L_X12Y139_SLICE_X17Y139_CO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D = CLBLM_L_X12Y139_SLICE_X17Y139_DO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_BMUX = CLBLM_L_X12Y139_SLICE_X17Y139_BO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_A = CLBLM_L_X12Y140_SLICE_X16Y140_AO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_B = CLBLM_L_X12Y140_SLICE_X16Y140_BO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_C = CLBLM_L_X12Y140_SLICE_X16Y140_CO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_D = CLBLM_L_X12Y140_SLICE_X16Y140_DO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_AMUX = CLBLM_L_X12Y140_SLICE_X16Y140_AO5;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_BMUX = CLBLM_L_X12Y140_SLICE_X16Y140_BO5;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_CMUX = CLBLM_L_X12Y140_SLICE_X16Y140_CO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_A = CLBLM_L_X12Y140_SLICE_X17Y140_AO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_B = CLBLM_L_X12Y140_SLICE_X17Y140_BO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_C = CLBLM_L_X12Y140_SLICE_X17Y140_CO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_D = CLBLM_L_X12Y140_SLICE_X17Y140_DO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_A = CLBLM_L_X12Y141_SLICE_X16Y141_AO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_B = CLBLM_L_X12Y141_SLICE_X16Y141_BO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_C = CLBLM_L_X12Y141_SLICE_X16Y141_CO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_D = CLBLM_L_X12Y141_SLICE_X16Y141_DO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_BMUX = CLBLM_L_X12Y141_SLICE_X16Y141_BO6;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_A = CLBLM_L_X12Y141_SLICE_X17Y141_AO6;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_B = CLBLM_L_X12Y141_SLICE_X17Y141_BO6;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_C = CLBLM_L_X12Y141_SLICE_X17Y141_CO6;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_D = CLBLM_L_X12Y141_SLICE_X17Y141_DO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_A = CLBLM_L_X12Y142_SLICE_X16Y142_AO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_B = CLBLM_L_X12Y142_SLICE_X16Y142_BO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_C = CLBLM_L_X12Y142_SLICE_X16Y142_CO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_D = CLBLM_L_X12Y142_SLICE_X16Y142_DO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_AMUX = CLBLM_L_X12Y142_SLICE_X16Y142_AO5;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_BMUX = CLBLM_L_X12Y142_SLICE_X16Y142_BO5;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_A = CLBLM_L_X12Y142_SLICE_X17Y142_AO6;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_B = CLBLM_L_X12Y142_SLICE_X17Y142_BO6;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_C = CLBLM_L_X12Y142_SLICE_X17Y142_CO6;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_D = CLBLM_L_X12Y142_SLICE_X17Y142_DO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A = CLBLM_L_X12Y143_SLICE_X16Y143_AO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B = CLBLM_L_X12Y143_SLICE_X16Y143_BO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C = CLBLM_L_X12Y143_SLICE_X16Y143_CO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D = CLBLM_L_X12Y143_SLICE_X16Y143_DO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_AMUX = CLBLM_L_X12Y143_SLICE_X16Y143_AO5;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A = CLBLM_L_X12Y143_SLICE_X17Y143_AO6;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B = CLBLM_L_X12Y143_SLICE_X17Y143_BO6;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C = CLBLM_L_X12Y143_SLICE_X17Y143_CO6;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D = CLBLM_L_X12Y143_SLICE_X17Y143_DO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A = CLBLM_R_X3Y130_SLICE_X2Y130_AO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B = CLBLM_R_X3Y130_SLICE_X2Y130_BO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C = CLBLM_R_X3Y130_SLICE_X2Y130_CO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D = CLBLM_R_X3Y130_SLICE_X2Y130_DO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A = CLBLM_R_X3Y130_SLICE_X3Y130_AO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B = CLBLM_R_X3Y130_SLICE_X3Y130_BO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C = CLBLM_R_X3Y130_SLICE_X3Y130_CO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D = CLBLM_R_X3Y130_SLICE_X3Y130_DO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A = CLBLM_R_X3Y131_SLICE_X2Y131_AO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B = CLBLM_R_X3Y131_SLICE_X2Y131_BO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C = CLBLM_R_X3Y131_SLICE_X2Y131_CO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D = CLBLM_R_X3Y131_SLICE_X2Y131_DO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A = CLBLM_R_X3Y131_SLICE_X3Y131_AO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B = CLBLM_R_X3Y131_SLICE_X3Y131_BO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C = CLBLM_R_X3Y131_SLICE_X3Y131_CO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D = CLBLM_R_X3Y131_SLICE_X3Y131_DO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_BMUX = CLBLM_R_X3Y131_SLICE_X3Y131_B5Q;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A = CLBLM_R_X3Y132_SLICE_X2Y132_AO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B = CLBLM_R_X3Y132_SLICE_X2Y132_BO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C = CLBLM_R_X3Y132_SLICE_X2Y132_CO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D = CLBLM_R_X3Y132_SLICE_X2Y132_DO6;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_CMUX = CLBLM_R_X3Y132_SLICE_X2Y132_CO5;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A = CLBLM_R_X3Y132_SLICE_X3Y132_AO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B = CLBLM_R_X3Y132_SLICE_X3Y132_BO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C = CLBLM_R_X3Y132_SLICE_X3Y132_CO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D = CLBLM_R_X3Y132_SLICE_X3Y132_DO6;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_DMUX = CLBLM_R_X3Y132_SLICE_X3Y132_D5Q;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A = CLBLM_R_X3Y133_SLICE_X2Y133_AO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B = CLBLM_R_X3Y133_SLICE_X2Y133_BO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C = CLBLM_R_X3Y133_SLICE_X2Y133_CO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D = CLBLM_R_X3Y133_SLICE_X2Y133_DO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_DMUX = CLBLM_R_X3Y133_SLICE_X2Y133_DO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A = CLBLM_R_X3Y133_SLICE_X3Y133_AO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B = CLBLM_R_X3Y133_SLICE_X3Y133_BO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C = CLBLM_R_X3Y133_SLICE_X3Y133_CO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D = CLBLM_R_X3Y133_SLICE_X3Y133_DO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_BMUX = CLBLM_R_X3Y133_SLICE_X3Y133_B5Q;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_A = CLBLM_R_X3Y134_SLICE_X2Y134_AO6;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_B = CLBLM_R_X3Y134_SLICE_X2Y134_BO6;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_C = CLBLM_R_X3Y134_SLICE_X2Y134_CO6;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_D = CLBLM_R_X3Y134_SLICE_X2Y134_DO6;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_AMUX = CLBLM_R_X3Y134_SLICE_X2Y134_AO5;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_A = CLBLM_R_X3Y134_SLICE_X3Y134_AO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_B = CLBLM_R_X3Y134_SLICE_X3Y134_BO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_C = CLBLM_R_X3Y134_SLICE_X3Y134_CO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_D = CLBLM_R_X3Y134_SLICE_X3Y134_DO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_AMUX = CLBLM_R_X3Y134_SLICE_X3Y134_A5Q;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_A = CLBLM_R_X3Y135_SLICE_X2Y135_AO6;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_B = CLBLM_R_X3Y135_SLICE_X2Y135_BO6;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_C = CLBLM_R_X3Y135_SLICE_X2Y135_CO6;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_D = CLBLM_R_X3Y135_SLICE_X2Y135_DO6;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_A = CLBLM_R_X3Y135_SLICE_X3Y135_AO6;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_B = CLBLM_R_X3Y135_SLICE_X3Y135_BO6;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_C = CLBLM_R_X3Y135_SLICE_X3Y135_CO6;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_D = CLBLM_R_X3Y135_SLICE_X3Y135_DO6;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_AMUX = CLBLM_R_X3Y135_SLICE_X3Y135_A5Q;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_A = CLBLM_R_X3Y136_SLICE_X2Y136_AO6;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_B = CLBLM_R_X3Y136_SLICE_X2Y136_BO6;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_C = CLBLM_R_X3Y136_SLICE_X2Y136_CO6;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_D = CLBLM_R_X3Y136_SLICE_X2Y136_DO6;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_AMUX = CLBLM_R_X3Y136_SLICE_X2Y136_A5Q;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_BMUX = CLBLM_R_X3Y136_SLICE_X2Y136_B5Q;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_A = CLBLM_R_X3Y136_SLICE_X3Y136_AO6;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_B = CLBLM_R_X3Y136_SLICE_X3Y136_BO6;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_C = CLBLM_R_X3Y136_SLICE_X3Y136_CO6;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_D = CLBLM_R_X3Y136_SLICE_X3Y136_DO6;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_BMUX = CLBLM_R_X3Y136_SLICE_X3Y136_B5Q;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_CMUX = CLBLM_R_X3Y136_SLICE_X3Y136_C5Q;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_DMUX = CLBLM_R_X3Y136_SLICE_X3Y136_D5Q;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A = CLBLM_R_X3Y137_SLICE_X2Y137_AO6;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B = CLBLM_R_X3Y137_SLICE_X2Y137_BO6;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C = CLBLM_R_X3Y137_SLICE_X2Y137_CO6;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D = CLBLM_R_X3Y137_SLICE_X2Y137_DO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A = CLBLM_R_X3Y137_SLICE_X3Y137_AO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B = CLBLM_R_X3Y137_SLICE_X3Y137_BO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C = CLBLM_R_X3Y137_SLICE_X3Y137_CO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D = CLBLM_R_X3Y137_SLICE_X3Y137_DO6;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_AMUX = CLBLM_R_X3Y137_SLICE_X3Y137_A5Q;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_BMUX = CLBLM_R_X3Y137_SLICE_X3Y137_B5Q;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_CMUX = CLBLM_R_X3Y137_SLICE_X3Y137_C5Q;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_DMUX = CLBLM_R_X3Y137_SLICE_X3Y137_D5Q;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A = CLBLM_R_X3Y138_SLICE_X2Y138_AO6;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B = CLBLM_R_X3Y138_SLICE_X2Y138_BO6;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C = CLBLM_R_X3Y138_SLICE_X2Y138_CO6;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D = CLBLM_R_X3Y138_SLICE_X2Y138_DO6;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A = CLBLM_R_X3Y138_SLICE_X3Y138_AO6;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B = CLBLM_R_X3Y138_SLICE_X3Y138_BO6;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C = CLBLM_R_X3Y138_SLICE_X3Y138_CO6;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D = CLBLM_R_X3Y138_SLICE_X3Y138_DO6;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_AMUX = CLBLM_R_X3Y138_SLICE_X3Y138_A5Q;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_BMUX = CLBLM_R_X3Y138_SLICE_X3Y138_BO5;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A = CLBLM_R_X3Y139_SLICE_X2Y139_AO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B = CLBLM_R_X3Y139_SLICE_X2Y139_BO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C = CLBLM_R_X3Y139_SLICE_X2Y139_CO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D = CLBLM_R_X3Y139_SLICE_X2Y139_DO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_CMUX = CLBLM_R_X3Y139_SLICE_X2Y139_C5Q;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A = CLBLM_R_X3Y139_SLICE_X3Y139_AO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B = CLBLM_R_X3Y139_SLICE_X3Y139_BO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C = CLBLM_R_X3Y139_SLICE_X3Y139_CO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D = CLBLM_R_X3Y139_SLICE_X3Y139_DO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_AMUX = CLBLM_R_X3Y139_SLICE_X3Y139_A5Q;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_A = CLBLM_R_X3Y140_SLICE_X2Y140_AO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_B = CLBLM_R_X3Y140_SLICE_X2Y140_BO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_C = CLBLM_R_X3Y140_SLICE_X2Y140_CO6;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_D = CLBLM_R_X3Y140_SLICE_X2Y140_DO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_A = CLBLM_R_X3Y140_SLICE_X3Y140_AO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_B = CLBLM_R_X3Y140_SLICE_X3Y140_BO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_C = CLBLM_R_X3Y140_SLICE_X3Y140_CO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_D = CLBLM_R_X3Y140_SLICE_X3Y140_DO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_CMUX = CLBLM_R_X3Y140_SLICE_X3Y140_C5Q;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A = CLBLM_R_X3Y141_SLICE_X2Y141_AO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B = CLBLM_R_X3Y141_SLICE_X2Y141_BO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C = CLBLM_R_X3Y141_SLICE_X2Y141_CO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D = CLBLM_R_X3Y141_SLICE_X2Y141_DO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_AMUX = CLBLM_R_X3Y141_SLICE_X2Y141_AO5;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_BMUX = CLBLM_R_X3Y141_SLICE_X2Y141_BO5;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A = CLBLM_R_X3Y141_SLICE_X3Y141_AO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B = CLBLM_R_X3Y141_SLICE_X3Y141_BO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C = CLBLM_R_X3Y141_SLICE_X3Y141_CO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D = CLBLM_R_X3Y141_SLICE_X3Y141_DO6;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_AMUX = CLBLM_R_X3Y141_SLICE_X3Y141_AO5;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A = CLBLM_R_X5Y126_SLICE_X6Y126_AO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B = CLBLM_R_X5Y126_SLICE_X6Y126_BO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C = CLBLM_R_X5Y126_SLICE_X6Y126_CO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D = CLBLM_R_X5Y126_SLICE_X6Y126_DO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_AMUX = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A = CLBLM_R_X5Y126_SLICE_X7Y126_AO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B = CLBLM_R_X5Y126_SLICE_X7Y126_BO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C = CLBLM_R_X5Y126_SLICE_X7Y126_CO6;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D = CLBLM_R_X5Y126_SLICE_X7Y126_DO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A = CLBLM_R_X5Y127_SLICE_X6Y127_AO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B = CLBLM_R_X5Y127_SLICE_X6Y127_BO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C = CLBLM_R_X5Y127_SLICE_X6Y127_CO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D = CLBLM_R_X5Y127_SLICE_X6Y127_DO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_DMUX = CLBLM_R_X5Y127_SLICE_X6Y127_DO5;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A = CLBLM_R_X5Y127_SLICE_X7Y127_AO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B = CLBLM_R_X5Y127_SLICE_X7Y127_BO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C = CLBLM_R_X5Y127_SLICE_X7Y127_CO6;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D = CLBLM_R_X5Y127_SLICE_X7Y127_DO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A = CLBLM_R_X5Y128_SLICE_X6Y128_AO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B = CLBLM_R_X5Y128_SLICE_X6Y128_BO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C = CLBLM_R_X5Y128_SLICE_X6Y128_CO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D = CLBLM_R_X5Y128_SLICE_X6Y128_DO6;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_CMUX = CLBLM_R_X5Y128_SLICE_X6Y128_CO5;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A = CLBLM_R_X5Y128_SLICE_X7Y128_AO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B = CLBLM_R_X5Y128_SLICE_X7Y128_BO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C = CLBLM_R_X5Y128_SLICE_X7Y128_CO6;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D = CLBLM_R_X5Y128_SLICE_X7Y128_DO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A = CLBLM_R_X5Y129_SLICE_X6Y129_AO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B = CLBLM_R_X5Y129_SLICE_X6Y129_BO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C = CLBLM_R_X5Y129_SLICE_X6Y129_CO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D = CLBLM_R_X5Y129_SLICE_X6Y129_DO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A = CLBLM_R_X5Y129_SLICE_X7Y129_AO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B = CLBLM_R_X5Y129_SLICE_X7Y129_BO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C = CLBLM_R_X5Y129_SLICE_X7Y129_CO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D = CLBLM_R_X5Y129_SLICE_X7Y129_DO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_BMUX = CLBLM_R_X5Y129_SLICE_X7Y129_B5Q;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A = CLBLM_R_X5Y130_SLICE_X6Y130_AO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B = CLBLM_R_X5Y130_SLICE_X6Y130_BO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C = CLBLM_R_X5Y130_SLICE_X6Y130_CO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D = CLBLM_R_X5Y130_SLICE_X6Y130_DO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_BMUX = CLBLM_R_X5Y130_SLICE_X6Y130_B5Q;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A = CLBLM_R_X5Y130_SLICE_X7Y130_AO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B = CLBLM_R_X5Y130_SLICE_X7Y130_BO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C = CLBLM_R_X5Y130_SLICE_X7Y130_CO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D = CLBLM_R_X5Y130_SLICE_X7Y130_DO6;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_DMUX = CLBLM_R_X5Y130_SLICE_X7Y130_D5Q;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A = CLBLM_R_X5Y131_SLICE_X6Y131_AO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B = CLBLM_R_X5Y131_SLICE_X6Y131_BO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C = CLBLM_R_X5Y131_SLICE_X6Y131_CO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D = CLBLM_R_X5Y131_SLICE_X6Y131_DO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_CMUX = CLBLM_R_X5Y131_SLICE_X6Y131_CO5;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A = CLBLM_R_X5Y131_SLICE_X7Y131_AO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B = CLBLM_R_X5Y131_SLICE_X7Y131_BO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C = CLBLM_R_X5Y131_SLICE_X7Y131_CO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D = CLBLM_R_X5Y131_SLICE_X7Y131_DO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_DMUX = CLBLM_R_X5Y131_SLICE_X7Y131_D5Q;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A = CLBLM_R_X5Y132_SLICE_X6Y132_AO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B = CLBLM_R_X5Y132_SLICE_X6Y132_BO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C = CLBLM_R_X5Y132_SLICE_X6Y132_CO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D = CLBLM_R_X5Y132_SLICE_X6Y132_DO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A = CLBLM_R_X5Y132_SLICE_X7Y132_AO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B = CLBLM_R_X5Y132_SLICE_X7Y132_BO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C = CLBLM_R_X5Y132_SLICE_X7Y132_CO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_CMUX = CLBLM_R_X5Y132_SLICE_X7Y132_C5Q;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A = CLBLM_R_X5Y133_SLICE_X6Y133_AO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B = CLBLM_R_X5Y133_SLICE_X6Y133_BO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C = CLBLM_R_X5Y133_SLICE_X6Y133_CO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D = CLBLM_R_X5Y133_SLICE_X6Y133_DO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_AMUX = CLBLM_R_X5Y133_SLICE_X6Y133_A5Q;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_BMUX = CLBLM_R_X5Y133_SLICE_X6Y133_B5Q;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_CMUX = CLBLM_R_X5Y133_SLICE_X6Y133_CO5;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A = CLBLM_R_X5Y133_SLICE_X7Y133_AO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B = CLBLM_R_X5Y133_SLICE_X7Y133_BO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C = CLBLM_R_X5Y133_SLICE_X7Y133_CO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D = CLBLM_R_X5Y133_SLICE_X7Y133_DO6;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_AMUX = CLBLM_R_X5Y133_SLICE_X7Y133_A5Q;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_BMUX = CLBLM_R_X5Y133_SLICE_X7Y133_B5Q;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_CMUX = CLBLM_R_X5Y133_SLICE_X7Y133_C5Q;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A = CLBLM_R_X5Y134_SLICE_X6Y134_AO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B = CLBLM_R_X5Y134_SLICE_X6Y134_BO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C = CLBLM_R_X5Y134_SLICE_X6Y134_CO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D = CLBLM_R_X5Y134_SLICE_X6Y134_DO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_AMUX = CLBLM_R_X5Y134_SLICE_X6Y134_A5Q;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_BMUX = CLBLM_R_X5Y134_SLICE_X6Y134_B5Q;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_CMUX = CLBLM_R_X5Y134_SLICE_X6Y134_C5Q;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A = CLBLM_R_X5Y134_SLICE_X7Y134_AO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B = CLBLM_R_X5Y134_SLICE_X7Y134_BO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C = CLBLM_R_X5Y134_SLICE_X7Y134_CO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D = CLBLM_R_X5Y134_SLICE_X7Y134_DO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_AMUX = CLBLM_R_X5Y134_SLICE_X7Y134_A5Q;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_DMUX = CLBLM_R_X5Y134_SLICE_X7Y134_D5Q;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A = CLBLM_R_X5Y135_SLICE_X6Y135_AO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B = CLBLM_R_X5Y135_SLICE_X6Y135_BO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C = CLBLM_R_X5Y135_SLICE_X6Y135_CO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D = CLBLM_R_X5Y135_SLICE_X6Y135_DO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_AMUX = CLBLM_R_X5Y135_SLICE_X6Y135_A5Q;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_BMUX = CLBLM_R_X5Y135_SLICE_X6Y135_B5Q;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_CMUX = CLBLM_R_X5Y135_SLICE_X6Y135_CO5;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A = CLBLM_R_X5Y135_SLICE_X7Y135_AO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B = CLBLM_R_X5Y135_SLICE_X7Y135_BO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C = CLBLM_R_X5Y135_SLICE_X7Y135_CO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D = CLBLM_R_X5Y135_SLICE_X7Y135_DO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_BMUX = CLBLM_R_X5Y135_SLICE_X7Y135_B5Q;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_DMUX = CLBLM_R_X5Y135_SLICE_X7Y135_D5Q;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A = CLBLM_R_X5Y136_SLICE_X6Y136_AO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B = CLBLM_R_X5Y136_SLICE_X6Y136_BO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C = CLBLM_R_X5Y136_SLICE_X6Y136_CO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D = CLBLM_R_X5Y136_SLICE_X6Y136_DO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_BMUX = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A = CLBLM_R_X5Y136_SLICE_X7Y136_AO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B = CLBLM_R_X5Y136_SLICE_X7Y136_BO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C = CLBLM_R_X5Y136_SLICE_X7Y136_CO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D = CLBLM_R_X5Y136_SLICE_X7Y136_DO6;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_CMUX = CLBLM_R_X5Y136_SLICE_X7Y136_C5Q;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_DMUX = CLBLM_R_X5Y136_SLICE_X7Y136_D5Q;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A = CLBLM_R_X5Y137_SLICE_X6Y137_AO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B = CLBLM_R_X5Y137_SLICE_X6Y137_BO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C = CLBLM_R_X5Y137_SLICE_X6Y137_CO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D = CLBLM_R_X5Y137_SLICE_X6Y137_DO6;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_DMUX = CLBLM_R_X5Y137_SLICE_X6Y137_DO5;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A = CLBLM_R_X5Y137_SLICE_X7Y137_AO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B = CLBLM_R_X5Y137_SLICE_X7Y137_BO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C = CLBLM_R_X5Y137_SLICE_X7Y137_CO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_AMUX = CLBLM_R_X5Y137_SLICE_X7Y137_A5Q;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_BMUX = CLBLM_R_X5Y137_SLICE_X7Y137_B5Q;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A = CLBLM_R_X5Y138_SLICE_X6Y138_AO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B = CLBLM_R_X5Y138_SLICE_X6Y138_BO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C = CLBLM_R_X5Y138_SLICE_X6Y138_CO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D = CLBLM_R_X5Y138_SLICE_X6Y138_DO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_BMUX = CLBLM_R_X5Y138_SLICE_X6Y138_B5Q;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_DMUX = CLBLM_R_X5Y138_SLICE_X6Y138_DO5;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A = CLBLM_R_X5Y138_SLICE_X7Y138_AO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B = CLBLM_R_X5Y138_SLICE_X7Y138_BO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C = CLBLM_R_X5Y138_SLICE_X7Y138_CO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D = CLBLM_R_X5Y138_SLICE_X7Y138_DO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_BMUX = CLBLM_R_X5Y138_SLICE_X7Y138_BO5;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A = CLBLM_R_X5Y139_SLICE_X6Y139_AO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B = CLBLM_R_X5Y139_SLICE_X6Y139_BO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C = CLBLM_R_X5Y139_SLICE_X6Y139_CO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D = CLBLM_R_X5Y139_SLICE_X6Y139_DO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_CMUX = CLBLM_R_X5Y139_SLICE_X6Y139_C5Q;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A = CLBLM_R_X5Y139_SLICE_X7Y139_AO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B = CLBLM_R_X5Y139_SLICE_X7Y139_BO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C = CLBLM_R_X5Y139_SLICE_X7Y139_CO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D = CLBLM_R_X5Y139_SLICE_X7Y139_DO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_AMUX = CLBLM_R_X5Y139_SLICE_X7Y139_A5Q;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_BMUX = CLBLM_R_X5Y139_SLICE_X7Y139_B5Q;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A = CLBLM_R_X5Y140_SLICE_X6Y140_AO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B = CLBLM_R_X5Y140_SLICE_X6Y140_BO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C = CLBLM_R_X5Y140_SLICE_X6Y140_CO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D = CLBLM_R_X5Y140_SLICE_X6Y140_DO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_AMUX = CLBLM_R_X5Y140_SLICE_X6Y140_A5Q;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_BMUX = CLBLM_R_X5Y140_SLICE_X6Y140_BO5;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A = CLBLM_R_X5Y140_SLICE_X7Y140_AO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B = CLBLM_R_X5Y140_SLICE_X7Y140_BO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C = CLBLM_R_X5Y140_SLICE_X7Y140_CO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D = CLBLM_R_X5Y140_SLICE_X7Y140_DO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_AMUX = CLBLM_R_X5Y140_SLICE_X7Y140_A5Q;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_BMUX = CLBLM_R_X5Y140_SLICE_X7Y140_B5Q;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A = CLBLM_R_X5Y141_SLICE_X6Y141_AO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B = CLBLM_R_X5Y141_SLICE_X6Y141_BO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C = CLBLM_R_X5Y141_SLICE_X6Y141_CO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D = CLBLM_R_X5Y141_SLICE_X6Y141_DO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A = CLBLM_R_X5Y141_SLICE_X7Y141_AO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B = CLBLM_R_X5Y141_SLICE_X7Y141_BO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C = CLBLM_R_X5Y141_SLICE_X7Y141_CO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D = CLBLM_R_X5Y141_SLICE_X7Y141_DO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_AMUX = CLBLM_R_X5Y141_SLICE_X7Y141_AO5;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A = CLBLM_R_X5Y142_SLICE_X6Y142_AO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B = CLBLM_R_X5Y142_SLICE_X6Y142_BO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C = CLBLM_R_X5Y142_SLICE_X6Y142_CO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D = CLBLM_R_X5Y142_SLICE_X6Y142_DO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_BMUX = CLBLM_R_X5Y142_SLICE_X6Y142_B5Q;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A = CLBLM_R_X5Y142_SLICE_X7Y142_AO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B = CLBLM_R_X5Y142_SLICE_X7Y142_BO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C = CLBLM_R_X5Y142_SLICE_X7Y142_CO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D = CLBLM_R_X5Y142_SLICE_X7Y142_DO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_BMUX = CLBLM_R_X5Y142_SLICE_X7Y142_BO5;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A = CLBLM_R_X5Y143_SLICE_X6Y143_AO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B = CLBLM_R_X5Y143_SLICE_X6Y143_BO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C = CLBLM_R_X5Y143_SLICE_X6Y143_CO6;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D = CLBLM_R_X5Y143_SLICE_X6Y143_DO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A = CLBLM_R_X5Y143_SLICE_X7Y143_AO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B = CLBLM_R_X5Y143_SLICE_X7Y143_BO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C = CLBLM_R_X5Y143_SLICE_X7Y143_CO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D = CLBLM_R_X5Y143_SLICE_X7Y143_DO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A = CLBLM_R_X7Y129_SLICE_X8Y129_AO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B = CLBLM_R_X7Y129_SLICE_X8Y129_BO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C = CLBLM_R_X7Y129_SLICE_X8Y129_CO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D = CLBLM_R_X7Y129_SLICE_X8Y129_DO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A = CLBLM_R_X7Y129_SLICE_X9Y129_AO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B = CLBLM_R_X7Y129_SLICE_X9Y129_BO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C = CLBLM_R_X7Y129_SLICE_X9Y129_CO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D = CLBLM_R_X7Y129_SLICE_X9Y129_DO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A = CLBLM_R_X7Y130_SLICE_X8Y130_AO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B = CLBLM_R_X7Y130_SLICE_X8Y130_BO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D = CLBLM_R_X7Y130_SLICE_X8Y130_DO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_CMUX = CLBLM_R_X7Y130_SLICE_X8Y130_CO5;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_DMUX = CLBLM_R_X7Y130_SLICE_X8Y130_DO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A = CLBLM_R_X7Y130_SLICE_X9Y130_AO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B = CLBLM_R_X7Y130_SLICE_X9Y130_BO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C = CLBLM_R_X7Y130_SLICE_X9Y130_CO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D = CLBLM_R_X7Y130_SLICE_X9Y130_DO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A = CLBLM_R_X7Y131_SLICE_X8Y131_AO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B = CLBLM_R_X7Y131_SLICE_X8Y131_BO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C = CLBLM_R_X7Y131_SLICE_X8Y131_CO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D = CLBLM_R_X7Y131_SLICE_X8Y131_DO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_AMUX = CLBLM_R_X7Y131_SLICE_X8Y131_A5Q;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_BMUX = CLBLM_R_X7Y131_SLICE_X8Y131_BO5;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_CMUX = CLBLM_R_X7Y131_SLICE_X8Y131_C5Q;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A = CLBLM_R_X7Y131_SLICE_X9Y131_AO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B = CLBLM_R_X7Y131_SLICE_X9Y131_BO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C = CLBLM_R_X7Y131_SLICE_X9Y131_CO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D = CLBLM_R_X7Y131_SLICE_X9Y131_DO6;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_DMUX = CLBLM_R_X7Y131_SLICE_X9Y131_D5Q;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A = CLBLM_R_X7Y132_SLICE_X8Y132_AO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B = CLBLM_R_X7Y132_SLICE_X8Y132_BO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C = CLBLM_R_X7Y132_SLICE_X8Y132_CO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D = CLBLM_R_X7Y132_SLICE_X8Y132_DO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_DMUX = CLBLM_R_X7Y132_SLICE_X8Y132_D5Q;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A = CLBLM_R_X7Y132_SLICE_X9Y132_AO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B = CLBLM_R_X7Y132_SLICE_X9Y132_BO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C = CLBLM_R_X7Y132_SLICE_X9Y132_CO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D = CLBLM_R_X7Y132_SLICE_X9Y132_DO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_AMUX = CLBLM_R_X7Y132_SLICE_X9Y132_A5Q;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_DMUX = CLBLM_R_X7Y132_SLICE_X9Y132_D5Q;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A = CLBLM_R_X7Y133_SLICE_X8Y133_AO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B = CLBLM_R_X7Y133_SLICE_X8Y133_BO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C = CLBLM_R_X7Y133_SLICE_X8Y133_CO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D = CLBLM_R_X7Y133_SLICE_X8Y133_DO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_AMUX = CLBLM_R_X7Y133_SLICE_X8Y133_A5Q;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_CMUX = CLBLM_R_X7Y133_SLICE_X8Y133_C5Q;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_DMUX = CLBLM_R_X7Y133_SLICE_X8Y133_D5Q;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A = CLBLM_R_X7Y133_SLICE_X9Y133_AO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B = CLBLM_R_X7Y133_SLICE_X9Y133_BO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C = CLBLM_R_X7Y133_SLICE_X9Y133_CO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D = CLBLM_R_X7Y133_SLICE_X9Y133_DO6;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_AMUX = CLBLM_R_X7Y133_SLICE_X9Y133_A5Q;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_BMUX = CLBLM_R_X7Y133_SLICE_X9Y133_B5Q;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_CMUX = CLBLM_R_X7Y133_SLICE_X9Y133_C5Q;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_DMUX = CLBLM_R_X7Y133_SLICE_X9Y133_D5Q;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A = CLBLM_R_X7Y134_SLICE_X8Y134_AO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B = CLBLM_R_X7Y134_SLICE_X8Y134_BO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C = CLBLM_R_X7Y134_SLICE_X8Y134_CO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D = CLBLM_R_X7Y134_SLICE_X8Y134_DO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_AMUX = CLBLM_R_X7Y134_SLICE_X8Y134_A5Q;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_BMUX = CLBLM_R_X7Y134_SLICE_X8Y134_B5Q;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_CMUX = CLBLM_R_X7Y134_SLICE_X8Y134_C5Q;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_DMUX = CLBLM_R_X7Y134_SLICE_X8Y134_DO5;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A = CLBLM_R_X7Y134_SLICE_X9Y134_AO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B = CLBLM_R_X7Y134_SLICE_X9Y134_BO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C = CLBLM_R_X7Y134_SLICE_X9Y134_CO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D = CLBLM_R_X7Y134_SLICE_X9Y134_DO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A = CLBLM_R_X7Y135_SLICE_X8Y135_AO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B = CLBLM_R_X7Y135_SLICE_X8Y135_BO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C = CLBLM_R_X7Y135_SLICE_X8Y135_CO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D = CLBLM_R_X7Y135_SLICE_X8Y135_DO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A = CLBLM_R_X7Y135_SLICE_X9Y135_AO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B = CLBLM_R_X7Y135_SLICE_X9Y135_BO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C = CLBLM_R_X7Y135_SLICE_X9Y135_CO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D = CLBLM_R_X7Y135_SLICE_X9Y135_DO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_AMUX = CLBLM_R_X7Y135_SLICE_X9Y135_A5Q;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_BMUX = CLBLM_R_X7Y135_SLICE_X9Y135_B5Q;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_CMUX = CLBLM_R_X7Y135_SLICE_X9Y135_C5Q;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_DMUX = CLBLM_R_X7Y135_SLICE_X9Y135_D5Q;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A = CLBLM_R_X7Y136_SLICE_X8Y136_AO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B = CLBLM_R_X7Y136_SLICE_X8Y136_BO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C = CLBLM_R_X7Y136_SLICE_X8Y136_CO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D = CLBLM_R_X7Y136_SLICE_X8Y136_DO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_AMUX = CLBLM_R_X7Y136_SLICE_X8Y136_A5Q;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_BMUX = CLBLM_R_X7Y136_SLICE_X8Y136_B5Q;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_CMUX = CLBLM_R_X7Y136_SLICE_X8Y136_C5Q;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_DMUX = CLBLM_R_X7Y136_SLICE_X8Y136_D5Q;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A = CLBLM_R_X7Y136_SLICE_X9Y136_AO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B = CLBLM_R_X7Y136_SLICE_X9Y136_BO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C = CLBLM_R_X7Y136_SLICE_X9Y136_CO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D = CLBLM_R_X7Y136_SLICE_X9Y136_DO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_AMUX = CLBLM_R_X7Y136_SLICE_X9Y136_A5Q;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_DMUX = CLBLM_R_X7Y136_SLICE_X9Y136_D5Q;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A = CLBLM_R_X7Y137_SLICE_X8Y137_AO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B = CLBLM_R_X7Y137_SLICE_X8Y137_BO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C = CLBLM_R_X7Y137_SLICE_X8Y137_CO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D = CLBLM_R_X7Y137_SLICE_X8Y137_DO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_BMUX = CLBLM_R_X7Y137_SLICE_X8Y137_B5Q;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_CMUX = CLBLM_R_X7Y137_SLICE_X8Y137_C5Q;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_DMUX = CLBLM_R_X7Y137_SLICE_X8Y137_D5Q;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A = CLBLM_R_X7Y137_SLICE_X9Y137_AO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B = CLBLM_R_X7Y137_SLICE_X9Y137_BO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C = CLBLM_R_X7Y137_SLICE_X9Y137_CO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D = CLBLM_R_X7Y137_SLICE_X9Y137_DO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_DMUX = CLBLM_R_X7Y137_SLICE_X9Y137_D5Q;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A = CLBLM_R_X7Y138_SLICE_X8Y138_AO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B = CLBLM_R_X7Y138_SLICE_X8Y138_BO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C = CLBLM_R_X7Y138_SLICE_X8Y138_CO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D = CLBLM_R_X7Y138_SLICE_X8Y138_DO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_BMUX = CLBLM_R_X7Y138_SLICE_X8Y138_B5Q;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_DMUX = CLBLM_R_X7Y138_SLICE_X8Y138_D5Q;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A = CLBLM_R_X7Y138_SLICE_X9Y138_AO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B = CLBLM_R_X7Y138_SLICE_X9Y138_BO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C = CLBLM_R_X7Y138_SLICE_X9Y138_CO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D = CLBLM_R_X7Y138_SLICE_X9Y138_DO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_AMUX = CLBLM_R_X7Y138_SLICE_X9Y138_A5Q;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_BMUX = CLBLM_R_X7Y138_SLICE_X9Y138_B5Q;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_CMUX = CLBLM_R_X7Y138_SLICE_X9Y138_C5Q;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A = CLBLM_R_X7Y139_SLICE_X8Y139_AO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B = CLBLM_R_X7Y139_SLICE_X8Y139_BO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C = CLBLM_R_X7Y139_SLICE_X8Y139_CO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D = CLBLM_R_X7Y139_SLICE_X8Y139_DO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_AMUX = CLBLM_R_X7Y139_SLICE_X8Y139_AO5;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A = CLBLM_R_X7Y139_SLICE_X9Y139_AO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B = CLBLM_R_X7Y139_SLICE_X9Y139_BO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C = CLBLM_R_X7Y139_SLICE_X9Y139_CO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A = CLBLM_R_X7Y140_SLICE_X8Y140_AO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B = CLBLM_R_X7Y140_SLICE_X8Y140_BO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C = CLBLM_R_X7Y140_SLICE_X8Y140_CO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D = CLBLM_R_X7Y140_SLICE_X8Y140_DO6;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_BMUX = CLBLM_R_X7Y140_SLICE_X8Y140_B5Q;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_CMUX = CLBLM_R_X7Y140_SLICE_X8Y140_C5Q;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_DMUX = CLBLM_R_X7Y140_SLICE_X8Y140_D5Q;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A = CLBLM_R_X7Y140_SLICE_X9Y140_AO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B = CLBLM_R_X7Y140_SLICE_X9Y140_BO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C = CLBLM_R_X7Y140_SLICE_X9Y140_CO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D = CLBLM_R_X7Y140_SLICE_X9Y140_DO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_DMUX = CLBLM_R_X7Y140_SLICE_X9Y140_D5Q;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A = CLBLM_R_X7Y141_SLICE_X8Y141_AO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B = CLBLM_R_X7Y141_SLICE_X8Y141_BO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C = CLBLM_R_X7Y141_SLICE_X8Y141_CO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_AMUX = CLBLM_R_X7Y141_SLICE_X8Y141_A5Q;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_BMUX = CLBLM_R_X7Y141_SLICE_X8Y141_BO5;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A = CLBLM_R_X7Y141_SLICE_X9Y141_AO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B = CLBLM_R_X7Y141_SLICE_X9Y141_BO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C = CLBLM_R_X7Y141_SLICE_X9Y141_CO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D = CLBLM_R_X7Y141_SLICE_X9Y141_DO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_AMUX = CLBLM_R_X7Y141_SLICE_X9Y141_A5Q;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A = CLBLM_R_X7Y142_SLICE_X8Y142_AO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B = CLBLM_R_X7Y142_SLICE_X8Y142_BO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C = CLBLM_R_X7Y142_SLICE_X8Y142_CO6;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D = CLBLM_R_X7Y142_SLICE_X8Y142_DO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A = CLBLM_R_X7Y142_SLICE_X9Y142_AO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B = CLBLM_R_X7Y142_SLICE_X9Y142_BO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C = CLBLM_R_X7Y142_SLICE_X9Y142_CO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_DMUX = CLBLM_R_X7Y142_SLICE_X9Y142_DO5;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A = CLBLM_R_X7Y143_SLICE_X8Y143_AO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B = CLBLM_R_X7Y143_SLICE_X8Y143_BO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C = CLBLM_R_X7Y143_SLICE_X8Y143_CO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D = CLBLM_R_X7Y143_SLICE_X8Y143_DO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_AMUX = CLBLM_R_X7Y143_SLICE_X8Y143_A5Q;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_BMUX = CLBLM_R_X7Y143_SLICE_X8Y143_BO5;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A = CLBLM_R_X7Y143_SLICE_X9Y143_AO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B = CLBLM_R_X7Y143_SLICE_X9Y143_BO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C = CLBLM_R_X7Y143_SLICE_X9Y143_CO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D = CLBLM_R_X7Y143_SLICE_X9Y143_DO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_BMUX = CLBLM_R_X7Y143_SLICE_X9Y143_BO5;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A = CLBLM_R_X11Y131_SLICE_X14Y131_AO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B = CLBLM_R_X11Y131_SLICE_X14Y131_BO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D = CLBLM_R_X11Y131_SLICE_X14Y131_DO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_AMUX = CLBLM_R_X11Y131_SLICE_X14Y131_AO5;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A = CLBLM_R_X11Y131_SLICE_X15Y131_AO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B = CLBLM_R_X11Y131_SLICE_X15Y131_BO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C = CLBLM_R_X11Y131_SLICE_X15Y131_CO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D = CLBLM_R_X11Y131_SLICE_X15Y131_DO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A = CLBLM_R_X11Y132_SLICE_X14Y132_AO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B = CLBLM_R_X11Y132_SLICE_X14Y132_BO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C = CLBLM_R_X11Y132_SLICE_X14Y132_CO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D = CLBLM_R_X11Y132_SLICE_X14Y132_DO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A = CLBLM_R_X11Y132_SLICE_X15Y132_AO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B = CLBLM_R_X11Y132_SLICE_X15Y132_BO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C = CLBLM_R_X11Y132_SLICE_X15Y132_CO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D = CLBLM_R_X11Y132_SLICE_X15Y132_DO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_AMUX = CLBLM_R_X11Y132_SLICE_X15Y132_AO5;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_BMUX = CLBLM_R_X11Y132_SLICE_X15Y132_BO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A = CLBLM_R_X11Y133_SLICE_X14Y133_AO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B = CLBLM_R_X11Y133_SLICE_X14Y133_BO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C = CLBLM_R_X11Y133_SLICE_X14Y133_CO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D = CLBLM_R_X11Y133_SLICE_X14Y133_DO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_CMUX = CLBLM_R_X11Y133_SLICE_X14Y133_CO5;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_DMUX = CLBLM_R_X11Y133_SLICE_X14Y133_DO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A = CLBLM_R_X11Y133_SLICE_X15Y133_AO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B = CLBLM_R_X11Y133_SLICE_X15Y133_BO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C = CLBLM_R_X11Y133_SLICE_X15Y133_CO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D = CLBLM_R_X11Y133_SLICE_X15Y133_DO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A = CLBLM_R_X11Y134_SLICE_X14Y134_AO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B = CLBLM_R_X11Y134_SLICE_X14Y134_BO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C = CLBLM_R_X11Y134_SLICE_X14Y134_CO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D = CLBLM_R_X11Y134_SLICE_X14Y134_DO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_AMUX = CLBLM_R_X11Y134_SLICE_X14Y134_AO5;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A = CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B = CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C = CLBLM_R_X11Y134_SLICE_X15Y134_CO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D = CLBLM_R_X11Y134_SLICE_X15Y134_DO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_BMUX = CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A = CLBLM_R_X11Y135_SLICE_X14Y135_AO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B = CLBLM_R_X11Y135_SLICE_X14Y135_BO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C = CLBLM_R_X11Y135_SLICE_X14Y135_CO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D = CLBLM_R_X11Y135_SLICE_X14Y135_DO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A = CLBLM_R_X11Y135_SLICE_X15Y135_AO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B = CLBLM_R_X11Y135_SLICE_X15Y135_BO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C = CLBLM_R_X11Y135_SLICE_X15Y135_CO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D = CLBLM_R_X11Y135_SLICE_X15Y135_DO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A = CLBLM_R_X11Y136_SLICE_X14Y136_AO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B = CLBLM_R_X11Y136_SLICE_X14Y136_BO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C = CLBLM_R_X11Y136_SLICE_X14Y136_CO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D = CLBLM_R_X11Y136_SLICE_X14Y136_DO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_DMUX = CLBLM_R_X11Y136_SLICE_X14Y136_DO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A = CLBLM_R_X11Y136_SLICE_X15Y136_AO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B = CLBLM_R_X11Y136_SLICE_X15Y136_BO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C = CLBLM_R_X11Y136_SLICE_X15Y136_CO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D = CLBLM_R_X11Y136_SLICE_X15Y136_DO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_AMUX = CLBLM_R_X11Y136_SLICE_X15Y136_AO5;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A = CLBLM_R_X11Y137_SLICE_X14Y137_AO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B = CLBLM_R_X11Y137_SLICE_X14Y137_BO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C = CLBLM_R_X11Y137_SLICE_X14Y137_CO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D = CLBLM_R_X11Y137_SLICE_X14Y137_DO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_AMUX = CLBLM_R_X11Y137_SLICE_X14Y137_AO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A = CLBLM_R_X11Y137_SLICE_X15Y137_AO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B = CLBLM_R_X11Y137_SLICE_X15Y137_BO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C = CLBLM_R_X11Y137_SLICE_X15Y137_CO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D = CLBLM_R_X11Y137_SLICE_X15Y137_DO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A = CLBLM_R_X11Y138_SLICE_X14Y138_AO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B = CLBLM_R_X11Y138_SLICE_X14Y138_BO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C = CLBLM_R_X11Y138_SLICE_X14Y138_CO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D = CLBLM_R_X11Y138_SLICE_X14Y138_DO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A = CLBLM_R_X11Y138_SLICE_X15Y138_AO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B = CLBLM_R_X11Y138_SLICE_X15Y138_BO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C = CLBLM_R_X11Y138_SLICE_X15Y138_CO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D = CLBLM_R_X11Y138_SLICE_X15Y138_DO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A = CLBLM_R_X11Y139_SLICE_X14Y139_AO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B = CLBLM_R_X11Y139_SLICE_X14Y139_BO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C = CLBLM_R_X11Y139_SLICE_X14Y139_CO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D = CLBLM_R_X11Y139_SLICE_X14Y139_DO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_AMUX = CLBLM_R_X11Y139_SLICE_X14Y139_AO5;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A = CLBLM_R_X11Y139_SLICE_X15Y139_AO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B = CLBLM_R_X11Y139_SLICE_X15Y139_BO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C = CLBLM_R_X11Y139_SLICE_X15Y139_CO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D = CLBLM_R_X11Y139_SLICE_X15Y139_DO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_AMUX = CLBLM_R_X11Y139_SLICE_X15Y139_AO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_DMUX = CLBLM_R_X11Y139_SLICE_X15Y139_DO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A = CLBLM_R_X11Y140_SLICE_X14Y140_AO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B = CLBLM_R_X11Y140_SLICE_X14Y140_BO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C = CLBLM_R_X11Y140_SLICE_X14Y140_CO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D = CLBLM_R_X11Y140_SLICE_X14Y140_DO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_AMUX = CLBLM_R_X11Y140_SLICE_X14Y140_AO5;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_BMUX = CLBLM_R_X11Y140_SLICE_X14Y140_BO5;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A = CLBLM_R_X11Y140_SLICE_X15Y140_AO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B = CLBLM_R_X11Y140_SLICE_X15Y140_BO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C = CLBLM_R_X11Y140_SLICE_X15Y140_CO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D = CLBLM_R_X11Y140_SLICE_X15Y140_DO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_BMUX = CLBLM_R_X11Y140_SLICE_X15Y140_B5Q;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_CMUX = CLBLM_R_X11Y140_SLICE_X15Y140_CO5;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A = CLBLM_R_X11Y141_SLICE_X14Y141_AO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B = CLBLM_R_X11Y141_SLICE_X14Y141_BO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C = CLBLM_R_X11Y141_SLICE_X14Y141_CO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D = CLBLM_R_X11Y141_SLICE_X14Y141_DO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A = CLBLM_R_X11Y141_SLICE_X15Y141_AO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B = CLBLM_R_X11Y141_SLICE_X15Y141_BO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C = CLBLM_R_X11Y141_SLICE_X15Y141_CO6;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D = CLBLM_R_X11Y141_SLICE_X15Y141_DO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A = CLBLM_R_X11Y142_SLICE_X14Y142_AO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B = CLBLM_R_X11Y142_SLICE_X14Y142_BO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C = CLBLM_R_X11Y142_SLICE_X14Y142_CO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D = CLBLM_R_X11Y142_SLICE_X14Y142_DO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A = CLBLM_R_X11Y142_SLICE_X15Y142_AO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B = CLBLM_R_X11Y142_SLICE_X15Y142_BO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C = CLBLM_R_X11Y142_SLICE_X15Y142_CO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D = CLBLM_R_X11Y142_SLICE_X15Y142_DO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_AMUX = CLBLM_R_X11Y142_SLICE_X15Y142_AO5;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_A = CLBLM_R_X13Y134_SLICE_X18Y134_AO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_B = CLBLM_R_X13Y134_SLICE_X18Y134_BO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_C = CLBLM_R_X13Y134_SLICE_X18Y134_CO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_D = CLBLM_R_X13Y134_SLICE_X18Y134_DO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_DMUX = CLBLM_R_X13Y134_SLICE_X18Y134_DO6;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_A = CLBLM_R_X13Y134_SLICE_X19Y134_AO6;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_B = CLBLM_R_X13Y134_SLICE_X19Y134_BO6;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_C = CLBLM_R_X13Y134_SLICE_X19Y134_CO6;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_D = CLBLM_R_X13Y134_SLICE_X19Y134_DO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_A = CLBLM_R_X13Y137_SLICE_X18Y137_AO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_B = CLBLM_R_X13Y137_SLICE_X18Y137_BO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_C = CLBLM_R_X13Y137_SLICE_X18Y137_CO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_D = CLBLM_R_X13Y137_SLICE_X18Y137_DO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_AMUX = CLBLM_R_X13Y137_SLICE_X18Y137_AO5;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_BMUX = CLBLM_R_X13Y137_SLICE_X18Y137_BO5;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_A = CLBLM_R_X13Y137_SLICE_X19Y137_AO6;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_B = CLBLM_R_X13Y137_SLICE_X19Y137_BO6;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_C = CLBLM_R_X13Y137_SLICE_X19Y137_CO6;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_D = CLBLM_R_X13Y137_SLICE_X19Y137_DO6;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_A = CLBLM_R_X13Y138_SLICE_X18Y138_AO6;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_B = CLBLM_R_X13Y138_SLICE_X18Y138_BO6;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_C = CLBLM_R_X13Y138_SLICE_X18Y138_CO6;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_D = CLBLM_R_X13Y138_SLICE_X18Y138_DO6;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_AMUX = CLBLM_R_X13Y138_SLICE_X18Y138_AO5;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_BMUX = CLBLM_R_X13Y138_SLICE_X18Y138_BO5;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_A = CLBLM_R_X13Y138_SLICE_X19Y138_AO6;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_B = CLBLM_R_X13Y138_SLICE_X19Y138_BO6;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_C = CLBLM_R_X13Y138_SLICE_X19Y138_CO6;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_D = CLBLM_R_X13Y138_SLICE_X19Y138_DO6;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A = CLBLM_R_X103Y178_SLICE_X162Y178_AO6;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B = CLBLM_R_X103Y178_SLICE_X162Y178_BO6;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C = CLBLM_R_X103Y178_SLICE_X162Y178_CO6;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D = CLBLM_R_X103Y178_SLICE_X162Y178_DO6;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B = CLBLM_R_X103Y178_SLICE_X163Y178_BO6;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C = CLBLM_R_X103Y178_SLICE_X163Y178_CO6;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D = CLBLM_R_X103Y178_SLICE_X163Y178_DO6;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_O = LIOB33_X0Y51_IOB_X0Y51_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_O = LIOB33_X0Y53_IOB_X0Y53_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_O = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y65_OLOGIC_X0Y66_OQ = CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  assign LIOI3_X0Y65_OLOGIC_X0Y66_TQ = 1'b1;
  assign LIOI3_X0Y65_OLOGIC_X0Y65_OQ = CLBLL_L_X2Y133_SLICE_X1Y133_BO6;
  assign LIOI3_X0Y65_OLOGIC_X0Y65_TQ = 1'b1;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_O = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_OQ = CLBLM_R_X5Y129_SLICE_X7Y129_BQ;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_OQ = CLBLM_R_X3Y136_SLICE_X2Y136_BQ;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_OQ = CLBLM_R_X5Y130_SLICE_X7Y130_D5Q;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_OQ = CLBLM_L_X10Y134_SLICE_X12Y134_B5Q;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_OQ = CLBLL_L_X4Y132_SLICE_X5Y132_BQ;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_OQ = CLBLL_L_X4Y137_SLICE_X5Y137_B5Q;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_OQ = CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_OQ = CLBLL_L_X4Y130_SLICE_X4Y130_BQ;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_OQ = CLBLL_L_X4Y132_SLICE_X5Y132_A5Q;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_OQ = CLBLL_L_X4Y131_SLICE_X4Y131_D5Q;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_OQ = CLBLM_L_X10Y131_SLICE_X12Y131_D5Q;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_OQ = CLBLM_R_X5Y138_SLICE_X6Y138_B5Q;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_OQ = CLBLM_R_X5Y130_SLICE_X7Y130_CQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_OQ = CLBLM_L_X10Y130_SLICE_X12Y130_B5Q;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = CLBLL_L_X4Y136_SLICE_X4Y136_CQ;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = CLBLM_R_X7Y135_SLICE_X9Y135_C5Q;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = CLBLM_R_X3Y132_SLICE_X3Y132_BQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_OQ = CLBLM_R_X5Y133_SLICE_X7Y133_AQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_OQ = CLBLM_L_X8Y138_SLICE_X10Y138_CQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_OQ = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_OQ = CLBLM_L_X10Y140_SLICE_X13Y140_D5Q;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_OQ = CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_OQ = CLBLM_R_X3Y132_SLICE_X3Y132_BQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_OQ = CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_OQ = CLBLL_L_X4Y133_SLICE_X4Y133_BO5;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = CLBLM_L_X8Y141_SLICE_X11Y141_BQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_OQ = CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = CLBLM_R_X3Y137_SLICE_X3Y137_D5Q;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = CLBLM_R_X3Y139_SLICE_X2Y139_C5Q;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_OQ = CLBLM_R_X3Y132_SLICE_X3Y132_BQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_OQ = CLBLL_L_X4Y134_SLICE_X5Y134_DQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_OQ = CLBLM_R_X3Y141_SLICE_X3Y141_BO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_OQ = CLBLM_R_X3Y137_SLICE_X2Y137_DO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_OQ = CLBLL_L_X4Y141_SLICE_X5Y141_DO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_OQ = CLBLL_L_X4Y139_SLICE_X5Y139_DO5;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_OQ = CLBLM_R_X5Y133_SLICE_X7Y133_A5Q;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_OQ = CLBLM_R_X3Y132_SLICE_X3Y132_BQ;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_OQ = CLBLM_L_X10Y137_SLICE_X13Y137_AQ;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_OQ = CLBLM_L_X10Y140_SLICE_X12Y140_AQ;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_OQ = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_OQ = CLBLM_L_X8Y135_SLICE_X11Y135_AQ;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_OQ = CLBLM_R_X3Y134_SLICE_X2Y134_AQ;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_OQ = CLBLM_R_X3Y132_SLICE_X3Y132_BQ;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_OQ = CLBLL_L_X4Y142_SLICE_X5Y142_CO5;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_OQ = CLBLM_R_X5Y140_SLICE_X6Y140_A5Q;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_OQ = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_OQ = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_OQ = RIOB33_X105Y101_IOB_X1Y101_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_OQ = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_OQ = RIOB33_X105Y119_IOB_X1Y120_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_OQ = RIOB33_X105Y119_IOB_X1Y119_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_OQ = RIOB33_X105Y121_IOB_X1Y122_I;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_OQ = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_OQ = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_OQ = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_OQ = RIOB33_X105Y125_IOB_X1Y125_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_OQ = RIOB33_X105Y123_IOB_X1Y124_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_OQ = RIOB33_X105Y127_IOB_X1Y127_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_OQ = RIOB33_X105Y125_IOB_X1Y126_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_OQ = RIOB33_X105Y131_IOB_X1Y132_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_OQ = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_OQ = RIOB33_X105Y119_IOB_X1Y120_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_OQ = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_OQ = CLBLM_R_X7Y143_SLICE_X8Y143_BO5;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_OQ = CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_OQ = CLBLM_R_X3Y141_SLICE_X2Y141_AO5;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_OQ = CLBLM_R_X3Y133_SLICE_X3Y133_CO6;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_OQ = CLBLL_L_X4Y143_SLICE_X4Y143_AO6;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_OQ = CLBLL_L_X4Y140_SLICE_X4Y140_DO6;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_OQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_OQ = CLBLM_R_X3Y141_SLICE_X2Y141_BO6;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_TQ = 1'b1;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ = CLBLM_R_X3Y136_SLICE_X2Y136_A5Q;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ = RIOB33_X105Y115_IOB_X1Y115_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ = 1'b1;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ = CLBLM_R_X3Y134_SLICE_X2Y134_AO5;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ = CLBLM_R_X5Y133_SLICE_X7Y133_CQ;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = CLBLM_R_X5Y138_SLICE_X7Y138_AQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = CLBLM_R_X3Y132_SLICE_X3Y132_BQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ = CLBLM_R_X3Y131_SLICE_X2Y131_AO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ = CLBLL_L_X2Y75_SLICE_X0Y75_AO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ = CLBLM_R_X7Y139_SLICE_X8Y139_AO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ = CLBLL_L_X4Y138_SLICE_X4Y138_AO5;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ = CLBLM_R_X3Y140_SLICE_X3Y140_AQ;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ = RIOB33_X105Y117_IOB_X1Y118_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ = RIOB33_X105Y129_IOB_X1Y129_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ = RIOB33_X105Y127_IOB_X1Y128_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ = RIOB33_X105Y103_IOB_X1Y103_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ = CLBLL_L_X4Y142_SLICE_X4Y142_BO6;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_OQ = CLBLL_L_X2Y134_SLICE_X1Y134_AO5;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ = CLBLM_R_X3Y141_SLICE_X2Y141_BQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ = CLBLL_L_X4Y130_SLICE_X4Y130_DQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = CLBLM_R_X3Y139_SLICE_X3Y139_A5Q;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = CLBLM_R_X7Y137_SLICE_X9Y137_D5Q;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ = RIOB33_X105Y101_IOB_X1Y102_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ = CLBLM_R_X5Y140_SLICE_X6Y140_BO5;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ = CLBLM_R_X3Y135_SLICE_X2Y135_AQ;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_O = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_O = RIOB33_X105Y123_IOB_X1Y124_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_O = RIOB33_X105Y135_IOB_X1Y136_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_O = RIOB33_X105Y135_IOB_X1Y135_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_O = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_O = RIOB33_X105Y139_IOB_X1Y139_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_O = RIOB33_X105Y141_IOB_X1Y142_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_O = RIOB33_X105Y141_IOB_X1Y141_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_O = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_O = RIOB33_X105Y145_IOB_X1Y145_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_O = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_O = RIOB33_X105Y147_IOB_X1Y147_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_OQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_TQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_OQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_OQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_OQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_OQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_OQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_OQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_OQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_OQ = CLBLM_R_X7Y140_SLICE_X9Y140_D5Q;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_OQ = CLBLM_R_X3Y141_SLICE_X3Y141_AO5;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_OQ = CLBLM_L_X10Y140_SLICE_X12Y140_AQ;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_OQ = CLBLM_R_X11Y142_SLICE_X15Y142_AO6;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_OQ = CLBLM_L_X8Y135_SLICE_X11Y135_AQ;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_OQ = CLBLM_L_X10Y137_SLICE_X13Y137_AQ;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_OQ = CLBLM_R_X3Y134_SLICE_X2Y134_AQ;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_OQ = CLBLM_R_X7Y141_SLICE_X9Y141_BO6;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_OQ = CLBLM_R_X5Y140_SLICE_X6Y140_BO5;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_OQ = CLBLM_R_X5Y140_SLICE_X6Y140_A5Q;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_OQ = CLBLM_R_X3Y138_SLICE_X3Y138_DO6;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_OQ = CLBLL_L_X4Y142_SLICE_X5Y142_CO5;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_OQ = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_OQ = CLBLM_L_X8Y140_SLICE_X11Y140_BQ;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_OQ = CLBLM_R_X3Y135_SLICE_X2Y135_AQ;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_OQ = CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_OQ = CLBLL_L_X4Y143_SLICE_X4Y143_AO6;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_OQ = 1'b0;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_OQ = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_OQ = CLBLM_R_X7Y141_SLICE_X8Y141_CO6;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_OQ = CLBLM_R_X11Y142_SLICE_X15Y142_AO5;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_OQ = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_OQ = CLBLM_L_X12Y142_SLICE_X16Y142_AO6;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_OQ = CLBLM_L_X12Y142_SLICE_X16Y142_BO5;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_OQ = CLBLM_L_X12Y142_SLICE_X16Y142_AO5;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_OQ = CLBLM_L_X12Y143_SLICE_X16Y143_AO6;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_OQ = CLBLM_L_X12Y143_SLICE_X16Y143_AO5;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_OQ = CLBLM_R_X11Y140_SLICE_X14Y140_AO5;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_TQ = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ = 1'b1;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_O = RIOB33_X105Y119_IOB_X1Y120_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O = RIOB33_X105Y119_IOB_X1Y119_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O = RIOB33_X105Y131_IOB_X1Y131_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O = RIOB33_X105Y143_IOB_X1Y144_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O = RIOB33_X105Y143_IOB_X1Y143_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ = CLBLM_R_X3Y140_SLICE_X3Y140_AQ;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ = CLBLL_L_X4Y141_SLICE_X5Y141_BO5;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ = CLBLM_R_X7Y143_SLICE_X8Y143_BO5;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ = CLBLM_L_X12Y142_SLICE_X16Y142_BO6;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ = CLBLM_R_X11Y142_SLICE_X14Y142_AO6;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O = RIOB33_X105Y137_IOB_X1Y137_I;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ = CLBLM_L_X10Y141_SLICE_X12Y141_BQ;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ = CLBLM_R_X7Y136_SLICE_X8Y136_D5Q;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ = CLBLL_L_X4Y141_SLICE_X5Y141_BO5;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_D1 = CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  assign LIOB33_X0Y147_IOB_X0Y148_O = CLBLL_L_X4Y141_SLICE_X5Y141_DO6;
  assign LIOB33_X0Y147_IOB_X0Y147_O = CLBLL_L_X4Y139_SLICE_X5Y139_DO5;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_D1 = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A1 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A3 = CLBLM_R_X7Y139_SLICE_X9Y139_AQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A4 = CLBLM_R_X11Y131_SLICE_X14Y131_BO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A5 = CLBLM_R_X7Y137_SLICE_X9Y137_AQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_A6 = CLBLM_R_X5Y139_SLICE_X7Y139_A5Q;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C4 = CLBLL_L_X4Y135_SLICE_X5Y135_CQ;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_T1 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C5 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B2 = CLBLM_R_X7Y139_SLICE_X9Y139_BQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B3 = CLBLM_R_X7Y137_SLICE_X9Y137_AQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B4 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B5 = CLBLM_L_X8Y140_SLICE_X10Y140_AQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_B6 = CLBLM_L_X12Y132_SLICE_X16Y132_AO6;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C6 = CLBLM_R_X7Y138_SLICE_X8Y138_D5Q;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_D1 = CLBLM_L_X8Y135_SLICE_X11Y135_AQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A1 = CLBLM_R_X5Y131_SLICE_X7Y131_CQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A2 = CLBLM_R_X5Y129_SLICE_X7Y129_BQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A3 = CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A5 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_A6 = CLBLM_R_X13Y134_SLICE_X18Y134_AO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C1 = CLBLM_R_X5Y138_SLICE_X6Y138_BQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C2 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C3 = CLBLM_R_X7Y134_SLICE_X8Y134_DO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B3 = CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B4 = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B5 = CLBLM_L_X8Y133_SLICE_X11Y133_BQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_B6 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D1 = CLBLM_R_X5Y140_SLICE_X6Y140_CQ;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C1 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C2 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C3 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C4 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C5 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_C6 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D4 = CLBLM_R_X5Y141_SLICE_X7Y141_CO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A1 = CLBLL_L_X4Y138_SLICE_X4Y138_CO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A2 = CLBLM_R_X7Y140_SLICE_X9Y140_DQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A3 = CLBLM_R_X5Y138_SLICE_X6Y138_BQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A4 = CLBLM_R_X7Y135_SLICE_X9Y135_DQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A5 = CLBLM_R_X7Y135_SLICE_X8Y135_AO6;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D1 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D2 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D3 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D4 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D5 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X7Y129_D6 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_A6 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_AX = CLBLM_L_X8Y137_SLICE_X10Y137_B5Q;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B1 = CLBLM_R_X5Y134_SLICE_X6Y134_DQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B2 = CLBLM_R_X5Y140_SLICE_X6Y140_CQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B3 = CLBLM_R_X3Y135_SLICE_X3Y135_DQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B4 = CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A1 = CLBLM_R_X5Y133_SLICE_X6Y133_B5Q;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A2 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A3 = CLBLM_R_X5Y129_SLICE_X6Y129_AQ;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A4 = CLBLM_R_X5Y130_SLICE_X6Y130_B5Q;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_A6 = CLBLM_R_X5Y130_SLICE_X6Y130_CO6;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C1 = CLBLM_R_X7Y138_SLICE_X9Y138_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C2 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C3 = CLBLL_L_X4Y139_SLICE_X4Y139_A5Q;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B1 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B2 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B3 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B4 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B5 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_B6 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A1 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A2 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A3 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A4 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A5 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_A6 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C1 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C2 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B1 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B2 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B3 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B4 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B5 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_B6 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C3 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C4 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C6 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C1 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C2 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C3 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C4 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C5 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_C6 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D1 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D2 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D3 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D4 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D5 = 1'b1;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_D6 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D1 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D2 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D3 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D4 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D5 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X0Y138_D6 = 1'b1;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D1 = CLBLM_L_X10Y137_SLICE_X12Y137_DO6;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A1 = CLBLM_R_X3Y137_SLICE_X3Y137_CQ;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A2 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A3 = CLBLM_R_X5Y138_SLICE_X6Y138_B5Q;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A4 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A5 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_A6 = 1'b1;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D4 = CLBLM_L_X10Y138_SLICE_X12Y138_DO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C1 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B1 = CLBLM_R_X3Y137_SLICE_X3Y137_CQ;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B2 = CLBLM_R_X3Y139_SLICE_X3Y139_BQ;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B3 = CLBLM_R_X5Y138_SLICE_X6Y138_B5Q;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B4 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B5 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_B6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C2 = 1'b1;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D6 = CLBLM_R_X11Y138_SLICE_X14Y138_BO6;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C1 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C2 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C3 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C4 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C5 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_C6 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C5 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C6 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D1 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D2 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D3 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D4 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D5 = 1'b1;
  assign CLBLL_L_X2Y138_SLICE_X1Y138_D6 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B3 = CLBLM_R_X3Y135_SLICE_X3Y135_BQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B4 = CLBLM_R_X5Y135_SLICE_X7Y135_BQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B5 = CLBLM_L_X8Y143_SLICE_X11Y143_AQ;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1 = 1'b1;
  assign LIOB33_X0Y151_IOB_X0Y152_O = CLBLM_R_X5Y133_SLICE_X7Y133_A5Q;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B6 = 1'b1;
  assign LIOB33_X0Y151_IOB_X0Y151_O = CLBLM_R_X3Y132_SLICE_X3Y132_BQ;
  assign RIOB33_SING_X105Y199_IOB_X1Y199_O = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1 = 1'b1;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_D = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_D = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D1 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D2 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D3 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C3 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D5 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C5 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D6 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C6 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A1 = CLBLM_R_X7Y135_SLICE_X9Y135_C5Q;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A2 = CLBLM_R_X7Y138_SLICE_X8Y138_D5Q;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A3 = CLBLM_R_X7Y140_SLICE_X9Y140_AQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A4 = CLBLM_L_X8Y138_SLICE_X11Y138_C5Q;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A5 = CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A5 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B2 = CLBLM_R_X7Y140_SLICE_X9Y140_BQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B3 = CLBLM_R_X7Y140_SLICE_X9Y140_AQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B4 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_B6 = CLBLM_R_X7Y134_SLICE_X8Y134_C5Q;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A1 = CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A2 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A3 = CLBLM_R_X5Y130_SLICE_X7Y130_AQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A4 = CLBLL_L_X4Y130_SLICE_X5Y130_A5Q;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_A6 = CLBLM_R_X7Y135_SLICE_X9Y135_C5Q;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C2 = CLBLM_R_X7Y140_SLICE_X9Y140_CQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_C3 = CLBLM_L_X10Y131_SLICE_X12Y131_D5Q;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B1 = CLBLL_L_X4Y134_SLICE_X4Y134_CQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B2 = CLBLM_R_X5Y130_SLICE_X7Y130_BQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B4 = CLBLL_L_X4Y134_SLICE_X4Y134_A5Q;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B5 = CLBLM_R_X5Y130_SLICE_X6Y130_B5Q;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_B6 = CLBLM_R_X7Y131_SLICE_X8Y131_A5Q;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D1 = CLBLM_R_X7Y133_SLICE_X9Y133_AQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C2 = CLBLM_R_X5Y130_SLICE_X7Y130_CQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C3 = CLBLM_R_X5Y139_SLICE_X7Y139_B5Q;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C4 = CLBLM_L_X8Y135_SLICE_X10Y135_CQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_C6 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D3 = CLBLM_L_X10Y141_SLICE_X13Y141_CQ;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D4 = CLBLM_R_X7Y136_SLICE_X8Y136_D5Q;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A1 = CLBLM_L_X8Y138_SLICE_X10Y138_CQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A2 = CLBLL_L_X4Y136_SLICE_X4Y136_D5Q;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A3 = CLBLM_R_X7Y140_SLICE_X8Y140_AQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A4 = CLBLM_R_X5Y135_SLICE_X7Y135_D5Q;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D1 = CLBLM_L_X10Y135_SLICE_X13Y135_AQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D2 = CLBLM_R_X7Y131_SLICE_X8Y131_C5Q;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D3 = CLBLL_L_X4Y136_SLICE_X4Y136_AQ;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D4 = CLBLM_R_X5Y133_SLICE_X7Y133_A5Q;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y130_SLICE_X7Y130_D6 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B4 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_A6 = CLBLM_R_X7Y141_SLICE_X9Y141_A5Q;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B5 = CLBLL_L_X4Y139_SLICE_X5Y139_C5Q;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_B2 = CLBLM_L_X8Y140_SLICE_X10Y140_D5Q;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A1 = CLBLL_L_X4Y130_SLICE_X5Y130_DO6;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A2 = CLBLM_R_X3Y131_SLICE_X3Y131_AQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A3 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A4 = CLBLM_R_X7Y131_SLICE_X8Y131_A5Q;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_A6 = CLBLM_R_X5Y131_SLICE_X6Y131_CO5;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B6 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C1 = CLBLM_R_X7Y133_SLICE_X8Y133_D5Q;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_C2 = CLBLM_R_X3Y139_SLICE_X2Y139_CQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B2 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B3 = CLBLL_L_X4Y130_SLICE_X4Y130_BQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B4 = CLBLM_R_X5Y133_SLICE_X6Y133_AQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B5 = CLBLM_L_X8Y132_SLICE_X10Y132_B5Q;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_B6 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D1 = CLBLL_L_X4Y140_SLICE_X5Y140_BQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D2 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C1 = CLBLM_R_X3Y131_SLICE_X3Y131_AQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C2 = CLBLM_R_X7Y131_SLICE_X8Y131_A5Q;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C3 = CLBLL_L_X4Y134_SLICE_X4Y134_CQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C4 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C5 = CLBLL_L_X4Y130_SLICE_X5Y130_AQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_C6 = CLBLM_R_X5Y130_SLICE_X7Y130_BQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D4 = CLBLM_R_X11Y141_SLICE_X14Y141_AQ;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D5 = CLBLL_L_X4Y136_SLICE_X5Y136_AQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y140_SLICE_X8Y140_D6 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_T1 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D1 = CLBLL_L_X4Y130_SLICE_X4Y130_BQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D2 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D3 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D4 = CLBLL_L_X4Y130_SLICE_X5Y130_B5Q;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D5 = 1'b1;
  assign CLBLM_R_X5Y130_SLICE_X6Y130_D6 = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C3 = CLBLM_R_X5Y142_SLICE_X7Y142_BO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C5 = CLBLM_R_X5Y141_SLICE_X7Y141_AO6;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C6 = CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  assign LIOB33_X0Y153_IOB_X0Y154_O = CLBLM_L_X10Y137_SLICE_X13Y137_AQ;
  assign LIOB33_X0Y153_IOB_X0Y153_O = CLBLM_L_X10Y140_SLICE_X12Y140_AQ;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_D1 = CLBLM_R_X11Y142_SLICE_X15Y142_AO6;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A1 = CLBLM_L_X10Y130_SLICE_X12Y130_B5Q;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A2 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A3 = CLBLM_L_X10Y133_SLICE_X12Y133_BQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A5 = CLBLM_R_X7Y135_SLICE_X9Y135_C5Q;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_A6 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B2 = CLBLM_R_X7Y134_SLICE_X8Y134_C5Q;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B3 = CLBLM_R_X3Y135_SLICE_X2Y135_AQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B4 = CLBLM_R_X7Y140_SLICE_X9Y140_BQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B5 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_B6 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A1 = CLBLL_L_X4Y135_SLICE_X4Y135_D5Q;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A2 = CLBLM_R_X5Y131_SLICE_X7Y131_DQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A3 = CLBLM_R_X5Y131_SLICE_X7Y131_AQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A5 = CLBLM_R_X5Y133_SLICE_X7Y133_AQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_A6 = CLBLL_L_X4Y133_SLICE_X5Y133_B5Q;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C1 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C2 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C3 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B1 = CLBLM_R_X5Y136_SLICE_X7Y136_DQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B2 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B4 = CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B5 = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_B6 = CLBLM_R_X5Y133_SLICE_X6Y133_A5Q;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D1 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C2 = CLBLM_R_X5Y131_SLICE_X7Y131_CQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C3 = CLBLL_L_X4Y135_SLICE_X5Y135_CQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C4 = CLBLL_L_X4Y140_SLICE_X5Y140_CQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C5 = CLBLM_R_X7Y138_SLICE_X9Y138_B5Q;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_C6 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D3 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D4 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A1 = CLBLM_R_X7Y135_SLICE_X9Y135_C5Q;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A4 = CLBLM_R_X5Y142_SLICE_X6Y142_CQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A5 = CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A6 = CLBLM_R_X5Y139_SLICE_X6Y139_CQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D2 = CLBLM_R_X5Y132_SLICE_X6Y132_AQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D3 = CLBLM_R_X5Y131_SLICE_X7Y131_DQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D4 = CLBLL_L_X4Y134_SLICE_X4Y134_DQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D5 = CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  assign CLBLM_R_X5Y131_SLICE_X7Y131_D6 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A5 = CLBLM_R_X7Y130_SLICE_X8Y130_CO5;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A6 = CLBLM_R_X5Y133_SLICE_X6Y133_A5Q;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_AX = CLBLM_R_X7Y142_SLICE_X9Y142_DO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B2 = CLBLL_L_X4Y140_SLICE_X5Y140_BQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B3 = CLBLM_R_X7Y140_SLICE_X9Y140_BQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A1 = CLBLM_R_X3Y131_SLICE_X3Y131_B5Q;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A2 = CLBLM_R_X11Y131_SLICE_X14Y131_BO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A3 = CLBLM_R_X5Y131_SLICE_X6Y131_AQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A4 = CLBLL_L_X4Y131_SLICE_X4Y131_AQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_A6 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C1 = CLBLL_L_X2Y138_SLICE_X1Y138_BO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C3 = CLBLL_L_X4Y140_SLICE_X5Y140_BQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B1 = CLBLM_R_X5Y131_SLICE_X6Y131_DO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B2 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B4 = CLBLM_L_X8Y135_SLICE_X10Y135_CQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B5 = CLBLM_R_X5Y129_SLICE_X6Y129_AQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_B6 = CLBLL_L_X4Y131_SLICE_X4Y131_AQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D1 = CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C1 = CLBLM_R_X7Y134_SLICE_X8Y134_AQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C2 = CLBLM_R_X5Y130_SLICE_X7Y130_BQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C3 = CLBLM_R_X7Y131_SLICE_X8Y131_A5Q;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C4 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C5 = CLBLM_L_X8Y132_SLICE_X10Y132_B5Q;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_C6 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B1 = CLBLM_R_X7Y132_SLICE_X8Y132_DQ;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D6 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D1 = CLBLL_L_X4Y130_SLICE_X5Y130_AQ;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D2 = CLBLL_L_X4Y134_SLICE_X4Y134_A5Q;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D3 = CLBLL_L_X4Y131_SLICE_X5Y131_CO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D4 = CLBLM_R_X5Y131_SLICE_X6Y131_CO6;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D5 = 1'b1;
  assign CLBLM_R_X5Y131_SLICE_X6Y131_D6 = CLBLL_L_X4Y131_SLICE_X5Y131_DO6;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_D1 = CLBLM_R_X3Y134_SLICE_X2Y134_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B6 = CLBLM_R_X5Y133_SLICE_X6Y133_A5Q;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_T1 = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_D1 = CLBLM_R_X3Y132_SLICE_X3Y132_BQ;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_T1 = 1'b1;
  assign LIOB33_X0Y155_IOB_X0Y156_O = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign LIOB33_X0Y155_IOB_X0Y155_O = CLBLM_L_X8Y135_SLICE_X11Y135_AQ;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1 = CLBLM_L_X12Y142_SLICE_X16Y142_BO6;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1 = CLBLM_R_X11Y142_SLICE_X14Y142_AO6;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_C4 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_C5 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_C6 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A1 = CLBLM_L_X8Y142_SLICE_X10Y142_CO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A2 = CLBLM_R_X7Y142_SLICE_X9Y142_BQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A3 = CLBLM_R_X7Y142_SLICE_X9Y142_AQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A4 = CLBLL_L_X4Y133_SLICE_X4Y133_BQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_A6 = CLBLM_R_X5Y140_SLICE_X7Y140_A5Q;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B1 = CLBLL_L_X4Y138_SLICE_X5Y138_DQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B2 = CLBLM_R_X7Y142_SLICE_X9Y142_BQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B4 = CLBLM_L_X8Y142_SLICE_X10Y142_CO6;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B5 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_B6 = CLBLM_R_X5Y140_SLICE_X7Y140_A5Q;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A2 = CLBLL_L_X4Y135_SLICE_X4Y135_D5Q;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A3 = CLBLM_R_X5Y132_SLICE_X7Y132_AQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A4 = CLBLM_R_X5Y134_SLICE_X7Y134_DQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A5 = CLBLM_L_X8Y131_SLICE_X11Y131_C5Q;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_A6 = CLBLM_R_X5Y133_SLICE_X7Y133_AQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C1 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C2 = CLBLM_R_X7Y142_SLICE_X9Y142_CQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C3 = CLBLM_L_X8Y141_SLICE_X11Y141_AQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B1 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B2 = CLBLM_R_X5Y132_SLICE_X7Y132_BQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B3 = CLBLM_L_X8Y140_SLICE_X11Y140_BQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B4 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_B6 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C2 = CLBLM_R_X5Y136_SLICE_X7Y136_DQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C3 = CLBLL_L_X4Y132_SLICE_X5Y132_A5Q;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C4 = CLBLL_L_X4Y134_SLICE_X4Y134_DQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C5 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_C6 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D3 = CLBLM_R_X7Y142_SLICE_X9Y142_BQ;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D4 = CLBLM_R_X7Y142_SLICE_X9Y142_AQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A1 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A2 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A3 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A4 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_D5 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D1 = CLBLM_R_X5Y134_SLICE_X6Y134_B5Q;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D2 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D3 = CLBLM_R_X5Y133_SLICE_X7Y133_CQ;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D4 = CLBLM_R_X7Y133_SLICE_X9Y133_DQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_D6 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D5 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X7Y132_D6 = CLBLL_L_X4Y131_SLICE_X4Y131_D5Q;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A6 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B1 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B2 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B3 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A1 = CLBLM_R_X5Y133_SLICE_X6Y133_DO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A2 = CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A3 = CLBLM_R_X5Y132_SLICE_X7Y132_C5Q;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A4 = CLBLM_R_X5Y132_SLICE_X6Y132_AQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_A6 = CLBLM_R_X5Y130_SLICE_X7Y130_DQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C1 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C2 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B1 = CLBLM_R_X5Y133_SLICE_X6Y133_DO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B2 = CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B3 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B4 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_B6 = CLBLM_R_X5Y130_SLICE_X7Y130_DQ;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D1 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D2 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D3 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C1 = CLBLL_L_X4Y130_SLICE_X4Y130_DQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C2 = CLBLL_L_X4Y132_SLICE_X5Y132_A5Q;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C3 = CLBLM_R_X5Y132_SLICE_X7Y132_DO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C4 = CLBLM_R_X5Y132_SLICE_X7Y132_CQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C5 = CLBLM_R_X5Y132_SLICE_X6Y132_DO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_C6 = CLBLL_L_X4Y133_SLICE_X4Y133_D5Q;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D4 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D5 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_D6 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D1 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D2 = CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D3 = CLBLM_R_X5Y130_SLICE_X6Y130_DO6;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D4 = CLBLL_L_X4Y130_SLICE_X4Y130_B5Q;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D5 = 1'b1;
  assign CLBLM_R_X5Y132_SLICE_X6Y132_D6 = CLBLM_R_X11Y140_SLICE_X15Y140_BQ;
  assign LIOB33_X0Y157_IOB_X0Y158_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOB33_X0Y157_IOB_X0Y157_O = CLBLM_R_X3Y140_SLICE_X3Y140_AQ;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_B5 = CLBLM_R_X11Y140_SLICE_X14Y140_AQ;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_B6 = RIOB33_X105Y139_IOB_X1Y140_I;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_C4 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_C5 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_C6 = 1'b1;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_D = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A1 = CLBLM_L_X8Y143_SLICE_X10Y143_CO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A2 = CLBLM_L_X8Y132_SLICE_X10Y132_BQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A3 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A4 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_A6 = CLBLM_R_X7Y143_SLICE_X9Y143_CO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B1 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B2 = CLBLM_R_X7Y133_SLICE_X8Y133_A5Q;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B3 = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B4 = CLBLM_L_X8Y141_SLICE_X11Y141_BQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B5 = CLBLM_L_X8Y143_SLICE_X10Y143_BO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_B6 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A1 = CLBLM_R_X5Y135_SLICE_X6Y135_A5Q;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A2 = CLBLM_R_X5Y134_SLICE_X7Y134_CQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A4 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A5 = CLBLM_L_X10Y131_SLICE_X12Y131_D5Q;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_A6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C1 = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C2 = CLBLM_R_X7Y133_SLICE_X8Y133_A5Q;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C3 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B1 = CLBLM_R_X7Y133_SLICE_X8Y133_CQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B2 = CLBLL_L_X4Y131_SLICE_X4Y131_D5Q;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B3 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B4 = CLBLM_L_X10Y140_SLICE_X13Y140_BQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_B6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D1 = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C2 = CLBLM_R_X3Y134_SLICE_X3Y134_A5Q;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C3 = CLBLM_R_X7Y134_SLICE_X8Y134_C5Q;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C4 = CLBLM_R_X5Y135_SLICE_X6Y135_A5Q;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C5 = CLBLM_R_X5Y133_SLICE_X7Y133_B5Q;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_C6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D3 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D4 = CLBLM_L_X8Y143_SLICE_X10Y143_BO5;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A1 = CLBLM_R_X7Y138_SLICE_X8Y138_B5Q;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A2 = CLBLM_R_X7Y143_SLICE_X9Y143_BO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A3 = CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A5 = CLBLM_R_X7Y143_SLICE_X8Y143_A5Q;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D2 = CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D3 = CLBLM_R_X3Y135_SLICE_X3Y135_BQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D4 = CLBLL_L_X4Y132_SLICE_X4Y132_AQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D5 = CLBLL_L_X4Y138_SLICE_X5Y138_DQ;
  assign CLBLM_R_X5Y133_SLICE_X7Y133_D6 = CLBLM_R_X3Y135_SLICE_X3Y135_CQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B4 = CLBLL_L_X4Y141_SLICE_X4Y141_AQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B5 = CLBLM_R_X7Y143_SLICE_X8Y143_A5Q;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_AX = CLBLM_R_X7Y143_SLICE_X8Y143_BO6;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B1 = CLBLM_R_X7Y143_SLICE_X9Y143_BO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A1 = CLBLM_R_X7Y133_SLICE_X9Y133_A5Q;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A2 = CLBLM_R_X5Y134_SLICE_X7Y134_D5Q;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A3 = CLBLM_R_X5Y137_SLICE_X6Y137_CQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A4 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_A6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C1 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C2 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C3 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B1 = CLBLM_R_X7Y135_SLICE_X8Y135_AQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B2 = CLBLM_R_X7Y139_SLICE_X9Y139_BQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B4 = CLBLL_L_X4Y133_SLICE_X5Y133_B5Q;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B5 = CLBLL_L_X4Y132_SLICE_X5Y132_CQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_B6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D1 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D2 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C1 = CLBLM_R_X7Y132_SLICE_X9Y132_DQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C2 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C4 = CLBLM_R_X5Y134_SLICE_X6Y134_C5Q;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C5 = CLBLM_R_X11Y134_SLICE_X14Y134_AO6;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_C6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D3 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D4 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D5 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_D6 = 1'b1;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D1 = CLBLL_L_X4Y137_SLICE_X5Y137_C5Q;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D2 = CLBLM_R_X5Y134_SLICE_X6Y134_CQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D3 = CLBLL_L_X4Y138_SLICE_X5Y138_DQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D4 = CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D5 = CLBLM_R_X3Y135_SLICE_X3Y135_BQ;
  assign CLBLM_R_X5Y133_SLICE_X6Y133_D6 = CLBLM_R_X3Y135_SLICE_X3Y135_CQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C4 = CLBLM_R_X11Y137_SLICE_X14Y137_AO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C5 = CLBLM_L_X12Y134_SLICE_X17Y134_DO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C6 = CLBLM_R_X11Y139_SLICE_X15Y139_DO6;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_D1 = CLBLL_L_X4Y142_SLICE_X5Y142_CO5;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D5 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_T1 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D6 = CLBLM_L_X8Y139_SLICE_X10Y139_CO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_D1 = CLBLM_R_X5Y129_SLICE_X7Y129_BQ;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_D1 = CLBLM_R_X5Y140_SLICE_X6Y140_A5Q;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_T1 = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_T1 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_D1 = CLBLM_R_X3Y136_SLICE_X2Y136_BQ;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_D1 = CLBLL_L_X2Y134_SLICE_X1Y134_AO5;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_OLOGIC_X0Y64_T1 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C4 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C5 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A1 = CLBLM_R_X5Y134_SLICE_X6Y134_DQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A2 = CLBLM_L_X10Y140_SLICE_X13Y140_BQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A3 = CLBLL_L_X4Y131_SLICE_X5Y131_AQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A5 = CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_A6 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_C6 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B1 = CLBLL_L_X4Y134_SLICE_X5Y134_CQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B2 = CLBLM_R_X5Y134_SLICE_X7Y134_BQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B3 = CLBLL_L_X4Y139_SLICE_X5Y139_CQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B4 = CLBLM_L_X8Y133_SLICE_X10Y133_C5Q;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_B6 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C1 = CLBLL_L_X4Y132_SLICE_X5Y132_C5Q;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C2 = CLBLM_L_X8Y134_SLICE_X10Y134_BO6;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C3 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C4 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C5 = CLBLM_L_X8Y139_SLICE_X11Y139_BQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B5 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B6 = CLBLM_R_X7Y140_SLICE_X8Y140_DQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y161_IOB_X0Y162_O = CLBLL_L_X4Y142_SLICE_X5Y142_CO5;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D2 = CLBLM_R_X7Y141_SLICE_X8Y141_A5Q;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D3 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D4 = CLBLM_L_X10Y133_SLICE_X13Y133_AQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D5 = CLBLM_R_X5Y134_SLICE_X6Y134_DQ;
  assign CLBLM_R_X5Y134_SLICE_X7Y134_D6 = 1'b1;
  assign LIOB33_X0Y161_IOB_X0Y161_O = CLBLM_R_X5Y140_SLICE_X6Y140_A5Q;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A1 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A2 = CLBLM_L_X10Y132_SLICE_X12Y132_AQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A3 = CLBLM_R_X11Y142_SLICE_X14Y142_AQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A5 = CLBLL_L_X4Y135_SLICE_X4Y135_C5Q;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_A6 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C1 = CLBLM_L_X12Y133_SLICE_X17Y133_AO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B1 = CLBLM_R_X7Y142_SLICE_X9Y142_CQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B2 = CLBLL_L_X4Y131_SLICE_X4Y131_D5Q;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B4 = CLBLM_R_X5Y133_SLICE_X6Y133_B5Q;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B5 = CLBLM_R_X7Y137_SLICE_X8Y137_AQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_B6 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D2 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C2 = CLBLM_R_X11Y138_SLICE_X14Y138_CO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C3 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C1 = CLBLM_R_X5Y134_SLICE_X6Y134_CQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C2 = CLBLM_R_X5Y130_SLICE_X7Y130_DQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C3 = 1'b1;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C4 = CLBLL_L_X4Y133_SLICE_X4Y133_A5Q;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C5 = CLBLM_R_X5Y137_SLICE_X6Y137_DO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D5 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C4 = CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C5 = CLBLM_R_X11Y139_SLICE_X14Y139_DO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y141_SLICE_X9Y141_D6 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_C6 = CLBLM_L_X10Y139_SLICE_X13Y139_DO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_CX = CLBLM_R_X5Y133_SLICE_X6Y133_CO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D2 = CLBLM_R_X5Y130_SLICE_X7Y130_DQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D3 = CLBLM_R_X5Y134_SLICE_X6Y134_DQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D4 = CLBLM_R_X5Y135_SLICE_X6Y135_CO6;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D5 = CLBLM_R_X5Y132_SLICE_X6Y132_AQ;
  assign CLBLM_R_X5Y134_SLICE_X6Y134_D6 = CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_D = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_D = RIOB33_X105Y145_IOB_X1Y145_I;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_A3 = CLBLM_R_X7Y141_SLICE_X8Y141_AQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D1 = CLBLM_L_X12Y135_SLICE_X17Y135_BO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D2 = CLBLM_L_X12Y139_SLICE_X16Y139_DO6;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D3 = CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D4 = CLBLL_L_X4Y130_SLICE_X5Y130_DO5;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D5 = CLBLM_L_X8Y139_SLICE_X10Y139_BO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_D6 = CLBLM_R_X3Y139_SLICE_X3Y139_BO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C3 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C4 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C5 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C6 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A6 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B4 = CLBLM_R_X7Y134_SLICE_X8Y134_C5Q;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B5 = CLBLL_L_X2Y138_SLICE_X1Y138_BO6;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_B6 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B1 = CLBLM_R_X13Y134_SLICE_X18Y134_AO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D2 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C4 = CLBLM_R_X7Y134_SLICE_X8Y134_C5Q;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D5 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D6 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_C6 = CLBLM_R_X7Y140_SLICE_X9Y140_BQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C2 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C3 = CLBLM_R_X7Y137_SLICE_X8Y137_CQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C4 = CLBLL_L_X4Y136_SLICE_X5Y136_D5Q;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C6 = CLBLM_L_X8Y134_SLICE_X10Y134_A5Q;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A1 = CLBLM_R_X5Y131_SLICE_X7Y131_AQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A3 = CLBLM_R_X5Y135_SLICE_X7Y135_AQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A4 = CLBLM_R_X11Y131_SLICE_X14Y131_BO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A5 = CLBLM_R_X5Y135_SLICE_X6Y135_AQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_A6 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOB33_X0Y163_IOB_X0Y163_O = CLBLM_R_X5Y140_SLICE_X6Y140_BO5;
  assign LIOB33_X0Y163_IOB_X0Y164_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B1 = CLBLM_R_X3Y137_SLICE_X3Y137_A5Q;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B2 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B3 = CLBLL_L_X4Y131_SLICE_X5Y131_B5Q;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B5 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_B6 = 1'b1;
  assign CLBLM_R_X7Y141_SLICE_X8Y141_D5 = CLBLM_R_X7Y141_SLICE_X8Y141_BO5;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C1 = CLBLM_R_X5Y139_SLICE_X7Y139_B5Q;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C2 = CLBLM_L_X8Y135_SLICE_X10Y135_AQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C3 = CLBLL_L_X4Y136_SLICE_X4Y136_AQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C4 = CLBLL_L_X4Y136_SLICE_X4Y136_CQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C5 = CLBLM_R_X11Y140_SLICE_X15Y140_CO6;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D1 = CLBLM_R_X5Y139_SLICE_X7Y139_AQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D2 = CLBLL_L_X4Y137_SLICE_X5Y137_C5Q;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D3 = CLBLL_L_X4Y132_SLICE_X5Y132_D5Q;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D4 = CLBLM_R_X7Y132_SLICE_X8Y132_CQ;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y135_SLICE_X7Y135_D6 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A1 = CLBLL_L_X4Y135_SLICE_X4Y135_CQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A3 = CLBLM_R_X7Y137_SLICE_X9Y137_D5Q;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A4 = CLBLM_R_X5Y135_SLICE_X7Y135_BQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A5 = CLBLM_R_X3Y135_SLICE_X3Y135_CQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_A6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B5 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B1 = CLBLL_L_X4Y134_SLICE_X5Y134_AQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B3 = CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B4 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B5 = CLBLM_L_X8Y135_SLICE_X10Y135_DQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_B6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B6 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C1 = CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C2 = CLBLM_R_X3Y135_SLICE_X3Y135_BQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C3 = CLBLM_R_X5Y134_SLICE_X6Y134_CQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C4 = CLBLM_R_X3Y135_SLICE_X3Y135_CQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C5 = CLBLM_R_X5Y135_SLICE_X6Y135_DO6;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_C6 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D1 = CLBLL_L_X4Y137_SLICE_X5Y137_C5Q;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D2 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D3 = CLBLL_L_X4Y138_SLICE_X5Y138_DQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D4 = CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D5 = 1'b1;
  assign CLBLM_R_X5Y135_SLICE_X6Y135_D6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C4 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C5 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D5 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1 = CLBLM_L_X10Y141_SLICE_X12Y141_BQ;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_D1 = 1'b0;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1 = 1'b1;
  assign LIOB33_X0Y165_IOB_X0Y166_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOB33_X0Y165_IOB_X0Y165_O = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A2 = CLBLM_R_X7Y133_SLICE_X8Y133_CQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A3 = CLBLM_R_X5Y136_SLICE_X7Y136_AQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A4 = CLBLL_L_X4Y135_SLICE_X4Y135_D5Q;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A5 = CLBLM_R_X5Y133_SLICE_X7Y133_AQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_A6 = CLBLL_L_X4Y142_SLICE_X4Y142_A5Q;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_D1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B1 = CLBLM_R_X7Y136_SLICE_X8Y136_CQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B2 = CLBLM_R_X5Y136_SLICE_X7Y136_BQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B4 = CLBLM_R_X7Y135_SLICE_X9Y135_C5Q;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B5 = CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_B6 = CLBLM_R_X11Y136_SLICE_X15Y136_AQ;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_T1 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_D1 = CLBLM_R_X5Y130_SLICE_X7Y130_D5Q;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C2 = CLBLM_R_X7Y136_SLICE_X9Y136_CQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C3 = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C4 = CLBLM_R_X5Y134_SLICE_X7Y134_CQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C5 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_C6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_D1 = CLBLM_R_X3Y141_SLICE_X3Y141_BO6;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_D1 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_T1 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D2 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D3 = CLBLL_L_X4Y136_SLICE_X5Y136_DQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D4 = CLBLM_R_X3Y141_SLICE_X2Y141_BQ;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D5 = CLBLM_R_X7Y136_SLICE_X8Y136_A5Q;
  assign CLBLM_R_X5Y136_SLICE_X7Y136_D6 = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_T1 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_D1 = CLBLM_L_X10Y134_SLICE_X12Y134_B5Q;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A1 = CLBLM_R_X5Y134_SLICE_X6Y134_B5Q;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A2 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A3 = CLBLM_R_X5Y136_SLICE_X6Y136_AQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A5 = CLBLM_R_X5Y136_SLICE_X7Y136_AQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_A6 = CLBLM_R_X11Y131_SLICE_X14Y131_BO6;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_T1 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B1 = CLBLM_R_X5Y141_SLICE_X6Y141_DQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B3 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B4 = CLBLL_L_X4Y133_SLICE_X4Y133_CQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B5 = CLBLM_L_X10Y140_SLICE_X13Y140_B5Q;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_B6 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C2 = CLBLL_L_X4Y134_SLICE_X4Y134_BQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C3 = CLBLM_L_X12Y132_SLICE_X16Y132_AO6;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C4 = CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C5 = CLBLM_R_X5Y136_SLICE_X6Y136_CQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_C6 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_T1 = 1'b1;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D2 = CLBLM_R_X5Y136_SLICE_X6Y136_CQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D3 = CLBLM_R_X3Y136_SLICE_X2Y136_CQ;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D4 = CLBLL_L_X4Y136_SLICE_X4Y136_B5Q;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D5 = CLBLL_L_X4Y134_SLICE_X4Y134_C5Q;
  assign CLBLM_R_X5Y136_SLICE_X6Y136_D6 = CLBLL_L_X4Y135_SLICE_X4Y135_AQ;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_D1 = CLBLM_R_X3Y137_SLICE_X2Y137_DO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_T1 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D1 = CLBLM_L_X10Y140_SLICE_X13Y140_C5Q;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_D = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_D = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOB33_X0Y167_IOB_X0Y168_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign LIOB33_X0Y167_IOB_X0Y167_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D2 = CLBLM_L_X8Y138_SLICE_X10Y138_BQ;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_C4 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_C5 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_C6 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A2 = CLBLM_R_X7Y137_SLICE_X8Y137_D5Q;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A3 = CLBLL_L_X4Y140_SLICE_X5Y140_AQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A4 = CLBLL_L_X4Y134_SLICE_X4Y134_C5Q;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A5 = CLBLM_L_X8Y137_SLICE_X10Y137_AQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_A6 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B1 = CLBLL_L_X4Y137_SLICE_X4Y137_DO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B2 = CLBLM_L_X8Y139_SLICE_X10Y139_AO6;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B4 = CLBLM_R_X5Y136_SLICE_X7Y136_D5Q;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B5 = CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_B6 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C1 = CLBLM_R_X5Y134_SLICE_X7Y134_A5Q;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C2 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C3 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C4 = CLBLM_R_X7Y138_SLICE_X8Y138_DQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C5 = CLBLM_R_X5Y135_SLICE_X7Y135_DQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_C6 = CLBLM_R_X7Y133_SLICE_X9Y133_BQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D1 = CLBLM_L_X8Y137_SLICE_X10Y137_CQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D2 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D3 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D4 = CLBLM_R_X3Y141_SLICE_X2Y141_BQ;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D5 = CLBLL_L_X4Y132_SLICE_X5Y132_C5Q;
  assign CLBLM_R_X5Y137_SLICE_X7Y137_D6 = CLBLM_R_X5Y136_SLICE_X7Y136_D5Q;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_D5 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A1 = CLBLM_R_X3Y136_SLICE_X2Y136_CQ;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_D6 = 1'b1;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A2 = CLBLM_R_X5Y137_SLICE_X6Y137_BQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A4 = CLBLL_L_X4Y134_SLICE_X5Y134_CQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A5 = CLBLL_L_X4Y135_SLICE_X4Y135_AQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_A6 = CLBLM_R_X11Y142_SLICE_X14Y142_AQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B2 = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B3 = CLBLL_L_X4Y131_SLICE_X5Y131_B5Q;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B4 = CLBLM_R_X5Y137_SLICE_X6Y137_CQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B5 = CLBLL_L_X4Y135_SLICE_X4Y135_AQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_B6 = CLBLM_R_X3Y136_SLICE_X2Y136_CQ;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_D = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C1 = CLBLL_L_X4Y135_SLICE_X4Y135_AQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C2 = CLBLM_R_X7Y137_SLICE_X8Y137_C5Q;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C3 = CLBLM_L_X12Y136_SLICE_X16Y136_A5Q;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C4 = CLBLM_R_X5Y136_SLICE_X6Y136_DQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_C6 = CLBLM_R_X3Y136_SLICE_X2Y136_CQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_D = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D1 = CLBLM_R_X3Y135_SLICE_X3Y135_CQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D2 = CLBLM_R_X3Y135_SLICE_X3Y135_BQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D3 = CLBLL_L_X4Y138_SLICE_X5Y138_DQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D4 = CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D5 = CLBLL_L_X4Y137_SLICE_X5Y137_C5Q;
  assign CLBLM_R_X5Y137_SLICE_X6Y137_D6 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_C4 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_C5 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_C6 = 1'b1;
  assign LIOB33_X0Y169_IOB_X0Y169_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOB33_X0Y169_IOB_X0Y170_O = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A1 = CLBLM_R_X5Y138_SLICE_X7Y138_DO6;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A3 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A4 = CLBLM_L_X8Y137_SLICE_X10Y137_C5Q;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A5 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_A6 = CLBLM_R_X5Y139_SLICE_X7Y139_CQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B1 = CLBLM_R_X5Y132_SLICE_X6Y132_AQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B2 = CLBLM_R_X5Y137_SLICE_X7Y137_BQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B3 = CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B4 = CLBLM_R_X5Y134_SLICE_X6Y134_CQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B5 = CLBLM_R_X7Y138_SLICE_X9Y138_B5Q;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_B6 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C1 = CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C2 = CLBLL_L_X4Y137_SLICE_X5Y137_C5Q;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C3 = CLBLM_R_X5Y134_SLICE_X6Y134_DQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C4 = CLBLM_R_X5Y140_SLICE_X6Y140_CQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C5 = CLBLM_R_X5Y138_SLICE_X7Y138_BO5;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_C6 = CLBLM_R_X5Y137_SLICE_X6Y137_DO5;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D1 = CLBLM_R_X3Y135_SLICE_X3Y135_DQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D2 = CLBLM_R_X5Y140_SLICE_X6Y140_CQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D3 = CLBLM_R_X7Y138_SLICE_X9Y138_B5Q;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D4 = CLBLM_R_X5Y134_SLICE_X6Y134_DQ;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D5 = CLBLM_R_X5Y138_SLICE_X7Y138_BO5;
  assign CLBLM_R_X5Y138_SLICE_X7Y138_D6 = CLBLM_R_X5Y137_SLICE_X7Y137_BQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A1 = CLBLM_R_X5Y139_SLICE_X7Y139_CQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A2 = CLBLM_R_X7Y133_SLICE_X9Y133_CQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A3 = CLBLM_R_X5Y138_SLICE_X7Y138_DO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A5 = CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_A6 = CLBLL_L_X4Y138_SLICE_X5Y138_B5Q;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B1 = CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B2 = CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B3 = CLBLM_L_X8Y138_SLICE_X10Y138_BQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B5 = CLBLL_L_X2Y138_SLICE_X1Y138_BO6;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_B6 = 1'b1;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C1 = CLBLM_R_X5Y140_SLICE_X6Y140_AQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C3 = CLBLM_R_X5Y137_SLICE_X6Y137_AQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C4 = CLBLM_R_X3Y136_SLICE_X2Y136_CQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C5 = CLBLL_L_X4Y135_SLICE_X4Y135_AQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_C6 = CLBLM_L_X10Y140_SLICE_X13Y140_BQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D1 = CLBLM_R_X5Y137_SLICE_X6Y137_DO5;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D2 = CLBLL_L_X4Y137_SLICE_X5Y137_C5Q;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D4 = CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D5 = CLBLM_R_X5Y137_SLICE_X6Y137_AQ;
  assign CLBLM_R_X5Y138_SLICE_X6Y138_D6 = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_D1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign LIOB33_X0Y179_IOB_X0Y180_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign LIOB33_X0Y179_IOB_X0Y179_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_T1 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D5 = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_D1 = CLBLL_L_X4Y132_SLICE_X5Y132_BQ;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C3 = CLBLM_L_X8Y140_SLICE_X10Y140_CQ;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_D1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C4 = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_D1 = 1'b1;
  assign RIOB33_X105Y161_IOB_X1Y162_O = CLBLM_R_X7Y140_SLICE_X9Y140_D5Q;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C5 = CLBLM_R_X7Y133_SLICE_X8Y133_A5Q;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_T1 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C6 = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_D1 = CLBLL_L_X4Y137_SLICE_X5Y137_B5Q;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1 = CLBLM_R_X3Y141_SLICE_X2Y141_BQ;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_D1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1 = CLBLL_L_X4Y130_SLICE_X4Y130_DQ;
  assign LIOB33_X0Y171_IOB_X0Y172_O = RIOB33_X105Y119_IOB_X1Y120_I;
  assign LIOB33_X0Y171_IOB_X0Y171_O = RIOB33_X105Y119_IOB_X1Y119_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D2 = CLBLM_R_X13Y137_SLICE_X18Y137_AO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D5 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D6 = CLBLM_L_X10Y133_SLICE_X12Y133_BQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A1 = CLBLM_R_X3Y136_SLICE_X2Y136_B5Q;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A2 = CLBLM_L_X8Y140_SLICE_X11Y140_CQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A4 = CLBLM_R_X5Y137_SLICE_X7Y137_BQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A5 = CLBLM_L_X8Y131_SLICE_X11Y131_CQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_A6 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C4 = CLBLM_R_X5Y140_SLICE_X7Y140_A5Q;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B1 = CLBLM_R_X3Y139_SLICE_X3Y139_DO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B2 = CLBLM_L_X8Y138_SLICE_X10Y138_C5Q;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B4 = CLBLM_R_X7Y136_SLICE_X8Y136_C5Q;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B5 = CLBLM_R_X5Y138_SLICE_X6Y138_CQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_B6 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_C6 = CLBLM_L_X10Y134_SLICE_X12Y134_AQ;
  assign LIOB33_X0Y197_IOB_X0Y198_O = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C1 = CLBLM_R_X5Y137_SLICE_X6Y137_DO5;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C2 = CLBLL_L_X4Y137_SLICE_X5Y137_C5Q;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C3 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C4 = CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C5 = CLBLM_R_X5Y137_SLICE_X7Y137_AQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D1 = CLBLM_R_X5Y140_SLICE_X7Y140_AQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D2 = CLBLM_R_X7Y140_SLICE_X8Y140_B5Q;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D3 = CLBLM_L_X8Y133_SLICE_X11Y133_BQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D4 = CLBLM_R_X3Y136_SLICE_X3Y136_CQ;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D5 = CLBLM_R_X7Y139_SLICE_X8Y139_CO6;
  assign CLBLM_R_X5Y139_SLICE_X7Y139_D6 = CLBLM_R_X5Y139_SLICE_X6Y139_C5Q;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B6 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A1 = CLBLM_R_X11Y140_SLICE_X15Y140_BQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A3 = CLBLM_R_X5Y139_SLICE_X6Y139_AQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A4 = CLBLM_L_X12Y132_SLICE_X16Y132_AO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A5 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_A6 = CLBLL_L_X4Y139_SLICE_X5Y139_AQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_BX = CLBLL_L_X4Y136_SLICE_X4Y136_BQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B1 = CLBLM_R_X5Y139_SLICE_X6Y139_DO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B2 = CLBLM_R_X5Y130_SLICE_X6Y130_AQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B3 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B4 = CLBLM_R_X7Y136_SLICE_X9Y136_BQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B5 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C1 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D2 = CLBLM_R_X3Y140_SLICE_X3Y140_CQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C1 = CLBLM_R_X5Y140_SLICE_X7Y140_AQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C2 = CLBLL_L_X4Y130_SLICE_X5Y130_AQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C4 = CLBLM_R_X5Y132_SLICE_X6Y132_AQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C5 = CLBLM_R_X7Y140_SLICE_X8Y140_DQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_C6 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C2 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C3 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C4 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D5 = CLBLM_L_X8Y142_SLICE_X10Y142_CO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D1 = CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D2 = CLBLL_L_X4Y138_SLICE_X5Y138_B5Q;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D3 = CLBLM_R_X5Y138_SLICE_X7Y138_DO6;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D4 = CLBLM_R_X5Y139_SLICE_X7Y139_CQ;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D5 = 1'b1;
  assign CLBLM_R_X5Y139_SLICE_X6Y139_D6 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X9Y142_D6 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C5 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_C6 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A1 = CLBLM_L_X8Y136_SLICE_X10Y136_AO5;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D5 = CLBLM_R_X7Y134_SLICE_X9Y134_CQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D6 = CLBLM_L_X12Y132_SLICE_X16Y132_AO6;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_CX = CLBLM_R_X5Y140_SLICE_X7Y140_CQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D1 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_A5 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D2 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D3 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B2 = CLBLM_L_X10Y140_SLICE_X12Y140_D5Q;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D4 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B3 = CLBLM_R_X5Y139_SLICE_X6Y139_C5Q;
  assign LIOB33_X0Y173_IOB_X0Y173_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOB33_X0Y173_IOB_X0Y174_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D5 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A1 = CLBLM_R_X7Y139_SLICE_X9Y139_AQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_D6 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A2 = CLBLM_L_X8Y132_SLICE_X11Y132_AQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A3 = CLBLM_L_X10Y132_SLICE_X12Y132_C5Q;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_DX = CLBLM_L_X8Y138_SLICE_X10Y138_A5Q;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B4 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B5 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_B6 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C3 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C4 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C6 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C3 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C4 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C5 = 1'b1;
  assign CLBLM_R_X7Y142_SLICE_X8Y142_C6 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_T1 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A1 = CLBLL_L_X4Y138_SLICE_X5Y138_DQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A2 = CLBLM_R_X5Y140_SLICE_X7Y140_BQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A4 = CLBLM_R_X3Y140_SLICE_X3Y140_DQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A5 = CLBLM_L_X10Y140_SLICE_X12Y140_DQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_A6 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B1 = CLBLM_R_X5Y138_SLICE_X7Y138_DO6;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B3 = CLBLM_R_X5Y140_SLICE_X7Y140_CQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B4 = CLBLL_L_X4Y142_SLICE_X5Y142_A5Q;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B5 = CLBLM_L_X10Y134_SLICE_X12Y134_A5Q;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_B6 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A1 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A2 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A3 = CLBLL_L_X4Y131_SLICE_X4Y131_D5Q;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A4 = CLBLM_R_X3Y130_SLICE_X3Y130_BO6;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A5 = CLBLM_R_X5Y133_SLICE_X7Y133_CQ;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_A6 = CLBLL_L_X4Y130_SLICE_X4Y130_BQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C1 = CLBLL_L_X4Y137_SLICE_X5Y137_C5Q;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C2 = CLBLM_R_X5Y135_SLICE_X7Y135_D5Q;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B1 = CLBLL_L_X4Y130_SLICE_X4Y130_DQ;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B2 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B3 = CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B4 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B5 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_B6 = CLBLL_L_X4Y132_SLICE_X5Y132_A5Q;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D1 = CLBLL_L_X4Y137_SLICE_X5Y137_C5Q;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C1 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C2 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C3 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C4 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C5 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_C6 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D3 = CLBLM_R_X5Y137_SLICE_X6Y137_DO5;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D4 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A1 = CLBLM_R_X5Y133_SLICE_X7Y133_AQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A2 = CLBLM_L_X8Y138_SLICE_X10Y138_DQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A3 = CLBLM_R_X5Y140_SLICE_X6Y140_AQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A5 = CLBLL_L_X4Y139_SLICE_X5Y139_C5Q;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_A6 = CLBLL_L_X4Y135_SLICE_X4Y135_D5Q;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D1 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D2 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D3 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D4 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D5 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X3Y130_D6 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_AX = CLBLM_R_X5Y140_SLICE_X6Y140_BO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B2 = CLBLM_R_X5Y139_SLICE_X7Y139_DO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B3 = CLBLM_R_X5Y131_SLICE_X6Y131_BQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B4 = CLBLM_R_X5Y137_SLICE_X7Y137_CO6;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B5 = CLBLM_L_X10Y137_SLICE_X13Y137_AQ;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A1 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A2 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A3 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A4 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A5 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_A6 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C1 = CLBLM_R_X5Y130_SLICE_X7Y130_DQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C2 = CLBLM_R_X5Y140_SLICE_X6Y140_CQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C3 = CLBLM_R_X5Y140_SLICE_X7Y140_DO6;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B1 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B2 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B3 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B4 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B5 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_B6 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D1 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D2 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C1 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C2 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C3 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C4 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C5 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_C6 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D3 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D4 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D5 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_D6 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D1 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D2 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D3 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D4 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D5 = 1'b1;
  assign CLBLM_R_X3Y130_SLICE_X2Y130_D6 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_T1 = 1'b1;
  assign LIOB33_X0Y175_IOB_X0Y176_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOB33_X0Y175_IOB_X0Y175_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_D1 = RIOB33_X105Y119_IOB_X1Y120_I;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_D = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_T1 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_D1 = CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_D1 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_T1 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_D1 = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_T1 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_D1 = CLBLL_L_X4Y130_SLICE_X4Y130_BQ;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = CLBLM_R_X3Y139_SLICE_X3Y139_A5Q;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_T1 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_D1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = CLBLM_R_X7Y137_SLICE_X9Y137_D5Q;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A1 = CLBLM_L_X8Y136_SLICE_X10Y136_BQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A2 = CLBLM_R_X7Y141_SLICE_X9Y141_A5Q;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A3 = CLBLM_R_X3Y135_SLICE_X2Y135_AQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A4 = CLBLM_R_X5Y141_SLICE_X7Y141_BO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A5 = CLBLM_L_X10Y130_SLICE_X12Y130_B5Q;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_A6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B1 = CLBLM_R_X5Y141_SLICE_X7Y141_DO6;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B2 = CLBLM_R_X3Y135_SLICE_X2Y135_AQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B3 = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B4 = CLBLM_L_X8Y136_SLICE_X10Y136_BQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B5 = CLBLL_L_X4Y140_SLICE_X4Y140_BO5;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_B6 = CLBLM_L_X10Y137_SLICE_X12Y137_AQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A1 = CLBLM_R_X5Y134_SLICE_X6Y134_AQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A2 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A3 = CLBLL_L_X4Y130_SLICE_X5Y130_CO5;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A4 = CLBLM_R_X3Y131_SLICE_X3Y131_AQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A5 = CLBLM_R_X5Y130_SLICE_X6Y130_B5Q;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C1 = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C2 = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C3 = CLBLM_R_X11Y139_SLICE_X14Y139_AO5;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B1 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B2 = CLBLM_R_X3Y131_SLICE_X3Y131_BQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B3 = CLBLM_R_X7Y138_SLICE_X9Y138_B5Q;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B4 = CLBLM_R_X5Y135_SLICE_X7Y135_AQ;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_B6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D1 = CLBLM_R_X5Y143_SLICE_X7Y143_AQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D2 = CLBLL_L_X4Y143_SLICE_X5Y143_DO6;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C2 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C3 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C4 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_C6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D3 = CLBLM_L_X10Y137_SLICE_X12Y137_AQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D4 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A1 = CLBLM_R_X5Y138_SLICE_X7Y138_DO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A2 = CLBLM_R_X5Y142_SLICE_X6Y142_BQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A3 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D2 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D3 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D4 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X3Y131_D6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_A6 = CLBLL_L_X4Y138_SLICE_X5Y138_B5Q;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B1 = CLBLM_R_X5Y141_SLICE_X6Y141_CQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B2 = CLBLM_L_X10Y140_SLICE_X13Y140_DQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B4 = CLBLM_R_X5Y139_SLICE_X7Y139_BQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A1 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A2 = CLBLM_R_X3Y131_SLICE_X2Y131_BQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A3 = CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A4 = CLBLM_R_X3Y131_SLICE_X3Y131_BQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_A6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C1 = CLBLM_R_X5Y141_SLICE_X6Y141_BQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C2 = CLBLM_R_X5Y139_SLICE_X7Y139_BQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C3 = CLBLM_R_X5Y142_SLICE_X6Y142_BQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B2 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B3 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B4 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_B6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D1 = CLBLL_L_X4Y140_SLICE_X4Y140_BO5;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D2 = CLBLM_R_X5Y141_SLICE_X7Y141_AO6;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_BX = CLBLM_R_X3Y132_SLICE_X2Y132_CO5;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D3 = CLBLM_R_X5Y141_SLICE_X6Y141_DQ;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C2 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C3 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C4 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_C6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D5 = CLBLM_R_X7Y140_SLICE_X8Y140_CQ;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_D6 = CLBLL_L_X4Y142_SLICE_X5Y142_A5Q;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y177_IOB_X0Y178_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign LIOB33_X0Y177_IOB_X0Y177_O = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D1 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D2 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D3 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D4 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D5 = 1'b1;
  assign CLBLM_R_X3Y131_SLICE_X2Y131_D6 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A5 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B2 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B3 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B4 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B5 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B6 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C1 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C2 = 1'b1;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_D = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C3 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C4 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_T1 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C5 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_C6 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A1 = CLBLM_R_X5Y142_SLICE_X7Y142_BO5;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A2 = CLBLL_L_X4Y137_SLICE_X5Y137_A5Q;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A3 = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A4 = CLBLM_R_X5Y142_SLICE_X7Y142_BO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A5 = CLBLM_R_X5Y141_SLICE_X7Y141_AO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B1 = CLBLM_R_X5Y141_SLICE_X6Y141_DQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B2 = CLBLL_L_X4Y140_SLICE_X4Y140_CO5;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B3 = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B4 = CLBLL_L_X4Y142_SLICE_X5Y142_A5Q;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B5 = CLBLL_L_X4Y140_SLICE_X4Y140_BO5;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_B6 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A1 = CLBLL_L_X4Y132_SLICE_X4Y132_CQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A2 = CLBLL_L_X4Y132_SLICE_X4Y132_AQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A3 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A4 = CLBLL_L_X4Y132_SLICE_X4Y132_BQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A5 = CLBLM_R_X7Y137_SLICE_X8Y137_B5Q;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C3 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_C4 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B1 = CLBLL_L_X4Y132_SLICE_X4Y132_CQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B2 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B3 = CLBLM_R_X3Y138_SLICE_X3Y138_A5Q;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B4 = CLBLL_L_X4Y132_SLICE_X4Y132_AQ;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D1 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B5 = CLBLL_L_X4Y132_SLICE_X4Y132_BQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D2 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C2 = CLBLM_R_X3Y132_SLICE_X3Y132_CQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C3 = CLBLL_L_X4Y132_SLICE_X4Y132_DQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C4 = CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D3 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C5 = CLBLM_R_X3Y139_SLICE_X3Y139_A5Q;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_C6 = CLBLM_L_X8Y132_SLICE_X11Y132_CO6;
  assign CLBLM_R_X5Y142_SLICE_X7Y142_D4 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A2 = CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A3 = CLBLM_R_X5Y142_SLICE_X6Y142_AQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A4 = CLBLM_R_X5Y135_SLICE_X6Y135_B5Q;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D5 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D2 = CLBLL_L_X4Y130_SLICE_X4Y130_B5Q;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D3 = CLBLM_R_X3Y135_SLICE_X3Y135_BQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D4 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D6 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D5 = CLBLM_R_X3Y133_SLICE_X2Y133_BQ;
  assign CLBLM_R_X3Y132_SLICE_X3Y132_D6 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_A6 = CLBLL_L_X4Y135_SLICE_X5Y135_CQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B1 = CLBLL_L_X4Y143_SLICE_X5Y143_AQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_B3 = CLBLM_R_X7Y140_SLICE_X8Y140_DQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A1 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A2 = CLBLL_L_X4Y135_SLICE_X5Y135_CQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A3 = CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A4 = CLBLL_L_X4Y135_SLICE_X4Y135_CQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_A6 = CLBLM_L_X8Y132_SLICE_X11Y132_BQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C1 = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_C2 = CLBLM_R_X5Y142_SLICE_X6Y142_CQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B1 = CLBLM_R_X3Y132_SLICE_X3Y132_DQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B2 = CLBLM_R_X3Y132_SLICE_X2Y132_BQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B3 = CLBLM_R_X7Y131_SLICE_X9Y131_D5Q;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B5 = CLBLM_L_X10Y140_SLICE_X13Y140_D5Q;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_B6 = CLBLM_R_X5Y133_SLICE_X6Y133_A5Q;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D1 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D2 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C2 = CLBLM_R_X3Y131_SLICE_X3Y131_BQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C3 = CLBLM_R_X3Y132_SLICE_X2Y132_BQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C4 = CLBLM_R_X3Y131_SLICE_X2Y131_BQ;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C5 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_C6 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D3 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D4 = 1'b1;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D5 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y142_SLICE_X6Y142_D6 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D1 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D2 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D3 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D4 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D5 = 1'b1;
  assign CLBLM_R_X3Y132_SLICE_X2Y132_D6 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A6 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B4 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B5 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B6 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C1 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C2 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C3 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C4 = 1'b1;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C5 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_C6 = 1'b1;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1 = 1'b1;
  assign LIOB33_X0Y181_IOB_X0Y182_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D1 = 1'b1;
  assign LIOB33_X0Y181_IOB_X0Y181_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D2 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D3 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D4 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D5 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A1 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_D6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A3 = CLBLM_R_X5Y143_SLICE_X7Y143_AQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A4 = CLBLL_L_X4Y143_SLICE_X5Y143_CO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A5 = CLBLM_R_X5Y141_SLICE_X7Y141_AO6;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_A6 = CLBLM_R_X7Y138_SLICE_X9Y138_BQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B1 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B2 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B3 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B4 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B5 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_B6 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A1 = CLBLL_L_X4Y130_SLICE_X4Y130_AQ;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A2 = CLBLL_L_X4Y133_SLICE_X4Y133_CQ;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A3 = CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A4 = CLBLM_R_X7Y131_SLICE_X9Y131_D5Q;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A5 = CLBLM_L_X10Y140_SLICE_X13Y140_D5Q;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C1 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_C2 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B1 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B2 = CLBLM_R_X7Y136_SLICE_X9Y136_A5Q;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B4 = CLBLL_L_X4Y132_SLICE_X5Y132_BQ;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B5 = CLBLL_L_X4Y134_SLICE_X4Y134_C5Q;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_B6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D1 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C1 = CLBLM_L_X8Y140_SLICE_X11Y140_BQ;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C2 = CLBLL_L_X4Y132_SLICE_X5Y132_CQ;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C3 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C4 = CLBLM_R_X5Y132_SLICE_X6Y132_CO6;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C5 = CLBLM_R_X3Y134_SLICE_X3Y134_AQ;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_C6 = CLBLM_R_X3Y134_SLICE_X3Y134_BQ;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D3 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X7Y143_D4 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A1 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A2 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A3 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A4 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A5 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D1 = CLBLM_R_X3Y131_SLICE_X2Y131_BQ;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D2 = CLBLM_R_X3Y131_SLICE_X3Y131_BQ;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D3 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D4 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D5 = CLBLM_R_X5Y135_SLICE_X6Y135_A5Q;
  assign CLBLM_R_X3Y133_SLICE_X3Y133_D6 = CLBLM_R_X3Y134_SLICE_X3Y134_BQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_A6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B1 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B2 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B3 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_B4 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A1 = CLBLM_R_X3Y141_SLICE_X2Y141_CO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A2 = CLBLL_L_X4Y133_SLICE_X5Y133_DQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A3 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A4 = CLBLM_R_X3Y133_SLICE_X2Y133_DO6;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_A6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C1 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C2 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_C3 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B1 = CLBLL_L_X4Y133_SLICE_X5Y133_CQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B2 = CLBLM_R_X3Y133_SLICE_X2Y133_BQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B3 = CLBLL_L_X4Y132_SLICE_X5Y132_DQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B4 = CLBLL_L_X4Y135_SLICE_X5Y135_CQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_B6 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D1 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D2 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D3 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C1 = CLBLM_L_X8Y140_SLICE_X11Y140_BQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C2 = CLBLM_R_X3Y131_SLICE_X2Y131_BQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C3 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C4 = CLBLM_R_X3Y134_SLICE_X3Y134_AQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C5 = CLBLM_R_X3Y131_SLICE_X3Y131_BQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_C6 = CLBLM_R_X3Y134_SLICE_X3Y134_BQ;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D6 = 1'b1;
  assign CLBLM_R_X5Y143_SLICE_X6Y143_D4 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1 = CLBLM_R_X5Y140_SLICE_X6Y140_BO5;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D1 = 1'b1;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D4 = CLBLM_R_X7Y134_SLICE_X8Y134_CQ;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X3Y133_SLICE_X2Y133_D6 = CLBLL_L_X4Y138_SLICE_X4Y138_BQ;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C1 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C5 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C6 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D2 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D5 = 1'b1;
  assign LIOB33_X0Y63_IOB_X0Y64_O = CLBLL_L_X2Y134_SLICE_X1Y134_AO5;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D6 = 1'b1;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_D = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_D = LIOB33_X0Y51_IOB_X0Y51_I;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign RIOB33_X105Y151_IOB_X1Y152_O = 1'b1;
  assign RIOB33_X105Y151_IOB_X1Y151_O = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOB33_X0Y183_IOB_X0Y184_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign LIOB33_X0Y183_IOB_X0Y183_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C4 = CLBLM_L_X8Y143_SLICE_X10Y143_BO5;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C5 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_A2 = CLBLM_R_X3Y134_SLICE_X2Y134_BO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_A3 = CLBLM_R_X11Y141_SLICE_X14Y141_AQ;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_A4 = CLBLM_L_X8Y139_SLICE_X11Y139_BQ;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_A5 = CLBLM_R_X3Y133_SLICE_X2Y133_CO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_A6 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_C6 = CLBLM_L_X8Y141_SLICE_X11Y141_BQ;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_B1 = CLBLM_R_X3Y134_SLICE_X3Y134_DO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_B2 = CLBLM_R_X5Y135_SLICE_X6Y135_A5Q;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_B3 = CLBLM_R_X3Y134_SLICE_X2Y134_AO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_B4 = CLBLM_R_X3Y140_SLICE_X3Y140_CQ;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_B6 = CLBLM_R_X3Y134_SLICE_X3Y134_CO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_C1 = CLBLM_L_X8Y140_SLICE_X11Y140_BQ;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_C2 = CLBLM_R_X3Y130_SLICE_X3Y130_AO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_C3 = CLBLM_R_X3Y134_SLICE_X3Y134_BQ;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_C4 = CLBLM_R_X3Y132_SLICE_X2Y132_CO6;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_C5 = CLBLM_R_X3Y134_SLICE_X3Y134_AQ;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_C6 = CLBLM_R_X7Y132_SLICE_X8Y132_D5Q;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B5 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B6 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_SING_X105Y150_IOB_X1Y150_O = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_D1 = CLBLM_L_X8Y140_SLICE_X11Y140_BQ;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_D2 = CLBLM_R_X7Y132_SLICE_X8Y132_D5Q;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_D3 = CLBLM_R_X3Y135_SLICE_X2Y135_DQ;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_D4 = CLBLM_R_X3Y134_SLICE_X3Y134_BQ;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_D5 = CLBLM_R_X3Y134_SLICE_X3Y134_AQ;
  assign CLBLM_R_X3Y134_SLICE_X3Y134_D6 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_A1 = CLBLM_R_X3Y134_SLICE_X3Y134_BQ;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_A2 = CLBLM_R_X3Y131_SLICE_X2Y131_AQ;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_A3 = CLBLM_L_X8Y140_SLICE_X11Y140_BQ;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_A4 = CLBLM_R_X3Y132_SLICE_X2Y132_CO6;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_A5 = CLBLM_R_X3Y134_SLICE_X3Y134_AQ;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_A6 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_AX = CLBLM_R_X3Y134_SLICE_X3Y134_AQ;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_B1 = CLBLM_R_X3Y134_SLICE_X3Y134_BQ;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_B2 = CLBLM_R_X7Y132_SLICE_X8Y132_D5Q;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_B3 = CLBLM_R_X3Y134_SLICE_X3Y134_AQ;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_B4 = CLBLM_R_X5Y135_SLICE_X6Y135_A5Q;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_B5 = CLBLM_R_X3Y130_SLICE_X3Y130_AO6;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_B6 = CLBLM_R_X3Y132_SLICE_X2Y132_CO6;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D2 = CLBLM_R_X7Y133_SLICE_X8Y133_A5Q;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_C1 = CLBLM_L_X8Y140_SLICE_X11Y140_BQ;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_C2 = CLBLM_R_X3Y134_SLICE_X3Y134_AQ;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_C3 = CLBLM_R_X7Y132_SLICE_X8Y132_D5Q;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_C4 = CLBLM_R_X3Y132_SLICE_X2Y132_CO6;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_C5 = CLBLM_R_X3Y134_SLICE_X2Y134_DO6;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_C6 = CLBLM_R_X3Y134_SLICE_X3Y134_BQ;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D5 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C4 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y143_SLICE_X9Y143_D6 = CLBLM_L_X8Y141_SLICE_X11Y141_BQ;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C5 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C6 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_D1 = CLBLM_L_X8Y140_SLICE_X11Y140_BQ;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_D2 = CLBLM_R_X3Y134_SLICE_X3Y134_AQ;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_D3 = CLBLM_R_X7Y137_SLICE_X9Y137_D5Q;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_D4 = 1'b1;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_D5 = CLBLM_R_X3Y135_SLICE_X2Y135_DQ;
  assign CLBLM_R_X3Y134_SLICE_X2Y134_D6 = CLBLM_R_X3Y134_SLICE_X3Y134_BQ;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_A6 = CLBLM_R_X7Y143_SLICE_X9Y143_DO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A1 = CLBLM_L_X10Y135_SLICE_X12Y135_B5Q;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A2 = CLBLM_L_X10Y138_SLICE_X13Y138_CQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A3 = CLBLL_L_X4Y134_SLICE_X4Y134_C5Q;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_B2 = CLBLM_R_X7Y143_SLICE_X9Y143_DO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOB33_X0Y65_IOB_X0Y66_O = CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  assign LIOB33_X0Y65_IOB_X0Y65_O = CLBLL_L_X2Y133_SLICE_X1Y133_BO6;
  assign LIOB33_X0Y111_IOB_X0Y112_O = CLBLL_L_X4Y132_SLICE_X5Y132_A5Q;
  assign LIOB33_X0Y111_IOB_X0Y111_O = CLBLL_L_X4Y131_SLICE_X4Y131_D5Q;
  assign RIOB33_X105Y153_IOB_X1Y154_O = 1'b1;
  assign RIOB33_X105Y153_IOB_X1Y153_O = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C4 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C5 = 1'b1;
  assign CLBLM_R_X7Y143_SLICE_X8Y143_C6 = 1'b1;
  assign LIOB33_X0Y185_IOB_X0Y186_O = RIOB33_X105Y119_IOB_X1Y120_I;
  assign LIOB33_X0Y185_IOB_X0Y185_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOB33_X0Y159_IOB_X0Y160_O = CLBLM_R_X3Y134_SLICE_X2Y134_AQ;
  assign LIOB33_X0Y159_IOB_X0Y159_O = CLBLM_R_X3Y132_SLICE_X3Y132_BQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_A1 = CLBLM_R_X3Y140_SLICE_X3Y140_C5Q;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_A2 = CLBLM_R_X3Y132_SLICE_X3Y132_DQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_A3 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_A5 = CLBLM_L_X12Y136_SLICE_X16Y136_AQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_A6 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_B1 = CLBLM_R_X5Y134_SLICE_X7Y134_A5Q;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_B2 = CLBLM_R_X3Y135_SLICE_X3Y135_BQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_B3 = CLBLM_R_X3Y135_SLICE_X3Y135_CQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_B5 = CLBLM_R_X5Y135_SLICE_X6Y135_DO6;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_B6 = CLBLM_R_X5Y130_SLICE_X7Y130_DQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_C2 = CLBLM_R_X5Y130_SLICE_X7Y130_DQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_C3 = CLBLM_R_X5Y135_SLICE_X6Y135_DO6;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_C4 = CLBLM_R_X3Y135_SLICE_X3Y135_A5Q;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_C5 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_C6 = CLBLM_R_X3Y135_SLICE_X3Y135_CQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_D1 = CLBLL_L_X4Y138_SLICE_X4Y138_DO6;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_D2 = CLBLM_R_X5Y130_SLICE_X7Y130_DQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_D3 = CLBLM_R_X3Y135_SLICE_X3Y135_DQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_D5 = CLBLM_R_X5Y138_SLICE_X7Y138_AQ;
  assign CLBLM_R_X3Y135_SLICE_X3Y135_D6 = CLBLM_R_X3Y133_SLICE_X3Y133_BQ;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_A1 = 1'b1;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_A2 = CLBLM_R_X7Y132_SLICE_X9Y132_BQ;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_A3 = CLBLM_R_X3Y135_SLICE_X2Y135_AQ;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_A4 = CLBLM_R_X3Y137_SLICE_X2Y137_BO6;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_A5 = CLBLL_L_X4Y135_SLICE_X5Y135_DO6;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_B1 = CLBLM_R_X7Y131_SLICE_X9Y131_D5Q;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_B2 = CLBLM_R_X3Y135_SLICE_X2Y135_BQ;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_B3 = CLBLM_R_X5Y139_SLICE_X7Y139_AQ;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_B4 = CLBLM_L_X10Y140_SLICE_X13Y140_D5Q;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_B5 = CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_C1 = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_C2 = CLBLM_R_X3Y135_SLICE_X2Y135_CQ;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_C3 = CLBLL_L_X4Y133_SLICE_X4Y133_DQ;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_C4 = CLBLM_L_X8Y138_SLICE_X10Y138_CQ;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_C6 = CLBLL_L_X4Y136_SLICE_X4Y136_D5Q;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_D1 = CLBLM_L_X8Y140_SLICE_X11Y140_BQ;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_D3 = CLBLM_R_X3Y134_SLICE_X3Y134_AQ;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_D4 = CLBLM_R_X7Y137_SLICE_X9Y137_D5Q;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_D5 = CLBLM_R_X3Y136_SLICE_X3Y136_CQ;
  assign CLBLM_R_X3Y135_SLICE_X2Y135_D6 = CLBLM_R_X3Y134_SLICE_X3Y134_BQ;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_D1 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_T1 = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_D1 = CLBLM_L_X10Y131_SLICE_X12Y131_D5Q;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_D1 = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_T1 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_D1 = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_T1 = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_D1 = CLBLM_R_X5Y138_SLICE_X6Y138_B5Q;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1 = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_T1 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_D1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_T1 = 1'b1;
  assign RIOB33_X105Y155_IOB_X1Y156_O = 1'b1;
  assign RIOB33_X105Y155_IOB_X1Y155_O = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1 = CLBLM_R_X3Y135_SLICE_X2Y135_AQ;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1 = 1'b1;
  assign LIOB33_X0Y187_IOB_X0Y188_O = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign LIOB33_X0Y187_IOB_X0Y187_O = CLBLM_R_X3Y135_SLICE_X2Y135_AQ;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B5 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_A1 = CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_A2 = CLBLM_R_X3Y138_SLICE_X2Y138_BQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_A3 = CLBLM_R_X3Y136_SLICE_X3Y136_AQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_A5 = CLBLM_L_X8Y139_SLICE_X11Y139_BQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_A6 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_B2 = CLBLM_R_X5Y136_SLICE_X7Y136_C5Q;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_B3 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_B4 = CLBLM_L_X10Y140_SLICE_X13Y140_BQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_B5 = CLBLL_L_X4Y133_SLICE_X5Y133_BQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_B6 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_C1 = CLBLM_R_X7Y136_SLICE_X9Y136_A5Q;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_C2 = CLBLL_L_X4Y134_SLICE_X5Y134_DQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_C3 = CLBLM_R_X7Y132_SLICE_X8Y132_BQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_C4 = CLBLM_R_X3Y135_SLICE_X3Y135_CQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_C6 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_D1 = CLBLM_R_X5Y136_SLICE_X7Y136_C5Q;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_D2 = CLBLL_L_X4Y134_SLICE_X4Y134_BQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_D4 = CLBLM_L_X10Y136_SLICE_X12Y136_CQ;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_D5 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_R_X3Y136_SLICE_X3Y136_D6 = 1'b1;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_D = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_A1 = CLBLM_R_X3Y138_SLICE_X3Y138_BO5;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_A2 = CLBLM_R_X3Y136_SLICE_X3Y136_D5Q;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_A3 = CLBLM_R_X3Y136_SLICE_X2Y136_AQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_A4 = CLBLM_R_X3Y139_SLICE_X3Y139_BQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_A6 = 1'b1;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_D = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_B1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_B2 = CLBLM_R_X3Y136_SLICE_X2Y136_BQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_B4 = CLBLL_L_X4Y136_SLICE_X4Y136_A5Q;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_B5 = CLBLL_L_X4Y139_SLICE_X4Y139_CQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_B6 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_C1 = CLBLL_L_X4Y135_SLICE_X4Y135_AQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_C2 = CLBLM_R_X3Y136_SLICE_X2Y136_CQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_C4 = CLBLL_L_X4Y130_SLICE_X4Y130_BQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_C5 = CLBLM_R_X3Y136_SLICE_X3Y136_DQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_C6 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_D1 = CLBLM_R_X3Y132_SLICE_X2Y132_AQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_D3 = CLBLM_R_X3Y136_SLICE_X2Y136_DQ;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_D4 = 1'b1;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_D5 = CLBLL_L_X4Y137_SLICE_X5Y137_B5Q;
  assign CLBLM_R_X3Y136_SLICE_X2Y136_D6 = CLBLM_R_X13Y134_SLICE_X18Y134_AO6;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A1 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A2 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A4 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A5 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A6 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_A3 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B1 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B2 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B3 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B4 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B5 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_B6 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C1 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C2 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C3 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C4 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C5 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_C6 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D1 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D2 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D3 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D4 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D5 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X17Y131_D6 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A1 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A2 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A3 = CLBLM_L_X8Y134_SLICE_X10Y134_A5Q;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A4 = CLBLL_L_X4Y136_SLICE_X5Y136_D5Q;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A5 = CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_A6 = CLBLM_R_X7Y137_SLICE_X8Y137_CQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B1 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B2 = CLBLL_L_X4Y136_SLICE_X5Y136_D5Q;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B3 = CLBLM_L_X8Y134_SLICE_X10Y134_A5Q;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B4 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B5 = CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_B6 = CLBLM_R_X7Y137_SLICE_X8Y137_CQ;
  assign RIOB33_X105Y157_IOB_X1Y157_O = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C1 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C2 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C3 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C4 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C5 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_C6 = 1'b1;
  assign RIOB33_X105Y157_IOB_X1Y158_O = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D1 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D2 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D3 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D4 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D5 = 1'b1;
  assign CLBLM_L_X12Y131_SLICE_X16Y131_D6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C2 = 1'b1;
  assign LIOB33_X0Y189_IOB_X0Y190_O = CLBLM_R_X7Y143_SLICE_X8Y143_BO5;
  assign LIOB33_X0Y189_IOB_X0Y189_O = CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C3 = CLBLM_R_X7Y134_SLICE_X8Y134_DO6;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A1 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A2 = CLBLM_R_X3Y136_SLICE_X2Y136_CQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A4 = CLBLM_R_X3Y135_SLICE_X3Y135_CQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A5 = CLBLM_L_X12Y136_SLICE_X16Y136_AQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_A6 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B2 = CLBLM_R_X5Y134_SLICE_X6Y134_AQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B3 = CLBLM_R_X3Y136_SLICE_X2Y136_AQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B5 = CLBLM_R_X3Y137_SLICE_X2Y137_AQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_B6 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C1 = CLBLL_L_X4Y134_SLICE_X4Y134_C5Q;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C2 = CLBLM_R_X3Y137_SLICE_X3Y137_CQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C3 = CLBLL_L_X4Y139_SLICE_X4Y139_BQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C5 = CLBLM_R_X5Y138_SLICE_X6Y138_B5Q;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_C6 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D2 = CLBLM_R_X3Y139_SLICE_X3Y139_A5Q;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D3 = CLBLM_R_X3Y137_SLICE_X3Y137_DQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D4 = CLBLM_L_X10Y140_SLICE_X13Y140_BQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D5 = CLBLM_R_X7Y139_SLICE_X8Y139_AQ;
  assign CLBLM_R_X3Y137_SLICE_X3Y137_D6 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D2 = CLBLM_R_X5Y134_SLICE_X6Y134_DQ;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_D1 = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D1 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A1 = CLBLL_L_X4Y135_SLICE_X5Y135_CQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A2 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A3 = CLBLM_R_X3Y137_SLICE_X2Y137_AQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A4 = CLBLM_R_X3Y137_SLICE_X3Y137_BQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A5 = CLBLM_R_X3Y137_SLICE_X3Y137_A5Q;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D3 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B1 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B2 = CLBLL_L_X2Y133_SLICE_X1Y133_AO6;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B3 = CLBLL_L_X2Y138_SLICE_X1Y138_AO6;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B4 = CLBLM_R_X3Y139_SLICE_X3Y139_BQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_B6 = CLBLM_R_X3Y137_SLICE_X2Y137_CO6;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D5 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C2 = CLBLM_R_X5Y137_SLICE_X7Y137_A5Q;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C4 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C5 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_C6 = CLBLM_R_X3Y138_SLICE_X2Y138_AQ;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D1 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D2 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D3 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D4 = CLBLM_R_X3Y136_SLICE_X3Y136_B5Q;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D5 = 1'b1;
  assign CLBLM_R_X3Y137_SLICE_X2Y137_D6 = CLBLM_R_X3Y137_SLICE_X3Y137_BQ;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A1 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A2 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A3 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A4 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A5 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_A6 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_T1 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B1 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B2 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B3 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B4 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B5 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_B6 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C1 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C2 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C3 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C4 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C5 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_C6 = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D1 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D2 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D3 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D4 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D5 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X17Y132_D6 = 1'b1;
  assign RIOB33_X105Y159_IOB_X1Y159_O = 1'b1;
  assign RIOB33_X105Y159_IOB_X1Y160_O = 1'b1;
  assign CLBLM_R_X7Y140_SLICE_X9Y140_D6 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A1 = CLBLM_R_X11Y140_SLICE_X14Y140_BO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A2 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A3 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A4 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A5 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_A6 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B1 = CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B2 = CLBLL_L_X4Y136_SLICE_X5Y136_D5Q;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B3 = CLBLM_L_X8Y134_SLICE_X10Y134_A5Q;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B4 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B5 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_B6 = CLBLM_R_X7Y137_SLICE_X8Y137_CQ;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C1 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C2 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C3 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C4 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C5 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_C6 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D1 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D2 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D3 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D4 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D5 = 1'b1;
  assign CLBLM_L_X12Y132_SLICE_X16Y132_D6 = 1'b1;
  assign LIOB33_X0Y191_IOB_X0Y191_O = CLBLM_R_X3Y133_SLICE_X3Y133_CO6;
  assign LIOB33_X0Y191_IOB_X0Y192_O = CLBLM_R_X3Y141_SLICE_X2Y141_AO5;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_D1 = RIOB33_X105Y125_IOB_X1Y125_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_T1 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_D1 = CLBLM_R_X5Y130_SLICE_X7Y130_CQ;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_D1 = RIOB33_X105Y123_IOB_X1Y124_I;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_T1 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_D1 = CLBLM_R_X7Y140_SLICE_X9Y140_D5Q;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_T1 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_D1 = CLBLM_L_X10Y130_SLICE_X12Y130_B5Q;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_T1 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_T1 = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_D1 = CLBLM_R_X3Y141_SLICE_X3Y141_AO5;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1 = CLBLM_R_X7Y136_SLICE_X8Y136_D5Q;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A2 = CLBLM_L_X10Y141_SLICE_X13Y141_BQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A3 = CLBLM_R_X3Y138_SLICE_X3Y138_AQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A4 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A5 = CLBLM_R_X3Y138_SLICE_X3Y138_A5Q;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_A6 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B1 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B2 = CLBLL_L_X4Y138_SLICE_X5Y138_AQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B3 = CLBLM_R_X3Y138_SLICE_X3Y138_AQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B4 = CLBLM_R_X3Y138_SLICE_X2Y138_BQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B5 = CLBLM_R_X3Y138_SLICE_X3Y138_A5Q;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_B6 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C1 = CLBLL_L_X4Y138_SLICE_X5Y138_AQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C2 = CLBLM_R_X3Y138_SLICE_X3Y138_AQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C3 = CLBLM_R_X3Y136_SLICE_X2Y136_AQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C4 = CLBLM_R_X3Y138_SLICE_X3Y138_A5Q;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C5 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_C6 = CLBLM_R_X3Y138_SLICE_X2Y138_BQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D1 = CLBLL_L_X4Y138_SLICE_X5Y138_AQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D2 = CLBLM_R_X3Y138_SLICE_X3Y138_AQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D3 = CLBLM_R_X3Y136_SLICE_X2Y136_AQ;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D4 = CLBLM_R_X3Y138_SLICE_X3Y138_A5Q;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D5 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_R_X3Y138_SLICE_X3Y138_D6 = CLBLM_R_X3Y138_SLICE_X2Y138_BQ;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A1 = CLBLM_R_X3Y141_SLICE_X2Y141_CO6;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A4 = CLBLM_R_X7Y135_SLICE_X9Y135_C5Q;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_A6 = CLBLM_R_X5Y137_SLICE_X7Y137_A5Q;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B1 = CLBLL_L_X4Y137_SLICE_X4Y137_CQ;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B2 = CLBLM_R_X3Y138_SLICE_X2Y138_BQ;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B3 = CLBLM_R_X3Y136_SLICE_X2Y136_AQ;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B5 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_B6 = CLBLM_R_X3Y138_SLICE_X3Y138_BO6;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C1 = CLBLM_R_X3Y141_SLICE_X2Y141_AQ;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C2 = CLBLM_R_X3Y138_SLICE_X2Y138_CQ;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C3 = 1'b1;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C4 = CLBLM_R_X13Y134_SLICE_X18Y134_AO6;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_C6 = CLBLM_R_X3Y133_SLICE_X2Y133_BQ;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D1 = CLBLM_R_X5Y137_SLICE_X7Y137_DO6;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D2 = CLBLM_R_X3Y137_SLICE_X3Y137_CQ;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D3 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D5 = CLBLM_R_X5Y138_SLICE_X6Y138_B5Q;
  assign CLBLM_R_X3Y138_SLICE_X2Y138_D6 = CLBLM_R_X3Y141_SLICE_X2Y141_AQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A1 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A2 = CLBLL_L_X4Y136_SLICE_X5Y136_D5Q;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A3 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A4 = CLBLM_L_X8Y134_SLICE_X10Y134_A5Q;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A5 = CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_A6 = CLBLM_R_X7Y137_SLICE_X8Y137_CQ;
  assign RIOB33_X105Y161_IOB_X1Y161_O = CLBLM_R_X3Y141_SLICE_X3Y141_AO5;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B1 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B2 = CLBLM_L_X8Y134_SLICE_X10Y134_A5Q;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B3 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B4 = CLBLL_L_X4Y136_SLICE_X5Y136_D5Q;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B5 = CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_B6 = CLBLM_R_X7Y137_SLICE_X8Y137_CQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C1 = CLBLM_R_X7Y132_SLICE_X9Y132_D5Q;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C2 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C3 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C4 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C5 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_C6 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D1 = CLBLM_L_X10Y132_SLICE_X12Y132_BQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D2 = CLBLM_R_X11Y133_SLICE_X14Y133_BQ;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D3 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D4 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D5 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X12Y133_SLICE_X17Y133_D6 = CLBLM_L_X12Y133_SLICE_X17Y133_BO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A1 = CLBLM_L_X12Y134_SLICE_X16Y134_CO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A2 = CLBLM_L_X12Y133_SLICE_X17Y133_DO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A3 = CLBLM_L_X8Y136_SLICE_X11Y136_CO5;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A4 = CLBLM_L_X12Y133_SLICE_X16Y133_BO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A5 = CLBLM_R_X3Y133_SLICE_X3Y133_BQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_A6 = CLBLM_L_X12Y133_SLICE_X16Y133_CO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C4 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C5 = 1'b1;
  assign LIOB33_X0Y193_IOB_X0Y193_O = CLBLL_L_X4Y142_SLICE_X4Y142_BO6;
  assign LIOB33_X0Y193_IOB_X0Y194_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B1 = CLBLM_R_X11Y133_SLICE_X15Y133_CO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B2 = CLBLM_R_X5Y133_SLICE_X6Y133_CO5;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B3 = CLBLM_L_X12Y133_SLICE_X17Y133_AO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B4 = CLBLM_L_X12Y135_SLICE_X17Y135_BO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B5 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_B6 = CLBLM_R_X13Y134_SLICE_X18Y134_DO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C6 = 1'b1;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_D = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C1 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C2 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C3 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C4 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C5 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_C6 = CLBLM_R_X5Y137_SLICE_X7Y137_AQ;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_D = LIOB33_X0Y55_IOB_X0Y55_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_D = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_D = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D1 = CLBLM_R_X3Y133_SLICE_X3Y133_BQ;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D2 = CLBLM_R_X3Y133_SLICE_X3Y133_B5Q;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D3 = CLBLM_L_X12Y133_SLICE_X17Y133_DO6;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D4 = 1'b1;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D5 = CLBLM_L_X8Y136_SLICE_X11Y136_CO5;
  assign CLBLM_L_X12Y133_SLICE_X16Y133_D6 = CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D5 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D6 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A4 = CLBLM_L_X10Y139_SLICE_X13Y139_A5Q;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A5 = CLBLM_R_X5Y143_SLICE_X7Y143_AQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D4 = CLBLM_L_X12Y139_SLICE_X17Y139_AO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A1 = CLBLM_R_X3Y139_SLICE_X2Y139_C5Q;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A2 = CLBLM_L_X10Y136_SLICE_X12Y136_CQ;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A4 = CLBLL_L_X4Y137_SLICE_X4Y137_AQ;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A5 = CLBLM_R_X5Y140_SLICE_X6Y140_CQ;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_A6 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B1 = CLBLM_R_X3Y138_SLICE_X2Y138_DO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B2 = CLBLM_R_X3Y137_SLICE_X2Y137_BO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B3 = CLBLL_L_X4Y139_SLICE_X4Y139_BQ;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B4 = CLBLM_R_X3Y139_SLICE_X2Y139_BQ;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B5 = CLBLM_R_X3Y139_SLICE_X2Y139_AQ;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_B6 = CLBLL_L_X4Y141_SLICE_X5Y141_CO6;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1 = CLBLL_L_X4Y141_SLICE_X5Y141_BO5;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_BX = CLBLM_R_X3Y141_SLICE_X3Y141_AO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C1 = CLBLM_R_X3Y139_SLICE_X2Y139_AQ;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C2 = CLBLL_L_X4Y139_SLICE_X4Y139_BQ;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C4 = CLBLL_L_X4Y141_SLICE_X5Y141_CO6;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C5 = CLBLM_R_X3Y135_SLICE_X2Y135_AQ;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_C6 = CLBLM_R_X3Y139_SLICE_X2Y139_BQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D5 = CLBLM_R_X5Y130_SLICE_X7Y130_DQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B4 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B5 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D1 = CLBLM_R_X3Y137_SLICE_X3Y137_D5Q;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D2 = CLBLM_L_X8Y141_SLICE_X11Y141_BQ;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D3 = CLBLM_R_X3Y136_SLICE_X3Y136_C5Q;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D4 = CLBLM_R_X3Y139_SLICE_X3Y139_A5Q;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D5 = CLBLM_R_X3Y139_SLICE_X2Y139_C5Q;
  assign CLBLM_R_X3Y139_SLICE_X3Y139_D6 = CLBLL_L_X4Y134_SLICE_X5Y134_DQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B6 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A2 = CLBLL_L_X2Y134_SLICE_X1Y134_AO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A3 = CLBLM_R_X3Y139_SLICE_X2Y139_AQ;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A4 = CLBLM_R_X3Y139_SLICE_X3Y139_CO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A5 = CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_A6 = CLBLM_R_X5Y136_SLICE_X6Y136_BQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D6 = CLBLM_L_X8Y143_SLICE_X10Y143_BO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B1 = CLBLL_L_X4Y135_SLICE_X5Y135_CQ;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B2 = CLBLM_R_X3Y139_SLICE_X2Y139_BQ;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B3 = CLBLM_R_X3Y139_SLICE_X2Y139_AQ;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B4 = CLBLM_R_X3Y139_SLICE_X3Y139_CO6;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_B6 = CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  assign RIOB33_X105Y163_IOB_X1Y163_O = CLBLM_R_X7Y136_SLICE_X8Y136_D5Q;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C1 = CLBLM_L_X8Y141_SLICE_X11Y141_BQ;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C2 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C3 = CLBLL_L_X4Y133_SLICE_X5Y133_CQ;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C4 = CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_C6 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C3 = 1'b1;
  assign RIOB33_X105Y163_IOB_X1Y164_O = CLBLM_L_X10Y141_SLICE_X12Y141_BQ;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C4 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C5 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D1 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D2 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D3 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D4 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D5 = 1'b1;
  assign CLBLM_R_X3Y139_SLICE_X2Y139_D6 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C6 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A1 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A2 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A3 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A4 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A5 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_A6 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B1 = CLBLM_R_X11Y131_SLICE_X14Y131_DO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B2 = CLBLM_L_X12Y134_SLICE_X16Y134_DO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B3 = CLBLM_R_X11Y140_SLICE_X14Y140_BO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B4 = CLBLM_L_X12Y135_SLICE_X16Y135_DO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B5 = CLBLM_L_X12Y134_SLICE_X17Y134_CO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_B6 = CLBLM_L_X12Y133_SLICE_X17Y133_CO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C1 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C2 = CLBLM_R_X3Y134_SLICE_X2Y134_AQ;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C3 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C4 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C5 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_C6 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign LIOB33_X0Y195_IOB_X0Y195_O = CLBLL_L_X4Y140_SLICE_X4Y140_DO6;
  assign LIOB33_X0Y195_IOB_X0Y196_O = CLBLL_L_X4Y143_SLICE_X4Y143_AO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D5 = CLBLM_L_X12Y135_SLICE_X17Y135_DO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D1 = CLBLM_R_X11Y132_SLICE_X15Y132_CO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D6 = CLBLM_L_X10Y132_SLICE_X13Y132_BO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D2 = CLBLM_R_X13Y134_SLICE_X18Y134_BO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D3 = CLBLM_L_X12Y133_SLICE_X16Y133_DO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D4 = CLBLM_L_X12Y133_SLICE_X17Y133_AO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D6 = CLBLM_L_X12Y134_SLICE_X17Y134_BO6;
  assign CLBLM_L_X12Y134_SLICE_X17Y134_D5 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1 = CLBLM_R_X7Y143_SLICE_X8Y143_BO5;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A1 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A2 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A3 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A4 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A5 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_A6 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_D1 = CLBLL_L_X4Y132_SLICE_X5Y132_A5Q;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B1 = CLBLM_R_X11Y131_SLICE_X14Y131_DO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B2 = CLBLM_L_X12Y135_SLICE_X16Y135_DO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B3 = CLBLM_R_X11Y133_SLICE_X14Y133_AQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B4 = CLBLM_R_X7Y132_SLICE_X9Y132_D5Q;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B5 = CLBLM_L_X12Y134_SLICE_X16Y134_AO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_B6 = CLBLM_R_X11Y136_SLICE_X15Y136_AO5;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D3 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D4 = 1'b1;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C1 = CLBLM_R_X11Y136_SLICE_X15Y136_AO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C2 = CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C3 = CLBLM_R_X3Y134_SLICE_X2Y134_AQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C4 = CLBLM_R_X3Y133_SLICE_X3Y133_B5Q;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C5 = CLBLM_R_X11Y140_SLICE_X14Y140_BO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_C6 = CLBLM_L_X12Y134_SLICE_X16Y134_BO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D1 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D2 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D3 = CLBLM_R_X11Y133_SLICE_X14Y133_AQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D4 = CLBLM_L_X12Y140_SLICE_X16Y140_AO5;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D5 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_L_X12Y134_SLICE_X16Y134_D6 = CLBLM_R_X5Y137_SLICE_X7Y137_AQ;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1 = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_T1 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B2 = CLBLM_L_X10Y136_SLICE_X12Y136_BQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B3 = CLBLM_L_X10Y136_SLICE_X12Y136_AQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B4 = CLBLL_L_X4Y135_SLICE_X5Y135_CQ;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_D1 = CLBLL_L_X4Y131_SLICE_X4Y131_D5Q;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_A1 = CLBLM_R_X3Y135_SLICE_X3Y135_AQ;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_A2 = CLBLL_L_X4Y140_SLICE_X4Y140_AO5;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_A3 = CLBLM_R_X3Y140_SLICE_X3Y140_AQ;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_A5 = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_A6 = CLBLM_R_X5Y142_SLICE_X6Y142_B5Q;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_T1 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_B1 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_B2 = CLBLM_R_X3Y135_SLICE_X2Y135_AQ;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_B3 = CLBLM_R_X3Y138_SLICE_X3Y138_AQ;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_B4 = CLBLM_R_X5Y133_SLICE_X7Y133_A5Q;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_B6 = CLBLM_R_X7Y136_SLICE_X8Y136_AQ;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_C2 = CLBLM_L_X10Y140_SLICE_X13Y140_BQ;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_C3 = CLBLM_L_X8Y142_SLICE_X11Y142_AQ;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_C4 = CLBLM_R_X3Y140_SLICE_X3Y140_BQ;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_C5 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_C6 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_D2 = CLBLM_R_X5Y130_SLICE_X7Y130_CQ;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_D3 = CLBLM_R_X3Y140_SLICE_X3Y140_DQ;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_D4 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_D5 = CLBLM_R_X5Y141_SLICE_X7Y141_AO6;
  assign CLBLM_R_X3Y140_SLICE_X3Y140_D6 = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_D1 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign RIOB33_X105Y165_IOB_X1Y165_O = CLBLM_R_X11Y142_SLICE_X15Y142_AO6;
  assign RIOB33_X105Y165_IOB_X1Y166_O = CLBLM_L_X10Y140_SLICE_X12Y140_AQ;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_A1 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_A2 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_A3 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_A4 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_A5 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_A6 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = CLBLL_L_X4Y136_SLICE_X4Y136_CQ;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_T1 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_B1 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_B2 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_B3 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_B4 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_B5 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_B6 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_D1 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_D1 = CLBLM_L_X10Y140_SLICE_X12Y140_AQ;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_C1 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_C2 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_C3 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_C4 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_C5 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_C6 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = CLBLM_R_X7Y135_SLICE_X9Y135_C5Q;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_T1 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_T1 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_D1 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_D2 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_D3 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_D4 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_D5 = 1'b1;
  assign CLBLM_R_X3Y140_SLICE_X2Y140_D6 = 1'b1;
  assign LIOB33_X0Y197_IOB_X0Y197_O = CLBLM_R_X3Y141_SLICE_X2Y141_BO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A1 = CLBLL_L_X4Y136_SLICE_X5Y136_D5Q;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A2 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A3 = CLBLM_R_X7Y137_SLICE_X8Y137_CQ;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A4 = CLBLM_L_X8Y134_SLICE_X10Y134_A5Q;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A5 = CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_A6 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C4 = CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B1 = CLBLM_R_X13Y138_SLICE_X18Y138_BO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B2 = CLBLM_L_X12Y135_SLICE_X17Y135_CO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B3 = CLBLM_R_X13Y134_SLICE_X18Y134_AO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B4 = CLBLM_L_X12Y136_SLICE_X17Y136_BO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B5 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_B6 = CLBLM_L_X12Y135_SLICE_X17Y135_AO5;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_T1 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C1 = CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C2 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C3 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C4 = CLBLM_R_X7Y137_SLICE_X8Y137_CQ;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C5 = CLBLL_L_X4Y136_SLICE_X5Y136_D5Q;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_C6 = CLBLM_L_X8Y134_SLICE_X10Y134_A5Q;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C5 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D1 = CLBLM_L_X12Y131_SLICE_X16Y131_AO6;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D2 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D3 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D4 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D5 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X12Y135_SLICE_X17Y135_D6 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A1 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A2 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A3 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A4 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A5 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_A6 = 1'b1;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B1 = CLBLM_L_X8Y136_SLICE_X11Y136_CO5;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B2 = CLBLM_R_X3Y140_SLICE_X3Y140_C5Q;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B3 = CLBLM_L_X10Y135_SLICE_X13Y135_AO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B4 = CLBLM_L_X10Y134_SLICE_X13Y134_DO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B5 = CLBLM_L_X12Y135_SLICE_X16Y135_AO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_B6 = CLBLM_L_X8Y137_SLICE_X10Y137_BQ;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_C6 = CLBLM_R_X5Y137_SLICE_X6Y137_DO5;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C1 = CLBLM_R_X11Y132_SLICE_X15Y132_AO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C2 = CLBLM_L_X8Y135_SLICE_X10Y135_CQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C3 = CLBLM_R_X11Y131_SLICE_X15Y131_AO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C4 = CLBLM_R_X5Y132_SLICE_X7Y132_CQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C5 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_C6 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D1 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D2 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D3 = CLBLL_L_X4Y142_SLICE_X4Y142_A5Q;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D4 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D5 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X12Y135_SLICE_X16Y135_D6 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_D1 = RIOB33_X105Y121_IOB_X1Y122_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_D = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_D = LIOB33_X0Y59_IOB_X0Y59_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_D = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_D = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B5 = CLBLM_R_X3Y135_SLICE_X3Y135_AQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A4 = CLBLL_L_X2Y138_SLICE_X1Y138_AO5;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A5 = CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_A6 = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_T1 = 1'b1;
  assign RIOB33_X105Y167_IOB_X1Y167_O = CLBLM_L_X10Y137_SLICE_X13Y137_AQ;
  assign RIOB33_X105Y167_IOB_X1Y168_O = CLBLM_L_X8Y135_SLICE_X11Y135_AQ;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B1 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B2 = CLBLM_R_X3Y136_SLICE_X2Y136_B5Q;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B3 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B4 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B5 = CLBLL_L_X4Y130_SLICE_X4Y130_D5Q;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_B6 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B6 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C1 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C2 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C3 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C4 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C5 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_C6 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D1 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D2 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D3 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D4 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D5 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X3Y141_D6 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A2 = CLBLL_L_X2Y138_SLICE_X1Y138_AO5;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A3 = CLBLM_R_X3Y141_SLICE_X2Y141_AQ;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A4 = CLBLL_L_X4Y142_SLICE_X5Y142_BQ;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_A6 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_AX = CLBLM_R_X3Y141_SLICE_X2Y141_BO5;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B2 = CLBLL_L_X2Y138_SLICE_X1Y138_AO5;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B5 = CLBLL_L_X4Y135_SLICE_X4Y135_AQ;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_B6 = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_D1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_BX = CLBLM_R_X3Y141_SLICE_X2Y141_AO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C1 = CLBLM_R_X7Y140_SLICE_X9Y140_BQ;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C2 = CLBLM_R_X3Y141_SLICE_X2Y141_AQ;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C3 = CLBLM_R_X3Y135_SLICE_X2Y135_AQ;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C4 = CLBLL_L_X2Y138_SLICE_X1Y138_AO5;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_C6 = CLBLM_R_X7Y141_SLICE_X8Y141_BO6;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D1 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D2 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D3 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D4 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D5 = 1'b1;
  assign CLBLM_R_X3Y141_SLICE_X2Y141_D6 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_A1 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_A2 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_A3 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_A4 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_A5 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_A6 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_B1 = CLBLL_L_X4Y136_SLICE_X5Y136_D5Q;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_B2 = CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_B3 = CLBLM_L_X8Y134_SLICE_X10Y134_A5Q;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_B4 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_B5 = CLBLM_L_X12Y139_SLICE_X16Y139_AO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_B6 = CLBLM_R_X7Y137_SLICE_X8Y137_CQ;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_C1 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_C2 = CLBLM_L_X12Y136_SLICE_X16Y136_CO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_C3 = CLBLM_L_X10Y136_SLICE_X12Y136_DO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_C4 = CLBLM_L_X12Y135_SLICE_X17Y135_BO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_C5 = CLBLM_L_X12Y136_SLICE_X17Y136_DO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_C6 = CLBLM_L_X12Y133_SLICE_X17Y133_AO6;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_T1 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_D1 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_D2 = CLBLM_R_X13Y137_SLICE_X18Y137_AO5;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_D3 = CLBLM_R_X11Y136_SLICE_X14Y136_AQ;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_D4 = CLBLM_R_X13Y138_SLICE_X18Y138_BO6;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_D5 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_L_X12Y136_SLICE_X17Y136_D6 = CLBLM_L_X12Y136_SLICE_X17Y136_BO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_A2 = CLBLM_R_X7Y134_SLICE_X8Y134_CQ;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_A3 = CLBLM_L_X12Y136_SLICE_X17Y136_CO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_A4 = CLBLM_L_X12Y138_SLICE_X16Y138_BO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_A5 = CLBLM_R_X11Y133_SLICE_X14Y133_BQ;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_A6 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_B1 = CLBLM_L_X10Y131_SLICE_X13Y131_CO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_B2 = CLBLM_L_X12Y136_SLICE_X17Y136_BO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_B3 = CLBLM_L_X12Y136_SLICE_X16Y136_AQ;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_B4 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_B5 = CLBLM_L_X10Y136_SLICE_X12Y136_C5Q;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_B6 = CLBLM_R_X11Y134_SLICE_X14Y134_AO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_C1 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_C2 = CLBLM_L_X12Y135_SLICE_X16Y135_CO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_C3 = CLBLM_L_X12Y136_SLICE_X17Y136_BO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_C4 = CLBLM_L_X12Y136_SLICE_X16Y136_A5Q;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_C5 = CLBLM_R_X7Y136_SLICE_X8Y136_BQ;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_C6 = CLBLM_R_X11Y134_SLICE_X14Y134_AO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_D1 = CLBLM_L_X10Y136_SLICE_X12Y136_C5Q;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_D2 = CLBLM_L_X12Y136_SLICE_X16Y136_AQ;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_D3 = CLBLM_L_X12Y136_SLICE_X17Y136_BO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_D4 = CLBLM_R_X11Y134_SLICE_X14Y134_AO6;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_D5 = 1'b1;
  assign CLBLM_L_X12Y136_SLICE_X16Y136_D6 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign LIOB33_X0Y109_IOB_X0Y110_O = CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  assign RIOB33_X105Y169_IOB_X1Y170_O = CLBLM_R_X3Y140_SLICE_X3Y140_AQ;
  assign RIOB33_X105Y169_IOB_X1Y169_O = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign LIOB33_X0Y109_IOB_X0Y109_O = CLBLL_L_X4Y130_SLICE_X4Y130_BQ;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A1 = CLBLM_L_X8Y140_SLICE_X10Y140_CQ;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A2 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A3 = CLBLM_L_X12Y135_SLICE_X17Y135_CO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A4 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_A6 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B1 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B2 = CLBLM_R_X11Y140_SLICE_X14Y140_BO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B3 = CLBLM_L_X12Y131_SLICE_X16Y131_AO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B4 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B5 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_B6 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C1 = CLBLM_L_X12Y133_SLICE_X17Y133_AO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C2 = CLBLM_L_X12Y137_SLICE_X16Y137_CO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C3 = CLBLM_L_X12Y135_SLICE_X17Y135_BO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C5 = CLBLM_L_X12Y137_SLICE_X17Y137_DO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_C6 = CLBLM_L_X12Y140_SLICE_X16Y140_BO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D1 = CLBLM_L_X12Y137_SLICE_X17Y137_AO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D2 = CLBLM_L_X10Y136_SLICE_X13Y136_BQ;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D3 = CLBLM_R_X13Y137_SLICE_X18Y137_AO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D4 = CLBLM_L_X12Y139_SLICE_X17Y139_AO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D5 = CLBLM_R_X13Y134_SLICE_X18Y134_AO6;
  assign CLBLM_L_X12Y137_SLICE_X17Y137_D6 = CLBLM_L_X10Y137_SLICE_X12Y137_BQ;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A1 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A2 = CLBLM_R_X5Y129_SLICE_X7Y129_AQ;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A3 = CLBLM_R_X7Y139_SLICE_X8Y139_AQ;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A4 = CLBLM_L_X12Y136_SLICE_X17Y136_BO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A5 = CLBLM_L_X12Y135_SLICE_X17Y135_CO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_A6 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_D1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B1 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B2 = CLBLM_L_X12Y135_SLICE_X17Y135_BO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B3 = CLBLM_L_X12Y133_SLICE_X17Y133_AO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B4 = CLBLM_R_X11Y137_SLICE_X15Y137_AO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B5 = CLBLM_L_X12Y137_SLICE_X16Y137_AO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_B6 = CLBLM_L_X12Y140_SLICE_X16Y140_BO6;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_T1 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C1 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C2 = CLBLM_R_X3Y136_SLICE_X2Y136_DQ;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C3 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C4 = CLBLM_L_X12Y136_SLICE_X17Y136_BO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C5 = CLBLM_L_X12Y140_SLICE_X16Y140_AQ;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_C6 = CLBLM_L_X12Y135_SLICE_X17Y135_CO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_D1 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D1 = CLBLM_L_X12Y137_SLICE_X16Y137_AO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D2 = CLBLM_R_X13Y137_SLICE_X18Y137_DO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D3 = CLBLM_L_X12Y135_SLICE_X17Y135_BO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D4 = CLBLM_R_X11Y132_SLICE_X14Y132_CO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D5 = CLBLM_L_X12Y133_SLICE_X17Y133_AO6;
  assign CLBLM_L_X12Y137_SLICE_X16Y137_D6 = CLBLM_R_X11Y137_SLICE_X15Y137_AO6;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_D1 = CLBLM_L_X8Y135_SLICE_X11Y135_AQ;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_T1 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = CLBLM_R_X3Y132_SLICE_X3Y132_BQ;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_T1 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_D1 = CLBLM_L_X10Y137_SLICE_X13Y137_AQ;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_D1 = CLBLM_R_X5Y140_SLICE_X6Y140_A5Q;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1 = CLBLM_R_X5Y133_SLICE_X7Y133_CQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_D1 = CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1 = 1'b1;
  assign RIOB33_X105Y171_IOB_X1Y172_O = CLBLM_R_X3Y134_SLICE_X2Y134_AQ;
  assign RIOB33_X105Y171_IOB_X1Y171_O = CLBLM_R_X7Y141_SLICE_X9Y141_BO6;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_T1 = 1'b1;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_D = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_D = LIOB33_X0Y61_IOB_X0Y61_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_D = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_D = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_A1 = CLBLM_L_X12Y135_SLICE_X17Y135_AO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_A2 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_A3 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_A4 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_A5 = CLBLM_L_X12Y131_SLICE_X16Y131_AO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_A6 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_B1 = CLBLM_L_X12Y136_SLICE_X16Y136_DO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_B2 = CLBLM_L_X12Y133_SLICE_X17Y133_AO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_B3 = CLBLM_L_X12Y135_SLICE_X17Y135_BO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_B4 = CLBLM_L_X12Y138_SLICE_X17Y138_DO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_B5 = CLBLM_L_X10Y131_SLICE_X13Y131_CO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_B6 = CLBLM_L_X12Y139_SLICE_X17Y139_CO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_C1 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_C2 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_C3 = CLBLM_R_X11Y140_SLICE_X15Y140_AQ;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_C4 = CLBLM_L_X12Y136_SLICE_X17Y136_AO5;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_C5 = CLBLM_L_X12Y135_SLICE_X17Y135_AO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_C6 = CLBLM_R_X13Y138_SLICE_X18Y138_BO5;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_D1 = CLBLM_L_X12Y138_SLICE_X17Y138_CO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_D2 = 1'b1;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_D3 = CLBLM_R_X11Y138_SLICE_X14Y138_AQ;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_D4 = CLBLM_L_X10Y141_SLICE_X13Y141_BQ;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_D5 = CLBLM_R_X13Y137_SLICE_X18Y137_AO6;
  assign CLBLM_L_X12Y138_SLICE_X17Y138_D6 = CLBLM_L_X12Y137_SLICE_X17Y137_BO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_A1 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_A2 = CLBLM_L_X12Y135_SLICE_X17Y135_CO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_A3 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_A4 = RIOB33_X105Y137_IOB_X1Y138_I;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_A5 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_A6 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_D1 = CLBLM_R_X3Y141_SLICE_X2Y141_AO5;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_B1 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_B2 = CLBLM_L_X12Y136_SLICE_X16Y136_BO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_B3 = CLBLM_L_X12Y133_SLICE_X17Y133_AO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_B4 = CLBLM_R_X11Y138_SLICE_X14Y138_AO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_B5 = CLBLM_L_X10Y137_SLICE_X12Y137_BO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_B6 = CLBLM_L_X12Y138_SLICE_X16Y138_CO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C4 = CLBLM_L_X10Y131_SLICE_X12Y131_D5Q;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_D = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_C1 = CLBLM_L_X12Y135_SLICE_X17Y135_BO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_C2 = CLBLM_L_X12Y140_SLICE_X16Y140_DO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_C3 = CLBLM_L_X10Y141_SLICE_X13Y141_BQ;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_C4 = CLBLM_L_X12Y139_SLICE_X16Y139_AO5;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_C5 = CLBLM_L_X12Y138_SLICE_X16Y138_DO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_C6 = CLBLM_L_X12Y137_SLICE_X17Y137_BO6;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_T1 = 1'b1;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_D = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_D1 = CLBLM_R_X13Y137_SLICE_X18Y137_AO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_D2 = CLBLM_R_X13Y138_SLICE_X18Y138_BO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_D3 = CLBLM_R_X11Y140_SLICE_X15Y140_AQ;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_D4 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_D5 = CLBLM_R_X13Y138_SLICE_X18Y138_AO6;
  assign CLBLM_L_X12Y138_SLICE_X16Y138_D6 = CLBLM_R_X11Y138_SLICE_X14Y138_AQ;
  assign RIOB33_X105Y173_IOB_X1Y174_O = CLBLM_R_X5Y140_SLICE_X6Y140_BO5;
  assign RIOB33_X105Y173_IOB_X1Y173_O = CLBLM_R_X5Y140_SLICE_X6Y140_A5Q;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C5 = CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C6 = CLBLM_R_X11Y140_SLICE_X14Y140_BO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A1 = CLBLM_L_X12Y135_SLICE_X17Y135_AO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A2 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A3 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A4 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A5 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_A6 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_T1 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B1 = CLBLM_L_X12Y135_SLICE_X17Y135_AO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B2 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B3 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B4 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B5 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_B6 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C1 = CLBLM_L_X8Y140_SLICE_X11Y140_CQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D1 = CLBLM_R_X11Y133_SLICE_X14Y133_CO5;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C2 = CLBLM_L_X12Y139_SLICE_X16Y139_AO5;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C3 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C4 = CLBLM_L_X12Y136_SLICE_X17Y136_BO6;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C5 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D2 = CLBLM_L_X8Y137_SLICE_X11Y137_CQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_C6 = CLBLM_L_X12Y140_SLICE_X16Y140_BO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D3 = CLBLM_R_X3Y137_SLICE_X3Y137_DQ;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D1 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D2 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D3 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D4 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D5 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X17Y139_D6 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A1 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A2 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A3 = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A4 = CLBLM_R_X11Y140_SLICE_X14Y140_CQ;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A5 = CLBLM_L_X12Y135_SLICE_X17Y135_CO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_A6 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B2 = CLBLM_R_X13Y138_SLICE_X18Y138_BO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B3 = CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B4 = CLBLM_R_X13Y137_SLICE_X18Y137_BO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B5 = CLBLM_R_X13Y138_SLICE_X18Y138_AO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_B6 = RIOB33_X105Y139_IOB_X1Y140_I;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C1 = CLBLM_R_X13Y134_SLICE_X18Y134_AO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C2 = CLBLM_R_X3Y138_SLICE_X2Y138_CQ;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C3 = CLBLM_L_X12Y139_SLICE_X17Y139_BO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C4 = CLBLM_R_X13Y138_SLICE_X18Y138_AO5;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C5 = CLBLM_L_X12Y140_SLICE_X16Y140_BO5;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_C6 = CLBLM_L_X12Y136_SLICE_X17Y136_BO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A1 = CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D3 = CLBLM_R_X13Y138_SLICE_X18Y138_BO6;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D2 = 1'b1;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D4 = CLBLM_R_X3Y138_SLICE_X2Y138_CQ;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D5 = CLBLM_L_X12Y140_SLICE_X16Y140_BO5;
  assign CLBLM_L_X12Y139_SLICE_X16Y139_D6 = CLBLM_L_X12Y136_SLICE_X17Y136_BO6;
  assign RIOB33_X105Y175_IOB_X1Y176_O = CLBLM_R_X3Y138_SLICE_X3Y138_DO6;
  assign RIOB33_X105Y175_IOB_X1Y175_O = CLBLL_L_X4Y142_SLICE_X5Y142_CO5;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_D1 = RIOB33_X105Y119_IOB_X1Y120_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_T1 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_D1 = CLBLM_R_X5Y133_SLICE_X7Y133_AQ;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_D1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_T1 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_D1 = CLBLM_R_X3Y134_SLICE_X2Y134_AQ;
  assign LIOI3_X0Y65_OLOGIC_X0Y66_D1 = CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_T1 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_D1 = CLBLM_L_X8Y138_SLICE_X10Y138_CQ;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_T1 = 1'b1;
  assign LIOI3_X0Y65_OLOGIC_X0Y66_T1 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_T1 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_D1 = CLBLM_R_X7Y141_SLICE_X9Y141_BO6;
  assign LIOI3_X0Y65_OLOGIC_X0Y65_D1 = CLBLL_L_X2Y133_SLICE_X1Y133_BO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = CLBLM_R_X5Y138_SLICE_X7Y138_AQ;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_T1 = 1'b1;
  assign LIOI3_X0Y65_OLOGIC_X0Y65_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = CLBLM_R_X3Y132_SLICE_X3Y132_BQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_A1 = CLBLM_R_X13Y138_SLICE_X18Y138_CO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_A2 = CLBLM_R_X11Y140_SLICE_X15Y140_CO5;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_A3 = CLBLM_L_X12Y140_SLICE_X16Y140_CO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_A4 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_A5 = CLBLM_L_X12Y140_SLICE_X16Y140_AQ;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_A6 = CLBLM_R_X13Y137_SLICE_X18Y137_CO6;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_B1 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_B2 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_B3 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_B4 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_B5 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_B6 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A1 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A2 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A3 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A4 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A5 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_A6 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_C1 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_C2 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_C3 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B1 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B2 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B3 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B4 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B5 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_B6 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_D1 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_D2 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C1 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C2 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C3 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C4 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C5 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_C6 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_D3 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_D4 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_D5 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_D6 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_A1 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_A2 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_A3 = CLBLM_L_X12Y135_SLICE_X17Y135_CO6;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D1 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D2 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D3 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D4 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D5 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X13Y130_D6 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_A5 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_A6 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_B6 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_AX = CLBLM_R_X11Y140_SLICE_X14Y140_DQ;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_B1 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_B2 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A1 = CLBLM_R_X7Y135_SLICE_X9Y135_B5Q;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A2 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A3 = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A5 = CLBLM_L_X10Y130_SLICE_X12Y130_C5Q;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_C1 = CLBLM_R_X7Y139_SLICE_X8Y139_AQ;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_C2 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_C3 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B1 = CLBLM_L_X10Y135_SLICE_X12Y135_A5Q;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B2 = CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B3 = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B4 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_B6 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_D1 = CLBLM_L_X12Y135_SLICE_X17Y135_CO6;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C1 = CLBLM_R_X7Y135_SLICE_X9Y135_AQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C4 = CLBLM_L_X10Y138_SLICE_X12Y138_BQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C5 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_C6 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_D2 = CLBLM_L_X12Y136_SLICE_X17Y136_BO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_D3 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_D4 = CLBLM_L_X8Y140_SLICE_X11Y140_CQ;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_D6 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D1 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D2 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D3 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D4 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D5 = 1'b1;
  assign CLBLM_L_X10Y130_SLICE_X12Y130_D6 = 1'b1;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_D = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_D = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_A1 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_A2 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_A3 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_A4 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_A5 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_A6 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_B1 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_B2 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_B3 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_B4 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_B5 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_B6 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_C1 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_C2 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_C3 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_C4 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_C5 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_C6 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_D1 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_D2 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_D3 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_D4 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_D5 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X19Y134_D6 = 1'b1;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_A1 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_A2 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_A3 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_A4 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_A5 = CLBLM_L_X12Y131_SLICE_X16Y131_AO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_A6 = CLBLM_R_X11Y140_SLICE_X14Y140_BO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_B1 = CLBLM_R_X13Y137_SLICE_X18Y137_BO5;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_B2 = CLBLM_R_X7Y131_SLICE_X8Y131_DQ;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_B3 = CLBLM_R_X13Y138_SLICE_X18Y138_AO5;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_B4 = CLBLM_L_X12Y136_SLICE_X17Y136_BO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_B5 = CLBLM_R_X13Y134_SLICE_X18Y134_AO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_B6 = CLBLM_R_X13Y134_SLICE_X18Y134_CO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_C1 = LIOB33_X0Y51_IOB_X0Y51_I;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_C2 = CLBLM_L_X12Y135_SLICE_X17Y135_AO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_C3 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_C4 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_C5 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_C6 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_D1 = LIOB33_X0Y51_IOB_X0Y51_I;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_D2 = CLBLM_R_X13Y138_SLICE_X18Y138_BO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_D3 = CLBLM_R_X13Y137_SLICE_X18Y137_BO5;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_D4 = CLBLM_L_X12Y136_SLICE_X17Y136_BO6;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_D5 = CLBLM_R_X7Y131_SLICE_X8Y131_DQ;
  assign CLBLM_R_X13Y134_SLICE_X18Y134_D6 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_A1 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_A2 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_A3 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_A4 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_A5 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_A6 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_B1 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_B2 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_B3 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_B4 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_B5 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_B6 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A2 = CLBLM_L_X10Y131_SLICE_X13Y131_BQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A3 = CLBLM_L_X10Y131_SLICE_X13Y131_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A4 = CLBLM_L_X8Y131_SLICE_X11Y131_D5Q;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A5 = CLBLM_R_X5Y133_SLICE_X7Y133_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_A6 = CLBLL_L_X4Y135_SLICE_X4Y135_D5Q;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_C1 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_C2 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_C3 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B2 = CLBLM_L_X10Y132_SLICE_X13Y132_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B3 = CLBLL_L_X4Y135_SLICE_X5Y135_CQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B4 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B5 = CLBLM_L_X10Y131_SLICE_X13Y131_BQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_B6 = CLBLM_R_X7Y131_SLICE_X9Y131_DQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_D1 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_D2 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C1 = CLBLM_R_X11Y131_SLICE_X14Y131_AO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C2 = CLBLM_R_X11Y131_SLICE_X14Y131_AO5;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C3 = CLBLM_R_X11Y132_SLICE_X15Y132_BO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C4 = CLBLL_L_X4Y130_SLICE_X5Y130_B5Q;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C5 = CLBLM_R_X7Y134_SLICE_X8Y134_AQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_C6 = CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_D3 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X17Y141_D4 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_A1 = CLBLM_L_X12Y141_SLICE_X16Y141_BO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_A2 = CLBLM_R_X7Y135_SLICE_X9Y135_DQ;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_A3 = CLBLM_R_X11Y138_SLICE_X14Y138_AQ;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_A4 = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_A5 = CLBLM_L_X12Y140_SLICE_X17Y140_AO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D1 = CLBLM_R_X11Y131_SLICE_X14Y131_AO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D2 = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D3 = CLBLM_R_X11Y132_SLICE_X15Y132_BO6;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D4 = CLBLM_L_X8Y139_SLICE_X11Y139_C5Q;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D5 = CLBLM_R_X7Y131_SLICE_X8Y131_CQ;
  assign CLBLM_L_X10Y131_SLICE_X13Y131_D6 = CLBLM_R_X11Y131_SLICE_X14Y131_AO5;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_B1 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_B2 = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_B3 = CLBLM_R_X11Y140_SLICE_X14Y140_BQ;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_B4 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A2 = CLBLM_L_X8Y131_SLICE_X11Y131_BQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A3 = CLBLM_L_X10Y131_SLICE_X12Y131_AQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A4 = CLBLM_L_X10Y131_SLICE_X12Y131_CQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A5 = CLBLM_R_X7Y131_SLICE_X9Y131_D5Q;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_A6 = CLBLM_L_X10Y140_SLICE_X13Y140_D5Q;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_C1 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_C2 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_C3 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B1 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B2 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B3 = CLBLL_L_X4Y131_SLICE_X5Y131_AQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B5 = CLBLM_L_X10Y131_SLICE_X12Y131_C5Q;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_B6 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_D1 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_D2 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C1 = CLBLM_L_X10Y132_SLICE_X12Y132_C5Q;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C2 = CLBLM_L_X10Y131_SLICE_X12Y131_CQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C3 = CLBLM_R_X3Y135_SLICE_X3Y135_DQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C4 = CLBLM_R_X3Y137_SLICE_X3Y137_B5Q;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_C6 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_D3 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_D4 = 1'b1;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_D5 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y141_SLICE_X16Y141_D6 = 1'b1;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D1 = CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D4 = CLBLM_L_X8Y131_SLICE_X11Y131_D5Q;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D5 = CLBLL_L_X4Y136_SLICE_X4Y136_CQ;
  assign CLBLM_L_X10Y131_SLICE_X12Y131_D6 = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_D1 = CLBLM_R_X7Y143_SLICE_X8Y143_BO5;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_T1 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_D1 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_D1 = CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_T1 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_A1 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_A2 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_A3 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_A4 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_A5 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_A6 = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_T1 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_D1 = CLBLM_R_X5Y140_SLICE_X6Y140_BO5;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_B1 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_B2 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_B3 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_B4 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_B5 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_B6 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_D1 = CLBLM_L_X10Y140_SLICE_X13Y140_D5Q;
  assign RIOB33_X105Y181_IOB_X1Y181_O = CLBLM_R_X7Y143_SLICE_X8Y143_BO5;
  assign RIOB33_X105Y181_IOB_X1Y182_O = CLBLL_L_X4Y141_SLICE_X5Y141_BO5;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A2 = CLBLL_L_X4Y134_SLICE_X5Y134_BQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A3 = CLBLM_L_X10Y132_SLICE_X13Y132_AQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A5 = CLBLM_L_X12Y132_SLICE_X16Y132_AO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_A6 = CLBLL_L_X4Y134_SLICE_X4Y134_C5Q;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_C1 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_C2 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_C3 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B1 = CLBLM_L_X8Y132_SLICE_X10Y132_B5Q;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B2 = CLBLL_L_X4Y132_SLICE_X5Y132_DQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B3 = CLBLM_R_X11Y131_SLICE_X14Y131_AO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B4 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B5 = CLBLM_L_X12Y132_SLICE_X16Y132_BO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_B6 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_D1 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_D2 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C1 = CLBLM_L_X12Y132_SLICE_X16Y132_BO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C2 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C3 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C4 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C5 = CLBLM_L_X8Y134_SLICE_X10Y134_AQ;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_C6 = CLBLM_R_X11Y131_SLICE_X15Y131_AO6;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_D3 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X17Y142_D4 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_A1 = CLBLM_L_X12Y133_SLICE_X16Y133_AO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_A2 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_A3 = CLBLM_L_X10Y139_SLICE_X13Y139_A5Q;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_A4 = CLBLM_R_X11Y135_SLICE_X15Y135_BO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_A5 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D1 = CLBLM_R_X11Y131_SLICE_X15Y131_AO6;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D2 = CLBLM_L_X8Y139_SLICE_X11Y139_C5Q;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D3 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D4 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D5 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X13Y132_D6 = CLBLM_R_X7Y131_SLICE_X8Y131_CQ;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_A6 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_B5 = CLBLM_L_X10Y139_SLICE_X13Y139_A5Q;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_B6 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_B1 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_B2 = CLBLM_L_X12Y138_SLICE_X16Y138_BO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_B3 = CLBLM_R_X11Y135_SLICE_X14Y135_AO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_B4 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A2 = CLBLM_L_X10Y132_SLICE_X12Y132_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A3 = CLBLM_L_X8Y132_SLICE_X11Y132_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A4 = CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A5 = CLBLM_L_X10Y131_SLICE_X12Y131_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_A6 = CLBLM_L_X8Y135_SLICE_X11Y135_BO6;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_C1 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_C2 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_C3 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B2 = CLBLM_L_X10Y132_SLICE_X12Y132_BQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B3 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B4 = CLBLM_R_X5Y130_SLICE_X7Y130_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B5 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_B6 = CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_D1 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_D2 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_D3 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C1 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C2 = CLBLM_R_X3Y135_SLICE_X2Y135_AQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C4 = CLBLM_L_X10Y131_SLICE_X12Y131_DQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C5 = CLBLM_L_X8Y131_SLICE_X11Y131_C5Q;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_C6 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_D4 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_D5 = 1'b1;
  assign CLBLM_L_X12Y142_SLICE_X16Y142_D6 = 1'b1;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D1 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D2 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D3 = CLBLM_R_X7Y132_SLICE_X9Y132_CQ;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D4 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D5 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X10Y132_SLICE_X12Y132_D6 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_D = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_D = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOB33_X105Y183_IOB_X1Y184_O = CLBLL_L_X4Y143_SLICE_X4Y143_AO6;
  assign RIOB33_X105Y183_IOB_X1Y183_O = 1'b0;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A1 = CLBLM_R_X3Y135_SLICE_X3Y135_CQ;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A3 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A4 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A5 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_A6 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A1 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B1 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B2 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B3 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B4 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B5 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_B6 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A2 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A3 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_A4 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C1 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C2 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C3 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C4 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C5 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_C6 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_B1 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A1 = CLBLM_R_X5Y133_SLICE_X7Y133_AQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A2 = CLBLM_R_X7Y133_SLICE_X8Y133_A5Q;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A3 = CLBLM_L_X10Y133_SLICE_X13Y133_AQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A5 = CLBLL_L_X4Y135_SLICE_X4Y135_D5Q;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D1 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D2 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D3 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D4 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D5 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X4Y129_D6 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_A6 = CLBLM_L_X8Y133_SLICE_X11Y133_B5Q;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B1 = CLBLM_L_X12Y136_SLICE_X17Y136_BO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B2 = CLBLM_R_X7Y133_SLICE_X9Y133_DQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B3 = CLBLM_R_X11Y132_SLICE_X15Y132_BO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B4 = CLBLM_L_X10Y132_SLICE_X13Y132_CO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B5 = CLBLM_R_X11Y141_SLICE_X14Y141_AQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_B6 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C1 = CLBLL_L_X4Y131_SLICE_X5Y131_B5Q;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C2 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C3 = CLBLM_R_X5Y134_SLICE_X6Y134_B5Q;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C4 = CLBLM_L_X12Y136_SLICE_X17Y136_BO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C5 = CLBLM_R_X11Y132_SLICE_X15Y132_BO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_C6 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X17Y143_D4 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A1 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A2 = CLBLM_L_X10Y139_SLICE_X13Y139_A5Q;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A3 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A4 = CLBLM_R_X11Y139_SLICE_X15Y139_BO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_A5 = CLBLM_L_X12Y136_SLICE_X17Y136_CO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D1 = CLBLM_R_X11Y131_SLICE_X14Y131_AO6;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D2 = CLBLM_R_X7Y137_SLICE_X8Y137_B5Q;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D3 = CLBLL_L_X4Y134_SLICE_X4Y134_A5Q;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D4 = CLBLM_L_X10Y133_SLICE_X13Y133_CO6;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B1 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B2 = 1'b1;
  assign CLBLM_L_X12Y143_SLICE_X16Y143_B3 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D5 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X13Y133_D6 = CLBLM_R_X11Y134_SLICE_X14Y134_AO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A1 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A2 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A3 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A4 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A5 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_A6 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A2 = CLBLM_L_X8Y133_SLICE_X10Y133_CQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A3 = CLBLM_R_X3Y131_SLICE_X2Y131_BQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_A5 = CLBLM_R_X11Y141_SLICE_X14Y141_AQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B1 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B5 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B6 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B2 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C1 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C2 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C3 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C4 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C5 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_C6 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B2 = CLBLM_L_X10Y133_SLICE_X12Y133_BQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B3 = CLBLM_L_X10Y131_SLICE_X13Y131_BQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B5 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_B6 = CLBLM_L_X8Y134_SLICE_X11Y134_B5Q;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C1 = CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D1 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D2 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D3 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D4 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D5 = 1'b1;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_D6 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_C5 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D1 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D2 = CLBLM_R_X7Y135_SLICE_X8Y135_AQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D3 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D5 = 1'b1;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D6 = CLBLM_L_X10Y130_SLICE_X12Y130_BQ;
  assign CLBLM_L_X10Y133_SLICE_X12Y133_D4 = CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_A1 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_A2 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_A3 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_A4 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_A5 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_A6 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_B1 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_B2 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_B3 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_B4 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_B5 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_B6 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_C1 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_C2 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_C3 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_C4 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_C5 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_C6 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_D1 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_D2 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_D3 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_D4 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_D5 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X19Y137_D6 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_A1 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_A2 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_A3 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_A4 = CLBLM_L_X12Y135_SLICE_X17Y135_CO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_A5 = CLBLM_R_X11Y136_SLICE_X15Y136_AQ;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_A6 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_B1 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_B2 = CLBLM_L_X12Y135_SLICE_X17Y135_CO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_B3 = CLBLM_L_X8Y136_SLICE_X10Y136_AQ;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_B4 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_B5 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_B6 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_C1 = CLBLM_R_X11Y136_SLICE_X15Y136_AQ;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_C2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_C3 = CLBLM_L_X10Y137_SLICE_X12Y137_BQ;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_C4 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_C5 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_C6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_D1 = CLBLM_R_X11Y142_SLICE_X15Y142_AO5;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_D1 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_D2 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_D3 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_D4 = CLBLM_L_X12Y135_SLICE_X17Y135_CO6;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_D5 = 1'b1;
  assign CLBLM_R_X13Y137_SLICE_X18Y137_D6 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign RIOB33_X105Y185_IOB_X1Y186_O = CLBLM_R_X7Y141_SLICE_X8Y141_DO6;
  assign RIOB33_X105Y185_IOB_X1Y185_O = CLBLM_R_X7Y141_SLICE_X8Y141_CO6;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_T1 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A1 = CLBLM_R_X5Y130_SLICE_X6Y130_CO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A2 = CLBLM_R_X5Y130_SLICE_X6Y130_B5Q;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A3 = CLBLL_L_X4Y130_SLICE_X4Y130_AQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A5 = CLBLM_R_X5Y129_SLICE_X6Y129_AQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_A6 = CLBLM_R_X7Y131_SLICE_X8Y131_C5Q;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B1 = CLBLM_R_X5Y133_SLICE_X7Y133_BQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B3 = CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B4 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B5 = CLBLL_L_X4Y138_SLICE_X4Y138_AQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_B6 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C1 = CLBLM_R_X5Y129_SLICE_X6Y129_AQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C2 = CLBLL_L_X4Y130_SLICE_X4Y130_AQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C3 = CLBLM_R_X5Y130_SLICE_X6Y130_CO6;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C4 = CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_C6 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A1 = CLBLM_L_X10Y136_SLICE_X13Y136_AQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D1 = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D2 = CLBLL_L_X4Y130_SLICE_X5Y130_A5Q;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D3 = CLBLM_R_X5Y133_SLICE_X7Y133_CQ;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D4 = CLBLM_R_X5Y133_SLICE_X7Y133_A5Q;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y130_SLICE_X4Y130_D6 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A2 = CLBLM_L_X8Y136_SLICE_X11Y136_BQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A3 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B1 = CLBLM_R_X7Y139_SLICE_X9Y139_AQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A5 = CLBLM_L_X10Y140_SLICE_X13Y140_B5Q;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_A6 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B2 = CLBLM_R_X11Y136_SLICE_X14Y136_CO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B3 = CLBLM_L_X8Y133_SLICE_X10Y133_AQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B4 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B5 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C1 = CLBLM_R_X5Y131_SLICE_X6Y131_AQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_B6 = CLBLM_R_X11Y140_SLICE_X14Y140_BO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C2 = CLBLM_L_X12Y134_SLICE_X16Y134_AO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C3 = CLBLL_L_X4Y136_SLICE_X5Y136_DQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C4 = CLBLM_R_X11Y136_SLICE_X15Y136_AO5;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C5 = CLBLM_L_X12Y134_SLICE_X16Y134_AO5;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_C6 = CLBLM_L_X8Y136_SLICE_X11Y136_BQ;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D1 = CLBLM_L_X10Y139_SLICE_X13Y139_AQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A1 = CLBLL_L_X4Y130_SLICE_X5Y130_DO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A2 = CLBLM_R_X3Y137_SLICE_X3Y137_D5Q;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A3 = CLBLL_L_X4Y130_SLICE_X5Y130_AQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A4 = CLBLM_R_X5Y130_SLICE_X6Y130_B5Q;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_A6 = CLBLL_L_X4Y130_SLICE_X5Y130_CO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D2 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D3 = CLBLM_L_X10Y133_SLICE_X12Y133_DO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_AX = CLBLL_L_X4Y130_SLICE_X4Y130_CO6;
  assign CLBLM_L_X10Y134_SLICE_X13Y134_D4 = CLBLM_R_X11Y136_SLICE_X15Y136_AO5;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B1 = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B2 = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B3 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B5 = CLBLL_L_X4Y141_SLICE_X4Y141_DQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_B6 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A6 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_A5 = CLBLM_L_X8Y135_SLICE_X10Y135_C5Q;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C1 = CLBLM_R_X5Y130_SLICE_X7Y130_BQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C2 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B1 = CLBLL_L_X4Y137_SLICE_X5Y137_A5Q;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B2 = CLBLM_R_X11Y141_SLICE_X14Y141_AQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B3 = CLBLM_L_X8Y134_SLICE_X11Y134_AQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C3 = CLBLL_L_X4Y134_SLICE_X4Y134_CQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C4 = CLBLM_R_X7Y131_SLICE_X8Y131_A5Q;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C5 = CLBLM_R_X3Y131_SLICE_X3Y131_AQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_C6 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B5 = CLBLM_L_X10Y139_SLICE_X13Y139_AQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_B6 = 1'b1;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D1 = CLBLL_L_X4Y130_SLICE_X4Y130_AQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D2 = CLBLL_L_X4Y130_SLICE_X5Y130_AQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D3 = CLBLM_R_X5Y129_SLICE_X6Y129_AQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D4 = CLBLM_R_X5Y130_SLICE_X6Y130_CO6;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D5 = CLBLL_L_X4Y131_SLICE_X4Y131_BQ;
  assign CLBLL_L_X4Y130_SLICE_X5Y130_D6 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C1 = CLBLM_R_X11Y133_SLICE_X15Y133_AO6;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C2 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C3 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C4 = CLBLM_L_X10Y135_SLICE_X13Y135_AQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C5 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_C6 = CLBLM_R_X7Y133_SLICE_X9Y133_AQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D1 = CLBLM_L_X10Y132_SLICE_X12Y132_AQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D2 = CLBLM_L_X10Y134_SLICE_X13Y134_A5Q;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D3 = CLBLM_L_X10Y134_SLICE_X12Y134_BQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D5 = 1'b1;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D6 = CLBLM_L_X8Y132_SLICE_X11Y132_BQ;
  assign CLBLM_L_X10Y134_SLICE_X12Y134_D4 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_T1 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_D1 = CLBLM_R_X3Y133_SLICE_X3Y133_CO6;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_D1 = CLBLM_R_X3Y138_SLICE_X3Y138_DO6;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_D1 = CLBLM_R_X3Y132_SLICE_X3Y132_BQ;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_D1 = CLBLL_L_X4Y142_SLICE_X5Y142_CO5;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_A1 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_A2 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_A3 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_A4 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_A5 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1 = CLBLM_R_X7Y139_SLICE_X8Y139_AO6;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_T1 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_B1 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_B2 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_B3 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_B4 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_B5 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1 = CLBLL_L_X4Y141_SLICE_X5Y141_BO5;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_C1 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_C2 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_C3 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_C4 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_C5 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1 = CLBLL_L_X4Y138_SLICE_X4Y138_AO5;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_D1 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_D2 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_D3 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_D4 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_D5 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X19Y138_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1 = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_A1 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_A2 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_A3 = CLBLM_L_X12Y135_SLICE_X17Y135_AO6;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_A4 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_A5 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_A6 = 1'b1;
  assign LIOB33_X0Y101_IOB_X0Y101_O = CLBLM_R_X3Y136_SLICE_X2Y136_BQ;
  assign LIOB33_X0Y101_IOB_X0Y102_O = CLBLM_R_X5Y129_SLICE_X7Y129_BQ;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_B1 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_B2 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_B3 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_B4 = CLBLM_L_X12Y135_SLICE_X17Y135_AO6;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_B5 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_B6 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_C1 = CLBLM_L_X8Y136_SLICE_X10Y136_AQ;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_C2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_C3 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_C4 = RIOB33_X105Y137_IOB_X1Y138_I;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_C5 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_C6 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_D1 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_D2 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_D3 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_D4 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_D5 = 1'b1;
  assign CLBLM_R_X13Y138_SLICE_X18Y138_D6 = 1'b1;
  assign RIOB33_X105Y187_IOB_X1Y187_O = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign RIOB33_X105Y187_IOB_X1Y188_O = CLBLL_L_X4Y141_SLICE_X5Y141_BO5;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A1 = CLBLM_R_X5Y141_SLICE_X6Y141_CQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A3 = CLBLL_L_X4Y131_SLICE_X4Y131_AQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A4 = CLBLM_R_X3Y132_SLICE_X3Y132_D5Q;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A5 = CLBLM_R_X5Y133_SLICE_X7Y133_AQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_A6 = CLBLL_L_X4Y135_SLICE_X4Y135_D5Q;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B1 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B2 = CLBLL_L_X4Y131_SLICE_X4Y131_BQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B3 = CLBLM_R_X5Y130_SLICE_X6Y130_B5Q;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B4 = CLBLL_L_X4Y132_SLICE_X4Y132_BQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B5 = CLBLL_L_X4Y130_SLICE_X4Y130_CO5;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C2 = CLBLL_L_X4Y131_SLICE_X4Y131_CQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C3 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C4 = CLBLM_R_X3Y131_SLICE_X3Y131_B5Q;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C5 = CLBLL_L_X4Y135_SLICE_X5Y135_CQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_C6 = CLBLM_R_X5Y130_SLICE_X7Y130_D5Q;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D2 = CLBLL_L_X4Y132_SLICE_X5Y132_A5Q;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D3 = CLBLL_L_X4Y131_SLICE_X4Y131_DQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D4 = CLBLM_R_X3Y132_SLICE_X3Y132_D5Q;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D5 = CLBLM_R_X3Y135_SLICE_X3Y135_DQ;
  assign CLBLL_L_X4Y131_SLICE_X4Y131_D6 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A1 = CLBLM_R_X7Y137_SLICE_X9Y137_BQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A2 = CLBLM_R_X11Y140_SLICE_X14Y140_BO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A3 = CLBLM_L_X8Y133_SLICE_X11Y133_CO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A4 = CLBLM_L_X10Y138_SLICE_X13Y138_CQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A5 = CLBLM_R_X11Y133_SLICE_X14Y133_CO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_A6 = CLBLM_L_X12Y136_SLICE_X17Y136_AO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_AX = CLBLM_L_X10Y136_SLICE_X13Y136_CO5;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B1 = CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B2 = CLBLM_L_X10Y137_SLICE_X12Y137_AQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B3 = CLBLM_R_X7Y139_SLICE_X9Y139_BQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B4 = CLBLM_L_X10Y135_SLICE_X12Y135_CO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B5 = CLBLM_R_X11Y136_SLICE_X15Y136_AO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_B6 = CLBLM_L_X12Y136_SLICE_X17Y136_AO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C1 = CLBLM_L_X12Y134_SLICE_X16Y134_AO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C2 = CLBLM_R_X5Y135_SLICE_X7Y135_AQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C3 = CLBLM_R_X5Y136_SLICE_X6Y136_CQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C4 = CLBLM_L_X12Y136_SLICE_X17Y136_AO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C5 = CLBLM_R_X3Y134_SLICE_X3Y134_A5Q;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_C6 = CLBLM_R_X11Y136_SLICE_X15Y136_AO5;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A1 = CLBLM_R_X7Y135_SLICE_X9Y135_C5Q;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A2 = CLBLL_L_X4Y133_SLICE_X5Y133_D5Q;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A3 = CLBLL_L_X4Y131_SLICE_X5Y131_AQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D1 = CLBLM_L_X8Y140_SLICE_X11Y140_AQ;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D2 = CLBLM_R_X5Y135_SLICE_X7Y135_B5Q;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D3 = CLBLM_R_X11Y131_SLICE_X14Y131_BO6;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D4 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D5 = CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  assign CLBLM_L_X10Y135_SLICE_X13Y135_D6 = CLBLM_R_X11Y140_SLICE_X14Y140_BO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A5 = CLBLL_L_X4Y131_SLICE_X5Y131_BQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_A6 = CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B1 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B3 = CLBLM_R_X11Y135_SLICE_X14Y135_AO6;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B4 = CLBLL_L_X4Y131_SLICE_X4Y131_BQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B5 = CLBLM_R_X5Y138_SLICE_X7Y138_AQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_B6 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A4 = CLBLM_L_X8Y135_SLICE_X10Y135_D5Q;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_A6 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C1 = CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C2 = CLBLM_R_X3Y137_SLICE_X3Y137_C5Q;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C3 = CLBLL_L_X4Y130_SLICE_X4Y130_AQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C4 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C5 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B1 = CLBLM_R_X7Y135_SLICE_X8Y135_AQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B2 = CLBLM_L_X12Y136_SLICE_X16Y136_A5Q;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B4 = CLBLM_R_X7Y140_SLICE_X8Y140_D5Q;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B5 = 1'b1;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_B6 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_C6 = CLBLM_R_X3Y131_SLICE_X3Y131_AQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D1 = CLBLM_L_X8Y134_SLICE_X10Y134_AQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C1 = CLBLM_L_X12Y132_SLICE_X16Y132_AO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C2 = CLBLM_R_X3Y135_SLICE_X2Y135_CQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C3 = CLBLM_L_X12Y135_SLICE_X16Y135_AO5;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C4 = CLBLM_L_X10Y132_SLICE_X12Y132_CQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C5 = CLBLM_L_X10Y135_SLICE_X12Y135_DO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_C6 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D2 = 1'b1;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D3 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D4 = CLBLM_L_X8Y139_SLICE_X11Y139_C5Q;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y131_SLICE_X5Y131_D6 = CLBLL_L_X4Y131_SLICE_X4Y131_BQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D1 = CLBLM_R_X7Y139_SLICE_X9Y139_BQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D2 = CLBLM_R_X11Y136_SLICE_X14Y136_CO6;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D3 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D4 = CLBLM_L_X10Y137_SLICE_X12Y137_AQ;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D5 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X10Y135_SLICE_X12Y135_D6 = CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  assign LIOB33_X0Y141_IOB_X0Y142_O = CLBLM_R_X3Y132_SLICE_X3Y132_BQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C4 = CLBLM_R_X5Y136_SLICE_X7Y136_CQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C6 = CLBLM_L_X8Y136_SLICE_X10Y136_AO6;
  assign LIOB33_X0Y103_IOB_X0Y104_O = CLBLM_R_X5Y130_SLICE_X7Y130_D5Q;
  assign LIOB33_X0Y103_IOB_X0Y103_O = CLBLM_L_X10Y134_SLICE_X12Y134_B5Q;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_D = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOB33_X105Y189_IOB_X1Y190_O = CLBLM_R_X11Y142_SLICE_X15Y142_AO5;
  assign RIOB33_X105Y189_IOB_X1Y189_O = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D2 = CLBLM_R_X5Y131_SLICE_X7Y131_AQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D5 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D6 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A1 = CLBLL_L_X4Y132_SLICE_X4Y132_CQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A2 = CLBLL_L_X4Y136_SLICE_X5Y136_D5Q;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A3 = CLBLL_L_X4Y132_SLICE_X4Y132_AQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A5 = CLBLL_L_X4Y132_SLICE_X4Y132_BQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_A6 = CLBLL_L_X4Y133_SLICE_X4Y133_AQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B1 = CLBLL_L_X4Y132_SLICE_X4Y132_CQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B2 = CLBLL_L_X4Y132_SLICE_X4Y132_BQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B3 = CLBLL_L_X4Y132_SLICE_X4Y132_AQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B5 = CLBLL_L_X4Y133_SLICE_X4Y133_C5Q;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_B6 = CLBLL_L_X4Y133_SLICE_X4Y133_AQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B2 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B3 = CLBLM_L_X8Y138_SLICE_X11Y138_AQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C1 = CLBLL_L_X4Y132_SLICE_X4Y132_BQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C2 = CLBLL_L_X4Y132_SLICE_X4Y132_CQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C3 = CLBLL_L_X4Y132_SLICE_X4Y132_AQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C5 = CLBLM_R_X3Y132_SLICE_X3Y132_CQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_C6 = CLBLL_L_X4Y133_SLICE_X4Y133_AQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D1 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D2 = CLBLM_L_X8Y132_SLICE_X11Y132_CO6;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D3 = CLBLL_L_X4Y132_SLICE_X4Y132_DQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D5 = CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  assign CLBLL_L_X4Y132_SLICE_X4Y132_D6 = CLBLM_R_X5Y133_SLICE_X6Y133_BQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A2 = CLBLM_R_X7Y140_SLICE_X8Y140_AQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A3 = CLBLM_L_X10Y136_SLICE_X13Y136_AQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A4 = CLBLM_L_X10Y137_SLICE_X13Y137_AQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A5 = CLBLM_L_X12Y132_SLICE_X16Y132_AO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_A6 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B2 = CLBLM_L_X10Y136_SLICE_X13Y136_BQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B3 = CLBLM_R_X11Y133_SLICE_X14Y133_AQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B4 = CLBLM_L_X8Y138_SLICE_X11Y138_CQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B5 = CLBLL_L_X4Y135_SLICE_X5Y135_CQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_B6 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C1 = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C1 = CLBLM_L_X12Y136_SLICE_X16Y136_AQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C2 = CLBLM_L_X10Y140_SLICE_X13Y140_B5Q;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C3 = CLBLM_R_X11Y142_SLICE_X14Y142_AQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C4 = CLBLL_L_X4Y131_SLICE_X5Y131_B5Q;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_C6 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A1 = CLBLL_L_X4Y136_SLICE_X5Y136_CQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A2 = CLBLL_L_X4Y130_SLICE_X4Y130_DQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A3 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A5 = CLBLM_L_X10Y140_SLICE_X13Y140_B5Q;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_A6 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D1 = CLBLM_R_X11Y136_SLICE_X14Y136_BO6;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B1 = CLBLL_L_X4Y136_SLICE_X5Y136_CQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B2 = CLBLL_L_X4Y132_SLICE_X5Y132_BQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B3 = CLBLM_R_X5Y141_SLICE_X6Y141_CQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B4 = CLBLL_L_X4Y131_SLICE_X5Y131_BQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_B6 = CLBLM_R_X5Y134_SLICE_X7Y134_BQ;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D2 = CLBLM_L_X10Y140_SLICE_X13Y140_B5Q;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D3 = CLBLM_R_X11Y134_SLICE_X14Y134_AO6;
  assign CLBLM_L_X10Y136_SLICE_X13Y136_D4 = CLBLM_R_X5Y136_SLICE_X6Y136_BQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C2 = CLBLM_R_X5Y128_SLICE_X6Y128_DO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A1 = CLBLM_L_X10Y140_SLICE_X13Y140_CQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A2 = CLBLL_L_X4Y135_SLICE_X5Y135_CQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C3 = CLBLM_R_X7Y140_SLICE_X9Y140_BQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C4 = CLBLM_R_X5Y134_SLICE_X7Y134_DQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C5 = CLBLL_L_X4Y132_SLICE_X5Y132_CQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_C6 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A3 = CLBLM_L_X10Y136_SLICE_X12Y136_AQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A4 = CLBLM_L_X8Y133_SLICE_X10Y133_CQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_A6 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D2 = CLBLL_L_X4Y133_SLICE_X4Y133_AQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D3 = CLBLM_L_X10Y140_SLICE_X13Y140_B5Q;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D4 = 1'b1;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D5 = CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  assign CLBLL_L_X4Y132_SLICE_X5Y132_D6 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B1 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C2 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_B6 = CLBLM_R_X7Y136_SLICE_X9Y136_DQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C3 = CLBLM_L_X10Y131_SLICE_X13Y131_AQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C4 = CLBLM_L_X12Y136_SLICE_X16Y136_AQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C5 = CLBLM_R_X5Y132_SLICE_X7Y132_CQ;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_C6 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C5 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C6 = 1'b1;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D1 = CLBLM_L_X10Y139_SLICE_X12Y139_CO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D2 = CLBLM_L_X10Y132_SLICE_X12Y132_DO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D3 = CLBLM_L_X8Y136_SLICE_X11Y136_DO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D4 = CLBLM_L_X10Y137_SLICE_X12Y137_AO5;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D5 = CLBLM_L_X10Y139_SLICE_X12Y139_DO6;
  assign CLBLM_L_X10Y136_SLICE_X12Y136_D6 = CLBLM_L_X8Y136_SLICE_X10Y136_BO6;
  assign LIOB33_X0Y105_IOB_X0Y106_O = CLBLL_L_X4Y132_SLICE_X5Y132_BQ;
  assign LIOB33_X0Y105_IOB_X0Y105_O = CLBLL_L_X4Y137_SLICE_X5Y137_B5Q;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D4 = CLBLM_R_X7Y132_SLICE_X9Y132_A5Q;
  assign RIOB33_X105Y191_IOB_X1Y192_O = CLBLM_L_X12Y142_SLICE_X16Y142_AO6;
  assign RIOB33_X105Y191_IOB_X1Y191_O = CLBLM_L_X12Y142_SLICE_X16Y142_BO5;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_D1 = CLBLL_L_X4Y143_SLICE_X4Y143_AO6;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_T1 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_D1 = CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_D1 = CLBLL_L_X4Y140_SLICE_X4Y140_DO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_T1 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_D1 = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_T1 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_D1 = CLBLL_L_X4Y133_SLICE_X4Y133_BO5;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_T1 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_T1 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_D1 = CLBLM_L_X8Y140_SLICE_X11Y140_BQ;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A1 = CLBLM_R_X5Y140_SLICE_X7Y140_B5Q;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A2 = CLBLM_R_X5Y133_SLICE_X6Y133_BQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A3 = CLBLL_L_X4Y134_SLICE_X4Y134_CQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A4 = CLBLM_R_X3Y133_SLICE_X2Y133_AQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1 = CLBLM_R_X3Y140_SLICE_X3Y140_AQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B1 = CLBLM_R_X5Y134_SLICE_X6Y134_C5Q;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B2 = CLBLL_L_X4Y133_SLICE_X4Y133_BQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B3 = CLBLM_R_X5Y135_SLICE_X7Y135_B5Q;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B4 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C2 = CLBLL_L_X4Y132_SLICE_X5Y132_D5Q;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C3 = CLBLM_R_X3Y137_SLICE_X3Y137_DQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C4 = CLBLL_L_X4Y132_SLICE_X4Y132_DQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C5 = CLBLM_R_X7Y138_SLICE_X9Y138_B5Q;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_C6 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D1 = CLBLM_R_X5Y132_SLICE_X7Y132_AQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D2 = CLBLM_R_X5Y137_SLICE_X7Y137_BQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D3 = CLBLL_L_X4Y133_SLICE_X4Y133_DQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D5 = CLBLL_L_X4Y130_SLICE_X4Y130_DQ;
  assign CLBLL_L_X4Y133_SLICE_X4Y133_D6 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A1 = CLBLM_R_X7Y133_SLICE_X8Y133_D5Q;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A3 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A4 = CLBLM_L_X10Y132_SLICE_X12Y132_CQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A5 = CLBLM_R_X7Y137_SLICE_X8Y137_DQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_A6 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B1 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B2 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B3 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B4 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B5 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_B6 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C1 = CLBLM_R_X11Y133_SLICE_X14Y133_CO6;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C2 = CLBLM_L_X10Y137_SLICE_X12Y137_CO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A2 = CLBLM_L_X10Y140_SLICE_X13Y140_D5Q;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A3 = CLBLL_L_X4Y133_SLICE_X5Y133_AQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A4 = CLBLM_R_X5Y132_SLICE_X7Y132_BQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A5 = CLBLL_L_X4Y133_SLICE_X5Y133_C5Q;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_A6 = CLBLM_R_X7Y131_SLICE_X9Y131_D5Q;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C3 = CLBLM_L_X10Y138_SLICE_X13Y138_DQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_C4 = CLBLM_R_X11Y136_SLICE_X15Y136_AO5;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B1 = CLBLM_R_X7Y131_SLICE_X8Y131_DQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B2 = CLBLM_R_X5Y130_SLICE_X7Y130_CQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B4 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B5 = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_B6 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D4 = CLBLM_L_X10Y140_SLICE_X12Y140_DQ;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D5 = CLBLM_L_X10Y137_SLICE_X13Y137_BO5;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C1 = CLBLM_L_X8Y134_SLICE_X10Y134_AQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C2 = 1'b1;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C3 = CLBLM_R_X3Y136_SLICE_X3Y136_AQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C5 = CLBLM_R_X5Y132_SLICE_X6Y132_AQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_C6 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X13Y137_D6 = CLBLM_L_X10Y137_SLICE_X13Y137_BO6;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A2 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A4 = CLBLM_R_X11Y140_SLICE_X14Y140_BO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A5 = CLBLM_L_X8Y136_SLICE_X10Y136_BQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A6 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_A3 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D1 = CLBLL_L_X4Y133_SLICE_X4Y133_D5Q;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_AX = CLBLM_R_X3Y137_SLICE_X3Y137_C5Q;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D2 = CLBLM_R_X7Y140_SLICE_X8Y140_D5Q;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B1 = CLBLM_R_X7Y135_SLICE_X8Y135_CO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B2 = CLBLM_L_X10Y137_SLICE_X13Y137_BO5;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B3 = CLBLM_L_X10Y136_SLICE_X12Y136_CQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B4 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B5 = CLBLM_L_X8Y136_SLICE_X11Y136_CO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_B6 = CLBLM_R_X7Y137_SLICE_X8Y137_AQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D3 = CLBLM_R_X5Y134_SLICE_X6Y134_C5Q;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D4 = CLBLM_R_X5Y132_SLICE_X6Y132_AQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_BX = CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  assign CLBLL_L_X4Y133_SLICE_X5Y133_D6 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C1 = CLBLM_L_X8Y135_SLICE_X10Y135_B5Q;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C2 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C3 = CLBLL_L_X4Y137_SLICE_X4Y137_C5Q;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C4 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C5 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_C6 = CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y107_IOB_X0Y108_O = CLBLM_R_X5Y130_SLICE_X6Y130_BQ;
  assign LIOB33_X0Y107_IOB_X0Y107_O = CLBLM_R_X5Y133_SLICE_X7Y133_CQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D1 = CLBLM_L_X8Y136_SLICE_X11Y136_CO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D2 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D3 = CLBLM_L_X10Y137_SLICE_X13Y137_BO5;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D4 = CLBLM_L_X10Y136_SLICE_X12Y136_CQ;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D5 = 1'b1;
  assign CLBLM_L_X10Y137_SLICE_X12Y137_D6 = CLBLM_R_X7Y137_SLICE_X8Y137_AQ;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_D = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_D = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOB33_X105Y193_IOB_X1Y194_O = CLBLM_L_X12Y142_SLICE_X16Y142_BO6;
  assign RIOB33_X105Y193_IOB_X1Y193_O = CLBLM_R_X11Y142_SLICE_X14Y142_AO6;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A1 = CLBLM_L_X8Y134_SLICE_X10Y134_A5Q;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A2 = CLBLM_R_X7Y137_SLICE_X8Y137_CQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A3 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A4 = CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A5 = CLBLL_L_X4Y136_SLICE_X5Y136_D5Q;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_A6 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B1 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B2 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B3 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B4 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B5 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_B6 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C1 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C2 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C3 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C4 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C5 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_C6 = 1'b1;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D1 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D2 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D3 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D4 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D5 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X15Y131_D6 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A1 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A2 = CLBLM_L_X12Y131_SLICE_X16Y131_AO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A3 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A4 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A5 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_A6 = 1'b1;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B1 = CLBLM_R_X11Y140_SLICE_X14Y140_BO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B2 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B3 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B4 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B5 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_B6 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C1 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C2 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C3 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C4 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C5 = CLBLM_R_X11Y140_SLICE_X14Y140_BO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_C6 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1 = CLBLM_R_X3Y136_SLICE_X2Y136_A5Q;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D1 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D2 = CLBLM_L_X10Y132_SLICE_X13Y132_AQ;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D3 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D4 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_A5 = CLBLM_R_X3Y141_SLICE_X2Y141_CO6;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D5 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_R_X11Y131_SLICE_X14Y131_D6 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_A6 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A1 = CLBLM_R_X7Y131_SLICE_X9Y131_D5Q;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A3 = CLBLL_L_X4Y134_SLICE_X4Y134_AQ;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A4 = CLBLL_L_X4Y137_SLICE_X5Y137_D5Q;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A5 = CLBLM_L_X10Y140_SLICE_X13Y140_D5Q;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_A6 = CLBLM_R_X5Y134_SLICE_X7Y134_D5Q;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_AX = CLBLL_L_X4Y140_SLICE_X4Y140_AO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B1 = CLBLM_R_X3Y135_SLICE_X3Y135_DQ;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B2 = CLBLL_L_X4Y134_SLICE_X4Y134_BQ;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B4 = CLBLM_L_X8Y138_SLICE_X10Y138_CQ;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B5 = CLBLL_L_X4Y133_SLICE_X5Y133_D5Q;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_B6 = CLBLL_L_X4Y136_SLICE_X4Y136_D5Q;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_B2 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C1 = CLBLM_L_X12Y133_SLICE_X16Y133_AO6;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C2 = CLBLL_L_X4Y134_SLICE_X4Y134_D5Q;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C3 = CLBLM_R_X5Y140_SLICE_X7Y140_B5Q;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C5 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_C6 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_B5 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_B6 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D1 = CLBLL_L_X4Y129_SLICE_X4Y129_AQ;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D2 = CLBLM_R_X7Y136_SLICE_X8Y136_AQ;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D3 = CLBLM_R_X3Y135_SLICE_X2Y135_AQ;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D5 = CLBLM_R_X3Y136_SLICE_X3Y136_B5Q;
  assign CLBLL_L_X4Y134_SLICE_X4Y134_D6 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A1 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A2 = CLBLM_L_X10Y134_SLICE_X12Y134_BQ;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A3 = CLBLM_L_X10Y138_SLICE_X13Y138_AQ;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A5 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_A6 = CLBLL_L_X4Y133_SLICE_X5Y133_AQ;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B2 = CLBLM_L_X12Y136_SLICE_X16Y136_A5Q;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B3 = CLBLM_R_X11Y137_SLICE_X14Y137_DO6;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B4 = CLBLM_R_X11Y140_SLICE_X15Y140_B5Q;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_B6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A1 = CLBLL_L_X4Y135_SLICE_X5Y135_BQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A2 = CLBLM_R_X5Y135_SLICE_X6Y135_BQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A3 = CLBLL_L_X4Y134_SLICE_X5Y134_AQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A4 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C1 = CLBLL_L_X4Y135_SLICE_X4Y135_D5Q;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C2 = CLBLM_L_X10Y138_SLICE_X13Y138_CQ;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C3 = CLBLM_R_X5Y133_SLICE_X7Y133_AQ;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C4 = CLBLM_R_X7Y138_SLICE_X9Y138_BQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_C6 = CLBLM_L_X8Y133_SLICE_X10Y133_BQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_A6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B1 = CLBLM_L_X8Y138_SLICE_X10Y138_CQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B2 = CLBLL_L_X4Y134_SLICE_X5Y134_BQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B3 = CLBLL_L_X4Y136_SLICE_X4Y136_D5Q;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B4 = CLBLM_R_X5Y135_SLICE_X6Y135_BQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_B6 = CLBLM_R_X5Y134_SLICE_X6Y134_BQ;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C1 = CLBLM_R_X5Y134_SLICE_X7Y134_BQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C2 = CLBLL_L_X4Y134_SLICE_X5Y134_CQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C3 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D5 = CLBLM_R_X5Y133_SLICE_X7Y133_AQ;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D6 = CLBLL_L_X4Y135_SLICE_X4Y135_D5Q;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C4 = CLBLL_L_X4Y139_SLICE_X5Y139_CQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_C6 = CLBLM_R_X3Y139_SLICE_X2Y139_BQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D3 = CLBLM_L_X10Y138_SLICE_X13Y138_DQ;
  assign CLBLM_L_X10Y138_SLICE_X13Y138_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A1 = CLBLM_L_X12Y132_SLICE_X16Y132_AO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A3 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A4 = CLBLM_L_X8Y140_SLICE_X10Y140_BQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A6 = 1'b1;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_A5 = CLBLM_L_X8Y133_SLICE_X10Y133_BQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D2 = CLBLM_R_X5Y134_SLICE_X6Y134_BQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D3 = CLBLM_R_X5Y138_SLICE_X6Y138_B5Q;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D4 = CLBLM_R_X3Y137_SLICE_X3Y137_D5Q;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D5 = CLBLM_R_X7Y140_SLICE_X9Y140_DQ;
  assign CLBLL_L_X4Y134_SLICE_X5Y134_D6 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B1 = CLBLM_R_X13Y134_SLICE_X18Y134_AO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B2 = CLBLM_L_X10Y138_SLICE_X12Y138_BQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B4 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B5 = CLBLM_R_X3Y137_SLICE_X2Y137_AQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_B6 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C1 = CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C2 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C3 = CLBLM_L_X10Y138_SLICE_X12Y138_AQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C4 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C5 = CLBLM_R_X7Y133_SLICE_X8Y133_D5Q;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_C6 = CLBLM_R_X11Y136_SLICE_X14Y136_CO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D1 = CLBLM_L_X12Y132_SLICE_X16Y132_AO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D2 = 1'b1;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D3 = CLBLM_R_X11Y136_SLICE_X15Y136_AO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D4 = CLBLM_L_X10Y138_SLICE_X12Y138_CO6;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D5 = CLBLL_L_X4Y138_SLICE_X4Y138_BQ;
  assign CLBLM_L_X10Y138_SLICE_X12Y138_D6 = CLBLM_L_X8Y140_SLICE_X10Y140_BQ;
  assign RIOB33_X105Y195_IOB_X1Y195_O = CLBLM_L_X12Y143_SLICE_X16Y143_AO6;
  assign RIOB33_X105Y195_IOB_X1Y196_O = CLBLM_L_X12Y142_SLICE_X16Y142_AO5;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A1 = CLBLL_L_X4Y136_SLICE_X5Y136_D5Q;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A2 = CLBLM_R_X7Y137_SLICE_X8Y137_CQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A3 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A4 = CLBLM_L_X8Y134_SLICE_X10Y134_A5Q;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A5 = CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_A6 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B1 = CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B2 = CLBLM_L_X12Y140_SLICE_X16Y140_AO5;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B3 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B4 = CLBLM_L_X8Y134_SLICE_X10Y134_A5Q;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B5 = CLBLM_R_X7Y137_SLICE_X8Y137_CQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_B6 = CLBLL_L_X4Y136_SLICE_X5Y136_D5Q;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C1 = CLBLM_R_X11Y134_SLICE_X14Y134_AO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C2 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C3 = CLBLM_R_X7Y132_SLICE_X9Y132_DQ;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C4 = CLBLM_L_X12Y136_SLICE_X17Y136_BO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C5 = CLBLM_R_X11Y132_SLICE_X15Y132_DO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_C6 = CLBLL_L_X4Y134_SLICE_X4Y134_C5Q;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D1 = CLBLM_R_X11Y132_SLICE_X15Y132_AO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D2 = CLBLM_R_X11Y131_SLICE_X15Y131_AO6;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D3 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D4 = CLBLL_L_X4Y133_SLICE_X4Y133_D5Q;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D5 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_R_X11Y132_SLICE_X15Y132_D6 = CLBLM_R_X3Y137_SLICE_X3Y137_C5Q;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A1 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A2 = CLBLM_L_X8Y138_SLICE_X10Y138_A5Q;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A3 = CLBLM_R_X11Y131_SLICE_X15Y131_AO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A4 = CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A5 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_A6 = CLBLM_L_X12Y132_SLICE_X16Y132_BO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_AX = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B1 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B2 = CLBLM_R_X11Y132_SLICE_X15Y132_BO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B3 = CLBLM_L_X12Y136_SLICE_X17Y136_BO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B4 = CLBLM_R_X11Y142_SLICE_X14Y142_AQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B5 = CLBLM_R_X11Y132_SLICE_X14Y132_AO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_B6 = CLBLL_L_X4Y130_SLICE_X4Y130_B5Q;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C1 = CLBLM_R_X11Y134_SLICE_X14Y134_AO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C2 = CLBLM_L_X10Y132_SLICE_X13Y132_DO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C3 = CLBLM_R_X11Y132_SLICE_X15Y132_BO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C4 = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C5 = CLBLM_R_X11Y132_SLICE_X14Y132_DO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_C6 = CLBLM_R_X7Y133_SLICE_X9Y133_CQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B4 = CLBLM_L_X10Y140_SLICE_X13Y140_D5Q;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_T1 = 1'b1;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D1 = CLBLM_L_X12Y131_SLICE_X16Y131_AO6;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D2 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D3 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D4 = CLBLM_L_X10Y140_SLICE_X13Y140_BQ;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D5 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_R_X11Y132_SLICE_X14Y132_D6 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A1 = CLBLM_R_X5Y135_SLICE_X7Y135_CQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A3 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A4 = CLBLL_L_X4Y133_SLICE_X4Y133_BQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A5 = CLBLM_R_X5Y134_SLICE_X6Y134_C5Q;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_A6 = CLBLL_L_X4Y138_SLICE_X4Y138_AO5;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C1 = CLBLM_L_X10Y139_SLICE_X13Y139_BQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C2 = CLBLM_L_X10Y139_SLICE_X13Y139_CQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B1 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B2 = CLBLL_L_X4Y135_SLICE_X4Y135_BQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B3 = CLBLM_R_X3Y132_SLICE_X3Y132_BQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B5 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_B6 = CLBLM_R_X5Y136_SLICE_X7Y136_BQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C1 = CLBLM_R_X3Y135_SLICE_X3Y135_BQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C2 = CLBLM_R_X5Y135_SLICE_X7Y135_B5Q;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C3 = CLBLL_L_X4Y141_SLICE_X4Y141_CQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C5 = CLBLL_L_X4Y134_SLICE_X4Y134_AQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_C6 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D1 = CLBLM_R_X5Y133_SLICE_X7Y133_AQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D2 = CLBLL_L_X4Y135_SLICE_X5Y135_C5Q;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D3 = CLBLM_R_X5Y136_SLICE_X7Y136_BQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D5 = CLBLM_R_X3Y135_SLICE_X3Y135_CQ;
  assign CLBLL_L_X4Y135_SLICE_X4Y135_D6 = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_D1 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = CLBLM_L_X8Y141_SLICE_X11Y141_BQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A1 = CLBLM_L_X10Y139_SLICE_X13Y139_AQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A2 = CLBLM_L_X10Y139_SLICE_X13Y139_BQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A4 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A5 = CLBLM_L_X10Y140_SLICE_X13Y140_AQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_A6 = CLBLM_R_X11Y131_SLICE_X14Y131_BO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_D1 = CLBLM_R_X3Y141_SLICE_X2Y141_BO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_AX = CLBLM_L_X10Y139_SLICE_X12Y139_AO6;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_D1 = CLBLM_R_X3Y135_SLICE_X2Y135_AQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A1 = CLBLM_R_X5Y137_SLICE_X7Y137_B5Q;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B5 = CLBLM_R_X7Y131_SLICE_X9Y131_D5Q;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B6 = CLBLM_R_X7Y136_SLICE_X8Y136_A5Q;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A4 = CLBLL_L_X4Y135_SLICE_X5Y135_AQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A5 = CLBLL_L_X4Y134_SLICE_X5Y134_AQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_A6 = CLBLL_L_X4Y135_SLICE_X5Y135_BQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B2 = CLBLM_L_X10Y139_SLICE_X13Y139_BQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_B3 = CLBLM_R_X11Y138_SLICE_X14Y138_AQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C4 = CLBLM_L_X10Y141_SLICE_X12Y141_CQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C5 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_C6 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B2 = CLBLL_L_X4Y137_SLICE_X5Y137_D5Q;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B4 = CLBLL_L_X4Y135_SLICE_X5Y135_AQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B5 = CLBLL_L_X4Y134_SLICE_X5Y134_AQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_B6 = CLBLL_L_X4Y135_SLICE_X5Y135_BQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C2 = CLBLM_R_X5Y129_SLICE_X7Y129_B5Q;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C3 = 1'b1;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C4 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C5 = CLBLM_R_X5Y134_SLICE_X6Y134_DQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_C6 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D6 = CLBLM_R_X7Y140_SLICE_X8Y140_D5Q;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D1 = CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D2 = CLBLM_R_X11Y136_SLICE_X15Y136_AO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D3 = CLBLM_L_X10Y135_SLICE_X13Y135_CO6;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D4 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLM_L_X10Y139_SLICE_X13Y139_D5 = CLBLM_R_X11Y140_SLICE_X14Y140_BO6;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D1 = CLBLL_L_X4Y134_SLICE_X5Y134_AQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D2 = CLBLL_L_X4Y135_SLICE_X5Y135_AQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D3 = CLBLL_L_X4Y135_SLICE_X5Y135_BQ;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D5 = CLBLL_L_X4Y134_SLICE_X5Y134_D5Q;
  assign CLBLL_L_X4Y135_SLICE_X5Y135_D6 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A1 = CLBLM_R_X5Y133_SLICE_X7Y133_AQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A2 = CLBLL_L_X4Y135_SLICE_X4Y135_D5Q;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A3 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A4 = CLBLM_R_X11Y140_SLICE_X14Y140_BO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_A6 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_AX = CLBLM_L_X10Y140_SLICE_X13Y140_AQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B1 = CLBLM_L_X8Y139_SLICE_X10Y139_DO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B2 = CLBLL_L_X4Y136_SLICE_X4Y136_BQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B3 = CLBLM_L_X10Y139_SLICE_X12Y139_AQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B4 = CLBLM_R_X11Y136_SLICE_X15Y136_AO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B5 = CLBLM_L_X12Y132_SLICE_X16Y132_AO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_B6 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C1 = CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C2 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C3 = CLBLM_L_X10Y135_SLICE_X12Y135_B5Q;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C4 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C5 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_C6 = CLBLM_L_X10Y133_SLICE_X12Y133_A5Q;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D1 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D2 = CLBLM_R_X11Y136_SLICE_X14Y136_CO6;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D3 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D4 = CLBLM_R_X5Y139_SLICE_X6Y139_AQ;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D5 = 1'b1;
  assign CLBLM_L_X10Y139_SLICE_X12Y139_D6 = CLBLM_R_X7Y136_SLICE_X9Y136_BQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1 = CLBLM_R_X3Y131_SLICE_X2Y131_AO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C1 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C2 = CLBLM_R_X7Y133_SLICE_X8Y133_A5Q;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A1 = CLBLM_L_X8Y134_SLICE_X10Y134_A5Q;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A2 = CLBLM_R_X7Y137_SLICE_X8Y137_CQ;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A3 = CLBLL_L_X4Y136_SLICE_X5Y136_D5Q;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A4 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A5 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_A6 = CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B1 = CLBLM_R_X7Y134_SLICE_X9Y134_DQ;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B2 = CLBLM_R_X11Y133_SLICE_X14Y133_DO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B3 = CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B4 = CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B5 = CLBLM_L_X10Y137_SLICE_X13Y137_DO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_B6 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C1 = CLBLM_R_X3Y137_SLICE_X3Y137_C5Q;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C2 = CLBLL_L_X4Y134_SLICE_X4Y134_C5Q;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C3 = CLBLM_R_X11Y132_SLICE_X15Y132_BO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C4 = CLBLM_L_X12Y135_SLICE_X17Y135_DO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C5 = CLBLM_R_X11Y131_SLICE_X14Y131_AO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_C6 = CLBLL_L_X4Y133_SLICE_X4Y133_D5Q;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D1 = CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D2 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D3 = CLBLM_R_X11Y133_SLICE_X14Y133_DO6;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D4 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D5 = CLBLM_R_X7Y134_SLICE_X9Y134_DQ;
  assign CLBLM_R_X11Y133_SLICE_X15Y133_D6 = CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A1 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A2 = CLBLM_R_X3Y133_SLICE_X3Y133_AQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A3 = CLBLM_R_X11Y133_SLICE_X14Y133_AQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A4 = CLBLM_R_X11Y131_SLICE_X14Y131_BO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_A6 = CLBLM_L_X10Y133_SLICE_X13Y133_AQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B1 = CLBLM_R_X7Y134_SLICE_X9Y134_CQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B2 = CLBLM_R_X11Y133_SLICE_X14Y133_BQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B4 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B5 = CLBLM_L_X8Y137_SLICE_X10Y137_AQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_B6 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1 = CLBLL_L_X2Y75_SLICE_X0Y75_AO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C1 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C2 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C3 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C4 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C5 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_C6 = 1'b1;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_D = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D1 = CLBLM_L_X12Y132_SLICE_X16Y132_BO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D2 = CLBLM_R_X11Y133_SLICE_X15Y133_AO6;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D3 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D4 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D5 = CLBLM_R_X5Y133_SLICE_X7Y133_B5Q;
  assign CLBLM_R_X11Y133_SLICE_X14Y133_D6 = CLBLM_L_X10Y140_SLICE_X12Y140_D5Q;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_D = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A1 = CLBLM_L_X8Y140_SLICE_X11Y140_DO6;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A2 = CLBLM_L_X10Y137_SLICE_X13Y137_AQ;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A4 = CLBLM_R_X3Y136_SLICE_X2Y136_A5Q;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A5 = CLBLL_L_X4Y133_SLICE_X5Y133_C5Q;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_A6 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B1 = CLBLM_L_X8Y138_SLICE_X10Y138_CQ;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B2 = CLBLL_L_X4Y136_SLICE_X4Y136_BQ;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B3 = CLBLL_L_X4Y135_SLICE_X5Y135_C5Q;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B4 = CLBLL_L_X4Y136_SLICE_X4Y136_D5Q;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_B6 = CLBLM_R_X3Y136_SLICE_X3Y136_DQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_BX = CLBLL_L_X4Y138_SLICE_X4Y138_BO6;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C1 = CLBLM_R_X11Y140_SLICE_X15Y140_CO6;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C2 = CLBLL_L_X4Y136_SLICE_X4Y136_CQ;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C3 = CLBLL_L_X4Y136_SLICE_X4Y136_AQ;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C5 = CLBLM_R_X3Y136_SLICE_X3Y136_C5Q;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_C6 = CLBLL_L_X4Y136_SLICE_X4Y136_D5Q;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D1 = CLBLM_R_X5Y129_SLICE_X6Y129_AQ;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D3 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D4 = CLBLM_L_X8Y138_SLICE_X10Y138_CQ;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D5 = CLBLM_L_X8Y137_SLICE_X10Y137_DQ;
  assign CLBLL_L_X4Y136_SLICE_X4Y136_D6 = 1'b1;
  assign LIOB33_X0Y113_IOB_X0Y114_O = CLBLM_R_X3Y141_SLICE_X2Y141_BQ;
  assign LIOB33_X0Y113_IOB_X0Y113_O = CLBLL_L_X4Y130_SLICE_X4Y130_DQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A1 = CLBLM_R_X5Y133_SLICE_X7Y133_AQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A3 = CLBLM_L_X10Y140_SLICE_X13Y140_AQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A4 = CLBLL_L_X4Y135_SLICE_X4Y135_D5Q;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A5 = CLBLL_L_X4Y140_SLICE_X5Y140_C5Q;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_A6 = CLBLM_L_X8Y133_SLICE_X11Y133_B5Q;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A1 = CLBLM_R_X3Y136_SLICE_X3Y136_AQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A2 = CLBLM_L_X8Y139_SLICE_X11Y139_BQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A3 = CLBLL_L_X4Y136_SLICE_X5Y136_AQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A5 = CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_A6 = CLBLL_L_X4Y136_SLICE_X5Y136_BQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B1 = CLBLM_L_X10Y134_SLICE_X13Y134_A5Q;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B1 = CLBLL_L_X4Y137_SLICE_X5Y137_DQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B2 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B3 = CLBLL_L_X4Y130_SLICE_X5Y130_B5Q;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B4 = CLBLL_L_X4Y136_SLICE_X5Y136_CQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_B6 = CLBLM_L_X8Y137_SLICE_X10Y137_DQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A1 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A4 = CLBLM_L_X8Y131_SLICE_X11Y131_BQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A5 = CLBLM_R_X7Y134_SLICE_X8Y134_DO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A2 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A6 = CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_A3 = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B1 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C2 = CLBLL_L_X4Y136_SLICE_X5Y136_CQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C3 = CLBLM_L_X8Y137_SLICE_X10Y137_DQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C4 = CLBLL_L_X4Y136_SLICE_X5Y136_BQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C5 = CLBLL_L_X4Y137_SLICE_X5Y137_DQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_C6 = CLBLM_R_X7Y137_SLICE_X8Y137_D5Q;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B4 = CLBLM_L_X8Y131_SLICE_X10Y131_BQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B5 = CLBLM_L_X8Y130_SLICE_X11Y130_AO6;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_B6 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D1 = CLBLL_L_X4Y140_SLICE_X5Y140_DQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D3 = 1'b1;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D4 = CLBLL_L_X4Y140_SLICE_X5Y140_CQ;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D5 = CLBLL_L_X4Y131_SLICE_X5Y131_B5Q;
  assign CLBLL_L_X4Y136_SLICE_X5Y136_D6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C4 = CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C5 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_C6 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D1 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D2 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D3 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D4 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X11Y130_D5 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B1 = CLBLM_L_X8Y130_SLICE_X11Y130_BO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B2 = CLBLM_L_X10Y137_SLICE_X13Y137_A5Q;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B3 = CLBLM_R_X7Y136_SLICE_X8Y136_C5Q;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A1 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A2 = CLBLL_L_X4Y134_SLICE_X5Y134_D5Q;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A3 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A5 = CLBLM_R_X5Y133_SLICE_X6Y133_A5Q;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_A6 = CLBLM_L_X8Y130_SLICE_X10Y130_CO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C1 = CLBLM_R_X11Y139_SLICE_X14Y139_AQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C2 = CLBLM_L_X10Y140_SLICE_X12Y140_CQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C3 = CLBLM_L_X10Y134_SLICE_X12Y134_AQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B1 = CLBLM_L_X8Y131_SLICE_X11Y131_BQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B2 = CLBLM_L_X8Y138_SLICE_X11Y138_AQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B3 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B4 = CLBLM_L_X8Y131_SLICE_X10Y131_BQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B5 = CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_B6 = CLBLM_R_X7Y130_SLICE_X8Y130_DO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D1 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D2 = CLBLM_L_X10Y140_SLICE_X12Y140_AQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C1 = CLBLM_L_X8Y138_SLICE_X11Y138_AQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C2 = CLBLM_L_X8Y131_SLICE_X11Y131_BQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C3 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C4 = CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C5 = CLBLM_R_X7Y130_SLICE_X8Y130_CO6;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_C6 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D6 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D1 = CLBLM_L_X8Y138_SLICE_X11Y138_AQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D2 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D3 = CLBLM_L_X8Y131_SLICE_X11Y131_BQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D4 = CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D5 = 1'b1;
  assign CLBLM_L_X8Y130_SLICE_X10Y130_D6 = CLBLM_R_X7Y130_SLICE_X8Y130_DO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C4 = CLBLM_L_X8Y138_SLICE_X10Y138_CQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C5 = CLBLM_R_X7Y135_SLICE_X9Y135_AQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A1 = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A2 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A3 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A4 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C6 = CLBLM_R_X7Y143_SLICE_X8Y143_A5Q;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A5 = CLBLM_L_X12Y135_SLICE_X17Y135_AO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_A6 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B1 = CLBLM_R_X11Y134_SLICE_X15Y134_DO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B2 = CLBLM_L_X12Y134_SLICE_X16Y134_AO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B3 = CLBLM_R_X11Y140_SLICE_X14Y140_BO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B4 = CLBLM_R_X11Y133_SLICE_X14Y133_CO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B5 = CLBLM_R_X5Y132_SLICE_X7Y132_AQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_B6 = CLBLM_L_X10Y134_SLICE_X13Y134_AQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C1 = CLBLM_R_X5Y132_SLICE_X7Y132_AQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C2 = CLBLM_L_X10Y134_SLICE_X13Y134_AQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C3 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C4 = CLBLM_R_X11Y140_SLICE_X14Y140_BO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C5 = CLBLM_R_X11Y133_SLICE_X14Y133_CO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_C6 = CLBLM_L_X12Y134_SLICE_X16Y134_AO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D1 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D2 = CLBLM_R_X11Y136_SLICE_X14Y136_CO6;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D3 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D4 = CLBLM_R_X5Y136_SLICE_X6Y136_AQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D5 = CLBLM_L_X10Y136_SLICE_X13Y136_AQ;
  assign CLBLM_R_X11Y134_SLICE_X15Y134_D6 = 1'b1;
  assign LIOB33_SING_X0Y100_IOB_X0Y100_O = CLBLM_R_X3Y136_SLICE_X2Y136_A5Q;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A1 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A2 = CLBLM_L_X10Y140_SLICE_X13Y140_DQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A3 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A4 = CLBLM_L_X10Y134_SLICE_X13Y134_A5Q;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A5 = CLBLM_L_X12Y132_SLICE_X16Y132_BO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_A6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B1 = CLBLM_L_X8Y133_SLICE_X10Y133_C5Q;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B2 = CLBLM_R_X7Y135_SLICE_X8Y135_BO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B3 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B4 = CLBLM_L_X8Y134_SLICE_X11Y134_AQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B5 = CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_B6 = CLBLM_R_X11Y134_SLICE_X14Y134_AO5;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C1 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C2 = CLBLM_L_X10Y134_SLICE_X12Y134_CO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C3 = CLBLM_R_X11Y134_SLICE_X15Y134_BO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C4 = CLBLM_L_X10Y139_SLICE_X12Y139_BO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C5 = CLBLM_R_X11Y134_SLICE_X14Y134_DO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D5 = CLBLL_L_X4Y138_SLICE_X4Y138_BQ;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_C6 = CLBLM_R_X7Y135_SLICE_X8Y135_BO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D6 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D1 = CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D2 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D3 = CLBLM_L_X8Y133_SLICE_X10Y133_C5Q;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D4 = CLBLM_R_X11Y134_SLICE_X14Y134_AO5;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D5 = 1'b1;
  assign CLBLM_R_X11Y134_SLICE_X14Y134_D6 = CLBLM_L_X8Y134_SLICE_X11Y134_AQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A1 = CLBLL_L_X4Y131_SLICE_X4Y131_DQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A2 = CLBLL_L_X4Y139_SLICE_X4Y139_DQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A3 = CLBLL_L_X4Y137_SLICE_X4Y137_AQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A4 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_A6 = CLBLL_L_X4Y135_SLICE_X5Y135_CQ;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_D = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B1 = CLBLL_L_X4Y135_SLICE_X4Y135_DQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B2 = CLBLL_L_X4Y137_SLICE_X4Y137_BQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B3 = CLBLL_L_X4Y137_SLICE_X5Y137_C5Q;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B4 = CLBLL_L_X4Y136_SLICE_X4Y136_D5Q;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_B6 = CLBLM_L_X8Y138_SLICE_X10Y138_CQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C1 = CLBLM_R_X3Y137_SLICE_X3Y137_AQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C2 = CLBLM_R_X3Y135_SLICE_X3Y135_DQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C4 = CLBLM_R_X5Y134_SLICE_X6Y134_A5Q;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C5 = CLBLL_L_X4Y138_SLICE_X5Y138_BQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_C6 = 1'b1;
  assign LIOB33_X0Y115_IOB_X0Y116_O = CLBLM_L_X10Y131_SLICE_X12Y131_D5Q;
  assign LIOB33_X0Y115_IOB_X0Y115_O = CLBLM_R_X5Y138_SLICE_X6Y138_B5Q;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D1 = CLBLM_R_X3Y135_SLICE_X3Y135_DQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D2 = CLBLM_R_X5Y138_SLICE_X7Y138_AQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D3 = CLBLM_R_X7Y138_SLICE_X9Y138_B5Q;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D4 = CLBLM_R_X5Y138_SLICE_X7Y138_CO6;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D5 = CLBLM_R_X5Y130_SLICE_X7Y130_DQ;
  assign CLBLL_L_X4Y137_SLICE_X4Y137_D6 = CLBLM_R_X5Y137_SLICE_X7Y137_BQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A1 = CLBLM_R_X7Y133_SLICE_X8Y133_A5Q;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A2 = CLBLL_L_X4Y137_SLICE_X5Y137_BQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A3 = CLBLM_R_X3Y135_SLICE_X2Y135_BQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A4 = CLBLM_R_X5Y131_SLICE_X6Y131_BQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A5 = CLBLM_L_X10Y137_SLICE_X13Y137_AQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_A6 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A2 = CLBLM_L_X8Y141_SLICE_X11Y141_BQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A3 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B1 = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B1 = CLBLL_L_X4Y137_SLICE_X5Y137_CQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B2 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B4 = CLBLM_R_X7Y138_SLICE_X9Y138_C5Q;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B5 = CLBLL_L_X4Y133_SLICE_X5Y133_AQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_B6 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B2 = CLBLM_L_X10Y141_SLICE_X13Y141_BQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B3 = CLBLL_L_X4Y135_SLICE_X5Y135_CQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A1 = CLBLM_R_X7Y133_SLICE_X9Y133_DQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A3 = CLBLM_L_X8Y130_SLICE_X10Y130_BO6;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A4 = CLBLM_R_X5Y133_SLICE_X6Y133_A5Q;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A5 = CLBLM_L_X10Y131_SLICE_X12Y131_C5Q;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C2 = CLBLM_L_X8Y137_SLICE_X10Y137_BQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C3 = CLBLM_R_X5Y130_SLICE_X7Y130_DQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C4 = CLBLM_R_X5Y136_SLICE_X6Y136_DQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_A6 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C5 = CLBLL_L_X4Y137_SLICE_X5Y137_C5Q;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_C6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B5 = CLBLM_L_X10Y136_SLICE_X13Y136_BQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B4 = CLBLM_R_X5Y133_SLICE_X6Y133_A5Q;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B2 = CLBLM_L_X8Y131_SLICE_X11Y131_BQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B3 = CLBLM_R_X5Y133_SLICE_X7Y133_C5Q;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_B6 = CLBLM_L_X8Y130_SLICE_X11Y130_CO6;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D1 = CLBLM_R_X5Y133_SLICE_X7Y133_A5Q;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D2 = CLBLM_R_X5Y138_SLICE_X6Y138_BQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D3 = CLBLL_L_X4Y137_SLICE_X5Y137_DQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D5 = CLBLL_L_X4Y138_SLICE_X5Y138_DQ;
  assign CLBLL_L_X4Y137_SLICE_X5Y137_D6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C1 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C2 = CLBLM_L_X8Y131_SLICE_X10Y131_BQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C4 = CLBLL_L_X4Y136_SLICE_X5Y136_DQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C5 = CLBLL_L_X4Y131_SLICE_X5Y131_B5Q;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_C6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D1 = CLBLM_R_X3Y135_SLICE_X3Y135_DQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D2 = CLBLM_L_X8Y133_SLICE_X11Y133_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D3 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D5 = CLBLM_L_X8Y131_SLICE_X11Y131_AQ;
  assign CLBLM_L_X8Y131_SLICE_X11Y131_D6 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A6 = CLBLM_L_X10Y141_SLICE_X13Y141_CQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B1 = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B3 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A1 = CLBLM_R_X7Y134_SLICE_X8Y134_DO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A2 = CLBLM_L_X8Y138_SLICE_X11Y138_BQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A3 = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A4 = CLBLM_R_X5Y133_SLICE_X6Y133_A5Q;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_A6 = CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C1 = CLBLM_L_X8Y138_SLICE_X11Y138_AQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C2 = CLBLM_L_X10Y142_SLICE_X12Y142_CO6;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C3 = CLBLM_L_X10Y142_SLICE_X12Y142_BO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B2 = CLBLM_R_X5Y133_SLICE_X6Y133_A5Q;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B3 = CLBLM_L_X8Y137_SLICE_X10Y137_C5Q;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B4 = CLBLM_L_X8Y130_SLICE_X10Y130_DO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B5 = CLBLM_L_X8Y140_SLICE_X10Y140_C5Q;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_B6 = CLBLM_L_X8Y131_SLICE_X10Y131_BQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D1 = CLBLM_R_X7Y142_SLICE_X9Y142_DO5;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D2 = CLBLM_L_X10Y141_SLICE_X12Y141_AQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C1 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C2 = CLBLM_L_X8Y131_SLICE_X10Y131_CQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C4 = CLBLM_R_X7Y131_SLICE_X9Y131_BQ;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C5 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_C6 = CLBLM_L_X8Y137_SLICE_X11Y137_D5Q;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D3 = CLBLM_L_X10Y134_SLICE_X12Y134_AQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D4 = CLBLM_L_X10Y141_SLICE_X13Y141_CQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D5 = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_D6 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D1 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D2 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D3 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D4 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D5 = 1'b1;
  assign CLBLM_L_X8Y131_SLICE_X10Y131_D6 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = CLBLM_R_X3Y137_SLICE_X3Y137_D5Q;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_D1 = CLBLL_L_X4Y143_SLICE_X4Y143_AO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = CLBLM_R_X3Y139_SLICE_X2Y139_C5Q;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_T1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D1 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A1 = CLBLM_L_X10Y136_SLICE_X13Y136_AQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D2 = CLBLM_R_X5Y136_SLICE_X7Y136_CQ;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A2 = CLBLM_L_X12Y136_SLICE_X17Y136_AO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A3 = CLBLM_L_X10Y134_SLICE_X12Y134_CO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A4 = CLBLM_R_X11Y134_SLICE_X15Y134_CO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A5 = CLBLM_R_X5Y136_SLICE_X6Y136_AQ;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_A6 = CLBLM_R_X11Y136_SLICE_X15Y136_AO5;
  assign LIOB33_SING_X0Y150_IOB_X0Y150_O = CLBLM_R_X3Y134_SLICE_X2Y134_AO5;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B1 = CLBLM_R_X11Y136_SLICE_X14Y136_DO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B2 = CLBLM_R_X11Y133_SLICE_X15Y133_BO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B3 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B4 = CLBLM_L_X12Y137_SLICE_X16Y137_BO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B5 = CLBLM_L_X12Y135_SLICE_X16Y135_BO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_B6 = CLBLM_L_X10Y131_SLICE_X13Y131_DO6;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D5 = CLBLM_R_X7Y137_SLICE_X9Y137_DQ;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_T1 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D6 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C2 = CLBLM_L_X10Y135_SLICE_X13Y135_AO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C3 = CLBLM_L_X10Y134_SLICE_X13Y134_DO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C4 = CLBLM_R_X11Y133_SLICE_X15Y133_DO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C5 = CLBLM_R_X11Y135_SLICE_X15Y135_DO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_C6 = CLBLM_L_X10Y137_SLICE_X13Y137_DO6;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D1 = CLBLM_L_X12Y135_SLICE_X16Y135_AO6;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D2 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D3 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D4 = CLBLM_L_X8Y137_SLICE_X10Y137_BQ;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D5 = CLBLM_R_X3Y140_SLICE_X3Y140_C5Q;
  assign CLBLM_R_X11Y135_SLICE_X15Y135_D6 = CLBLM_L_X8Y136_SLICE_X11Y136_CO5;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A1 = CLBLM_L_X12Y137_SLICE_X17Y137_CO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A2 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A3 = CLBLM_L_X10Y135_SLICE_X13Y135_BO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A4 = CLBLM_R_X11Y135_SLICE_X14Y135_BO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A5 = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_A6 = CLBLM_L_X10Y134_SLICE_X13Y134_CO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B1 = CLBLM_R_X7Y135_SLICE_X8Y135_DO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B2 = CLBLM_L_X8Y136_SLICE_X11Y136_CO5;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B3 = CLBLM_L_X8Y137_SLICE_X11Y137_DQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B4 = CLBLM_R_X7Y133_SLICE_X8Y133_BQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B5 = CLBLM_R_X11Y133_SLICE_X14Y133_CO5;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_B6 = CLBLM_L_X8Y136_SLICE_X10Y136_CO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C1 = CLBLM_L_X10Y135_SLICE_X12Y135_CO5;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C2 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C3 = CLBLM_R_X7Y135_SLICE_X8Y135_DO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C4 = CLBLM_L_X10Y134_SLICE_X13Y134_CO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C5 = CLBLM_R_X11Y135_SLICE_X14Y135_DO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_C6 = CLBLM_L_X10Y135_SLICE_X13Y135_DO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D1 = CLBLM_L_X8Y137_SLICE_X11Y137_DQ;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D2 = CLBLM_R_X11Y133_SLICE_X14Y133_CO5;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D3 = CLBLM_L_X8Y136_SLICE_X11Y136_CO5;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D4 = CLBLM_L_X8Y136_SLICE_X10Y136_CO6;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D5 = 1'b1;
  assign CLBLM_R_X11Y135_SLICE_X14Y135_D6 = CLBLM_R_X7Y133_SLICE_X8Y133_BQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A1 = CLBLM_R_X3Y137_SLICE_X3Y137_B5Q;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A2 = CLBLL_L_X4Y135_SLICE_X4Y135_AQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A3 = CLBLM_R_X3Y136_SLICE_X2Y136_CQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A5 = CLBLL_L_X4Y138_SLICE_X5Y138_CQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_A6 = 1'b1;
  assign LIOB33_X0Y117_IOB_X0Y117_O = CLBLM_L_X10Y130_SLICE_X12Y130_B5Q;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_AX = CLBLL_L_X4Y137_SLICE_X4Y137_BQ;
  assign LIOB33_X0Y117_IOB_X0Y118_O = CLBLM_R_X5Y130_SLICE_X7Y130_CQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B1 = CLBLM_R_X11Y141_SLICE_X14Y141_AQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B2 = CLBLM_R_X7Y131_SLICE_X9Y131_D5Q;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B3 = CLBLM_R_X3Y136_SLICE_X2Y136_CQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B5 = CLBLL_L_X4Y135_SLICE_X4Y135_AQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_B6 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_BX = CLBLL_L_X4Y138_SLICE_X5Y138_CQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C1 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C2 = CLBLM_R_X3Y139_SLICE_X3Y139_AQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C3 = CLBLM_R_X5Y139_SLICE_X7Y139_A5Q;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C4 = CLBLL_L_X4Y137_SLICE_X4Y137_CQ;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C5 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_C6 = CLBLL_L_X4Y133_SLICE_X4Y133_C5Q;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D1 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D2 = CLBLM_R_X7Y138_SLICE_X9Y138_B5Q;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D3 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D4 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D5 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X4Y138_D6 = CLBLM_R_X5Y138_SLICE_X7Y138_CO6;
  assign LIOB33_SING_X0Y199_IOB_X0Y199_O = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A1 = CLBLM_R_X5Y139_SLICE_X6Y139_CQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A3 = CLBLL_L_X4Y137_SLICE_X5Y137_CQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A4 = CLBLM_R_X3Y138_SLICE_X3Y138_CO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A5 = CLBLM_L_X12Y136_SLICE_X16Y136_AQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_A6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A1 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A2 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A3 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B1 = CLBLM_R_X5Y138_SLICE_X6Y138_CQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B3 = CLBLL_L_X4Y135_SLICE_X4Y135_AQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B4 = CLBLM_L_X12Y136_SLICE_X16Y136_AQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B5 = CLBLM_R_X3Y136_SLICE_X2Y136_CQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_B6 = CLBLM_L_X8Y140_SLICE_X11Y140_AQ;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A4 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A5 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_BX = CLBLM_R_X5Y138_SLICE_X6Y138_DO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C1 = CLBLL_L_X4Y138_SLICE_X5Y138_BQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C2 = CLBLL_L_X4Y135_SLICE_X4Y135_AQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C4 = CLBLM_L_X10Y138_SLICE_X13Y138_DQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C5 = CLBLM_R_X3Y136_SLICE_X2Y136_CQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_C6 = CLBLM_L_X10Y140_SLICE_X13Y140_B5Q;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A1 = CLBLM_L_X8Y135_SLICE_X11Y135_BO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A3 = CLBLM_L_X8Y132_SLICE_X11Y132_AQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A4 = CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A5 = CLBLM_L_X10Y134_SLICE_X12Y134_AQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_A6 = 1'b1;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_CX = CLBLL_L_X4Y138_SLICE_X4Y138_AO6;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D1 = CLBLM_R_X5Y138_SLICE_X6Y138_DO5;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D3 = CLBLL_L_X4Y138_SLICE_X5Y138_DQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D4 = CLBLM_R_X5Y138_SLICE_X7Y138_AQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D5 = CLBLM_R_X5Y130_SLICE_X7Y130_DQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_D6 = CLBLL_L_X4Y140_SLICE_X4Y140_AQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B2 = CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  assign CLBLL_L_X4Y138_SLICE_X5Y138_DX = CLBLL_L_X4Y140_SLICE_X4Y140_DO5;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B3 = CLBLM_L_X10Y132_SLICE_X12Y132_AQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B4 = CLBLM_L_X8Y135_SLICE_X10Y135_C5Q;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B5 = CLBLM_L_X8Y132_SLICE_X11Y132_BQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_B6 = CLBLM_L_X8Y132_SLICE_X11Y132_AO5;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C1 = CLBLM_L_X8Y132_SLICE_X11Y132_BQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C2 = CLBLM_L_X10Y132_SLICE_X12Y132_AQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C3 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C4 = CLBLM_L_X8Y135_SLICE_X11Y135_BO6;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C5 = CLBLM_L_X8Y132_SLICE_X11Y132_AQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_C6 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A1 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A2 = CLBLM_L_X10Y133_SLICE_X12Y133_A5Q;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D1 = CLBLM_L_X10Y133_SLICE_X12Y133_AQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D2 = CLBLL_L_X4Y132_SLICE_X4Y132_DQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D3 = CLBLM_R_X3Y132_SLICE_X3Y132_CQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D4 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D5 = CLBLL_L_X4Y132_SLICE_X5Y132_DQ;
  assign CLBLM_L_X8Y132_SLICE_X11Y132_D6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A5 = CLBLM_L_X8Y142_SLICE_X11Y142_CO5;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A6 = CLBLM_L_X8Y141_SLICE_X10Y141_CO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B1 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B2 = CLBLM_L_X8Y141_SLICE_X11Y141_BQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B3 = CLBLM_L_X10Y141_SLICE_X12Y141_C5Q;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A2 = CLBLM_R_X7Y132_SLICE_X9Y132_CQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A3 = CLBLL_L_X4Y136_SLICE_X4Y136_B5Q;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A4 = CLBLM_R_X11Y142_SLICE_X14Y142_AQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A5 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_A6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C1 = CLBLM_L_X8Y141_SLICE_X11Y141_BQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C2 = CLBLM_L_X10Y141_SLICE_X12Y141_CQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C3 = CLBLM_L_X8Y142_SLICE_X11Y142_DO6;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B1 = CLBLM_L_X10Y140_SLICE_X13Y140_B5Q;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B2 = CLBLL_L_X4Y131_SLICE_X4Y131_CQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B3 = CLBLM_L_X10Y134_SLICE_X12Y134_B5Q;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B5 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_B6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D1 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D2 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C1 = CLBLM_R_X7Y131_SLICE_X9Y131_D5Q;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C2 = CLBLM_L_X8Y132_SLICE_X10Y132_CQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C3 = CLBLM_L_X10Y130_SLICE_X12Y130_AQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C4 = CLBLM_L_X10Y140_SLICE_X13Y140_D5Q;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_C6 = CLBLM_R_X7Y135_SLICE_X9Y135_D5Q;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D3 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D4 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D5 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_D6 = 1'b1;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D1 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D2 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D3 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D4 = CLBLM_L_X8Y131_SLICE_X10Y131_CQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D5 = CLBLM_R_X7Y132_SLICE_X9Y132_AQ;
  assign CLBLM_L_X8Y132_SLICE_X10Y132_D6 = CLBLM_R_X11Y132_SLICE_X15Y132_AO5;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A1 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A2 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A3 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A4 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A5 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_A6 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_AX = CLBLM_R_X11Y136_SLICE_X14Y136_AQ;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B1 = CLBLM_L_X10Y136_SLICE_X13Y136_DO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B2 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B3 = CLBLM_R_X11Y135_SLICE_X15Y135_AO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B4 = CLBLM_R_X11Y134_SLICE_X14Y134_BO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B5 = CLBLM_R_X11Y138_SLICE_X15Y138_AO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_B6 = CLBLM_L_X10Y139_SLICE_X12Y139_BO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C1 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C2 = CLBLM_R_X11Y140_SLICE_X14Y140_BO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C3 = CLBLL_L_X4Y137_SLICE_X4Y137_AQ;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C4 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C5 = CLBLM_R_X11Y132_SLICE_X15Y132_AO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_C6 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D1 = CLBLM_R_X11Y138_SLICE_X15Y138_AO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D2 = CLBLM_R_X11Y134_SLICE_X14Y134_CO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D3 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D4 = CLBLM_L_X10Y136_SLICE_X13Y136_DO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D5 = CLBLM_L_X12Y137_SLICE_X16Y137_DO6;
  assign CLBLM_R_X11Y136_SLICE_X15Y136_D6 = CLBLM_R_X11Y135_SLICE_X15Y135_CO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A1 = CLBLM_R_X7Y138_SLICE_X8Y138_CQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A2 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A3 = CLBLM_R_X11Y136_SLICE_X14Y136_AQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A4 = CLBLM_L_X10Y136_SLICE_X12Y136_AQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A5 = CLBLM_R_X13Y134_SLICE_X18Y134_AO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B1 = CLBLM_R_X11Y140_SLICE_X15Y140_BQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B2 = CLBLM_L_X12Y131_SLICE_X16Y131_AO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B3 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B4 = CLBLL_L_X4Y140_SLICE_X4Y140_AQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B5 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_B6 = CLBLM_L_X12Y140_SLICE_X16Y140_AO5;
  assign LIOB33_X0Y119_IOB_X0Y119_O = CLBLM_R_X3Y132_SLICE_X3Y132_BQ;
  assign LIOB33_X0Y119_IOB_X0Y120_O = CLBLM_R_X5Y138_SLICE_X7Y138_AQ;
  assign RIOB33_X105Y197_IOB_X1Y198_O = CLBLM_L_X12Y143_SLICE_X16Y143_AO5;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C1 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C2 = CLBLM_R_X7Y137_SLICE_X8Y137_CQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C3 = CLBLL_L_X4Y136_SLICE_X5Y136_D5Q;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C4 = CLBLM_L_X8Y134_SLICE_X10Y134_A5Q;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C5 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_C6 = CLBLM_L_X10Y135_SLICE_X12Y135_AQ;
  assign RIOB33_X105Y197_IOB_X1Y197_O = CLBLM_R_X11Y140_SLICE_X14Y140_AO5;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D1 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D2 = CLBLM_R_X11Y134_SLICE_X14Y134_AO6;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D3 = CLBLM_R_X7Y133_SLICE_X9Y133_CQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D4 = CLBLM_L_X12Y136_SLICE_X17Y136_BO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A1 = CLBLM_R_X5Y137_SLICE_X7Y137_BQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A3 = CLBLM_R_X3Y139_SLICE_X3Y139_BO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A4 = CLBLM_R_X7Y137_SLICE_X8Y137_BQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A5 = CLBLM_R_X3Y136_SLICE_X3Y136_C5Q;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_A6 = 1'b1;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D5 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_R_X11Y136_SLICE_X14Y136_D6 = CLBLM_L_X10Y140_SLICE_X13Y140_BQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B1 = CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B2 = CLBLL_L_X4Y139_SLICE_X5Y139_DO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B3 = CLBLL_L_X4Y138_SLICE_X5Y138_AQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B5 = CLBLL_L_X4Y139_SLICE_X4Y139_BQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_B6 = CLBLL_L_X4Y141_SLICE_X5Y141_BO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C1 = CLBLL_L_X4Y137_SLICE_X4Y137_BQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C2 = CLBLL_L_X4Y139_SLICE_X4Y139_CQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C3 = CLBLM_L_X12Y132_SLICE_X16Y132_AO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C4 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C5 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D1 = CLBLM_R_X5Y141_SLICE_X7Y141_AO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D2 = CLBLM_R_X7Y136_SLICE_X8Y136_B5Q;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D3 = CLBLL_L_X4Y139_SLICE_X4Y139_DQ;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D4 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D5 = CLBLL_L_X4Y140_SLICE_X4Y140_CO6;
  assign CLBLL_L_X4Y139_SLICE_X4Y139_D6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_D = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A1 = CLBLM_R_X5Y130_SLICE_X6Y130_B5Q;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A2 = CLBLM_R_X7Y138_SLICE_X9Y138_C5Q;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A3 = CLBLL_L_X4Y139_SLICE_X5Y139_AQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A5 = CLBLL_L_X4Y136_SLICE_X4Y136_D5Q;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_A6 = CLBLM_L_X8Y138_SLICE_X10Y138_CQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B2 = CLBLL_L_X4Y139_SLICE_X5Y139_BQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B3 = CLBLL_L_X4Y140_SLICE_X5Y140_AQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B4 = CLBLM_R_X3Y139_SLICE_X2Y139_AQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B5 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_B6 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_D = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C1 = CLBLM_R_X5Y139_SLICE_X7Y139_BQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C2 = CLBLM_L_X8Y135_SLICE_X11Y135_AQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C3 = CLBLM_R_X5Y140_SLICE_X7Y140_B5Q;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C4 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_C6 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A1 = CLBLM_L_X8Y137_SLICE_X11Y137_CQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A2 = CLBLM_L_X10Y134_SLICE_X13Y134_AQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A3 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A5 = CLBLL_L_X4Y137_SLICE_X4Y137_C5Q;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D1 = CLBLM_R_X7Y140_SLICE_X8Y140_C5Q;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D2 = CLBLM_R_X3Y139_SLICE_X2Y139_AQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D3 = CLBLM_R_X5Y129_SLICE_X7Y129_B5Q;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D4 = CLBLM_R_X3Y139_SLICE_X2Y139_BQ;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D5 = 1'b1;
  assign CLBLL_L_X4Y139_SLICE_X5Y139_D6 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B1 = CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_A6 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B2 = CLBLM_R_X5Y137_SLICE_X7Y137_AQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B3 = CLBLM_R_X5Y130_SLICE_X7Y130_AQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C1 = CLBLM_R_X7Y133_SLICE_X9Y133_C5Q;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C2 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C3 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C4 = CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C5 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_C6 = CLBLM_L_X8Y137_SLICE_X11Y137_D5Q;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D1 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D2 = CLBLL_L_X4Y132_SLICE_X4Y132_DQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D3 = CLBLM_R_X3Y132_SLICE_X3Y132_CQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D4 = CLBLM_R_X5Y133_SLICE_X7Y133_B5Q;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D5 = CLBLM_R_X7Y134_SLICE_X8Y134_A5Q;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_D6 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A1 = CLBLM_L_X8Y131_SLICE_X11Y131_DQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A2 = CLBLL_L_X4Y136_SLICE_X4Y136_D5Q;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A3 = CLBLM_L_X8Y133_SLICE_X10Y133_AQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A4 = CLBLM_L_X10Y134_SLICE_X13Y134_AQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A5 = CLBLM_L_X8Y138_SLICE_X10Y138_CQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B1 = CLBLM_L_X8Y138_SLICE_X10Y138_CQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B2 = CLBLM_L_X8Y133_SLICE_X10Y133_BQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B3 = CLBLM_L_X10Y132_SLICE_X12Y132_BQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B4 = CLBLL_L_X4Y136_SLICE_X4Y136_D5Q;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B5 = CLBLM_R_X5Y131_SLICE_X7Y131_D5Q;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C1 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C2 = CLBLM_L_X8Y132_SLICE_X10Y132_CQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C3 = CLBLM_L_X8Y133_SLICE_X10Y133_C5Q;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C4 = CLBLM_R_X5Y134_SLICE_X6Y134_CQ;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D1 = CLBLM_L_X8Y136_SLICE_X11Y136_CO5;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D2 = CLBLM_L_X8Y134_SLICE_X10Y134_CO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D3 = CLBLM_L_X8Y132_SLICE_X10Y132_A5Q;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D4 = CLBLM_L_X8Y132_SLICE_X10Y132_DO6;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D5 = CLBLM_R_X11Y133_SLICE_X14Y133_CO5;
  assign CLBLM_L_X8Y133_SLICE_X10Y133_D6 = CLBLM_R_X5Y132_SLICE_X7Y132_BQ;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A1 = CLBLM_L_X12Y137_SLICE_X17Y137_AO5;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A2 = CLBLM_R_X7Y135_SLICE_X8Y135_BQ;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A3 = CLBLM_R_X11Y134_SLICE_X15Y134_AO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A4 = CLBLM_R_X13Y134_SLICE_X18Y134_AO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A5 = CLBLM_R_X13Y137_SLICE_X18Y137_AO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_A6 = CLBLL_L_X4Y131_SLICE_X4Y131_CQ;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B1 = CLBLM_L_X10Y131_SLICE_X12Y131_AQ;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B2 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B3 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B4 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B5 = CLBLM_L_X12Y138_SLICE_X16Y138_AO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_B6 = CLBLM_R_X11Y140_SLICE_X14Y140_BO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_C5 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C1 = CLBLM_L_X12Y139_SLICE_X16Y139_AO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C2 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C3 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C4 = CLBLM_R_X11Y140_SLICE_X14Y140_BO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C5 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_C6 = CLBLL_L_X4Y139_SLICE_X4Y139_CQ;
  assign LIOB33_X0Y121_IOB_X0Y121_O = CLBLM_R_X7Y135_SLICE_X9Y135_C5Q;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D1 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D2 = CLBLM_R_X11Y140_SLICE_X14Y140_BO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D3 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D4 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D5 = CLBLM_L_X10Y131_SLICE_X13Y131_AQ;
  assign CLBLM_R_X11Y137_SLICE_X15Y137_D6 = CLBLM_L_X10Y137_SLICE_X12Y137_AO6;
  assign CLBLM_R_X5Y129_SLICE_X6Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOB33_X0Y121_IOB_X0Y122_O = CLBLL_L_X4Y136_SLICE_X4Y136_CQ;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A1 = CLBLM_R_X11Y138_SLICE_X15Y138_CO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A2 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A3 = CLBLM_L_X8Y133_SLICE_X10Y133_DO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A4 = CLBLM_R_X11Y132_SLICE_X14Y132_BO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A5 = CLBLM_L_X12Y133_SLICE_X17Y133_AO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_A6 = CLBLM_R_X11Y137_SLICE_X14Y137_CO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B1 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B2 = CLBLM_R_X7Y136_SLICE_X8Y136_AQ;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B3 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B4 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B5 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_B6 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C1 = CLBLM_L_X10Y134_SLICE_X13Y134_BO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C2 = CLBLM_R_X11Y137_SLICE_X15Y137_CO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C3 = CLBLM_R_X11Y137_SLICE_X15Y137_DO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C4 = CLBLM_R_X11Y137_SLICE_X15Y137_BO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C5 = CLBLM_L_X8Y138_SLICE_X11Y138_DO6;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_C6 = CLBLM_R_X11Y137_SLICE_X14Y137_BO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_D1 = CLBLM_R_X3Y132_SLICE_X3Y132_BQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B3 = CLBLM_R_X11Y136_SLICE_X15Y136_BO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A1 = CLBLL_L_X4Y131_SLICE_X5Y131_B5Q;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A3 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A4 = CLBLL_L_X4Y141_SLICE_X4Y141_BQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A5 = CLBLL_L_X4Y141_SLICE_X4Y141_AQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_A6 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B4 = CLBLM_L_X10Y137_SLICE_X13Y137_A5Q;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_AX = CLBLM_R_X5Y133_SLICE_X7Y133_AQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B5 = CLBLM_R_X11Y135_SLICE_X15Y135_BO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B1 = CLBLL_L_X4Y141_SLICE_X4Y141_DQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B2 = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B3 = CLBLL_L_X4Y140_SLICE_X5Y140_DQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B4 = CLBLM_R_X3Y140_SLICE_X3Y140_DQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B5 = CLBLL_L_X4Y139_SLICE_X4Y139_DQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_B6 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_B6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_D1 = CLBLL_L_X4Y134_SLICE_X5Y134_DQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C1 = CLBLL_L_X4Y139_SLICE_X4Y139_DQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C2 = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C3 = CLBLL_L_X4Y141_SLICE_X4Y141_DQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C4 = CLBLM_R_X3Y140_SLICE_X3Y140_DQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C5 = CLBLL_L_X4Y140_SLICE_X5Y140_DQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_C6 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_T1 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_D1 = CLBLM_R_X7Y141_SLICE_X8Y141_CO6;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D1 = CLBLL_L_X4Y138_SLICE_X5Y138_C5Q;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D2 = CLBLL_L_X4Y139_SLICE_X4Y139_A5Q;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D3 = CLBLL_L_X4Y140_SLICE_X4Y140_AQ;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D4 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y140_SLICE_X4Y140_D6 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C1 = CLBLL_L_X4Y140_SLICE_X5Y140_C5Q;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_T1 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C3 = CLBLM_R_X5Y140_SLICE_X6Y140_CQ;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C4 = CLBLM_L_X12Y140_SLICE_X16Y140_AQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C5 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1 = CLBLL_L_X4Y142_SLICE_X4Y142_BO6;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_C6 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A1 = CLBLL_L_X4Y136_SLICE_X4Y136_DQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A2 = CLBLL_L_X4Y138_SLICE_X5Y138_B5Q;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A3 = CLBLL_L_X4Y140_SLICE_X5Y140_AQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A5 = CLBLM_R_X7Y135_SLICE_X9Y135_C5Q;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_A6 = CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B1 = CLBLL_L_X4Y136_SLICE_X4Y136_DQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B3 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B4 = CLBLM_R_X11Y132_SLICE_X14Y132_AQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B5 = CLBLM_R_X3Y135_SLICE_X2Y135_AQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_B6 = CLBLL_L_X4Y141_SLICE_X5Y141_CO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C1 = CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C2 = CLBLL_L_X4Y138_SLICE_X5Y138_DQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C3 = CLBLL_L_X4Y134_SLICE_X5Y134_BQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C5 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_C6 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_X105Y177_IOB_X1Y178_O = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A1 = CLBLM_R_X3Y134_SLICE_X3Y134_BQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D1 = CLBLL_L_X4Y139_SLICE_X5Y139_AQ;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D2 = 1'b1;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D4 = CLBLL_L_X4Y140_SLICE_X4Y140_BO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D5 = CLBLM_R_X5Y141_SLICE_X7Y141_AO6;
  assign CLBLL_L_X4Y140_SLICE_X5Y140_D6 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A2 = CLBLM_L_X10Y140_SLICE_X13Y140_D5Q;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A3 = CLBLM_L_X8Y134_SLICE_X11Y134_AQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A4 = CLBLM_R_X7Y136_SLICE_X9Y136_D5Q;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A5 = CLBLM_R_X7Y131_SLICE_X9Y131_D5Q;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B1 = CLBLM_R_X7Y140_SLICE_X9Y140_D5Q;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B2 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B3 = CLBLM_R_X7Y133_SLICE_X9Y133_C5Q;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B5 = CLBLM_R_X5Y133_SLICE_X7Y133_C5Q;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_B6 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C1 = CLBLM_R_X3Y133_SLICE_X3Y133_BQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C2 = CLBLM_L_X8Y135_SLICE_X11Y135_CO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C3 = CLBLM_L_X10Y134_SLICE_X12Y134_DO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C4 = CLBLM_L_X8Y135_SLICE_X11Y135_DO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C5 = CLBLM_L_X8Y133_SLICE_X11Y133_DO6;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_C6 = CLBLM_L_X8Y132_SLICE_X11Y132_AQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D3 = CLBLM_R_X3Y140_SLICE_X3Y140_AQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D4 = CLBLM_L_X8Y140_SLICE_X10Y140_AQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D5 = CLBLM_L_X10Y140_SLICE_X13Y140_B5Q;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D1 = CLBLL_L_X4Y136_SLICE_X5Y136_AQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D2 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D3 = CLBLM_R_X7Y137_SLICE_X8Y137_B5Q;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D4 = CLBLM_L_X8Y132_SLICE_X11Y132_AQ;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D5 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X11Y134_D6 = CLBLM_R_X5Y136_SLICE_X6Y136_BQ;
  assign CLBLM_L_X10Y140_SLICE_X13Y140_D6 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A1 = CLBLL_L_X4Y139_SLICE_X5Y139_CQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A2 = CLBLM_R_X11Y141_SLICE_X14Y141_AQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A3 = CLBLM_L_X8Y136_SLICE_X11Y136_B5Q;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A5 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_A6 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B1 = CLBLM_L_X8Y136_SLICE_X10Y136_DO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B2 = CLBLM_L_X8Y132_SLICE_X11Y132_BQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B3 = CLBLM_L_X8Y132_SLICE_X11Y132_DO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B4 = CLBLM_L_X8Y134_SLICE_X10Y134_DO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B5 = CLBLM_R_X7Y132_SLICE_X9Y132_DQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_B6 = CLBLM_L_X8Y134_SLICE_X11Y134_DO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C1 = CLBLM_R_X11Y133_SLICE_X15Y133_AO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C2 = CLBLM_R_X7Y132_SLICE_X9Y132_A5Q;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C3 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C4 = CLBLM_R_X7Y136_SLICE_X9Y136_A5Q;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C5 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_C6 = CLBLM_R_X5Y134_SLICE_X6Y134_A5Q;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A1 = CLBLM_L_X8Y130_SLICE_X11Y130_BO6;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A2 = CLBLM_L_X10Y140_SLICE_X12Y140_BQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D1 = CLBLM_L_X10Y132_SLICE_X12Y132_AQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D2 = CLBLM_R_X7Y136_SLICE_X8Y136_BQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D3 = CLBLM_R_X7Y136_SLICE_X9Y136_CQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D4 = 1'b1;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D5 = CLBLM_R_X3Y136_SLICE_X3Y136_AQ;
  assign CLBLM_L_X8Y134_SLICE_X10Y134_D6 = CLBLM_L_X8Y138_SLICE_X10Y138_A5Q;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A4 = CLBLM_R_X11Y140_SLICE_X15Y140_AQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A5 = CLBLM_L_X10Y140_SLICE_X12Y140_AQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_A6 = CLBLM_R_X5Y133_SLICE_X6Y133_A5Q;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_D = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_D = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A1 = CLBLM_R_X11Y140_SLICE_X15Y140_DO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A2 = CLBLM_L_X12Y139_SLICE_X16Y139_BO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A3 = CLBLM_L_X10Y136_SLICE_X12Y136_BQ;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A4 = CLBLM_L_X12Y133_SLICE_X17Y133_AO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A5 = CLBLM_L_X12Y135_SLICE_X17Y135_BO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_A6 = CLBLM_L_X12Y137_SLICE_X17Y137_BO6;
  assign LIOB33_X0Y123_IOB_X0Y123_O = CLBLM_R_X3Y132_SLICE_X3Y132_BQ;
  assign LIOB33_X0Y123_IOB_X0Y124_O = CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B1 = CLBLM_L_X12Y136_SLICE_X17Y136_AO5;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B2 = CLBLM_L_X12Y135_SLICE_X17Y135_CO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B3 = CLBLM_L_X12Y138_SLICE_X16Y138_AO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B4 = RIOB33_X105Y145_IOB_X1Y145_I;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B5 = CLBLM_L_X12Y131_SLICE_X16Y131_AO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_B6 = CLBLM_L_X10Y138_SLICE_X12Y138_BQ;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C1 = CLBLM_L_X12Y138_SLICE_X17Y138_AO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C2 = CLBLM_L_X12Y138_SLICE_X16Y138_AO5;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C3 = CLBLM_R_X11Y139_SLICE_X15Y139_AO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C4 = CLBLM_R_X11Y136_SLICE_X15Y136_CO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C5 = CLBLM_R_X13Y134_SLICE_X18Y134_AO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B5 = CLBLM_L_X10Y140_SLICE_X12Y140_BQ;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_C6 = CLBLM_R_X11Y138_SLICE_X15Y138_BO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_B6 = CLBLM_R_X5Y133_SLICE_X6Y133_A5Q;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D1 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D2 = CLBLM_L_X12Y137_SLICE_X17Y137_CO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D3 = CLBLM_R_X11Y138_SLICE_X14Y138_DO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D4 = CLBLM_L_X12Y138_SLICE_X17Y138_BO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D5 = CLBLM_L_X10Y133_SLICE_X13Y133_DO6;
  assign CLBLM_R_X11Y138_SLICE_X15Y138_D6 = CLBLM_R_X11Y135_SLICE_X14Y135_CO6;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y120_D = RIOB33_X105Y119_IOB_X1Y120_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A1 = CLBLM_L_X10Y139_SLICE_X13Y139_CQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A2 = CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A3 = CLBLM_L_X8Y138_SLICE_X10Y138_BQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A4 = CLBLM_L_X10Y137_SLICE_X13Y137_CO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A5 = CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_A6 = CLBLM_L_X10Y138_SLICE_X12Y138_DO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_AX = CLBLM_L_X10Y138_SLICE_X13Y138_AQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B1 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B2 = CLBLM_L_X12Y139_SLICE_X16Y139_AO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B3 = CLBLM_L_X8Y138_SLICE_X10Y138_BQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B4 = CLBLM_L_X12Y131_SLICE_X16Y131_BO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B5 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_B6 = CLBLM_L_X10Y139_SLICE_X13Y139_CQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C1 = CLBLM_L_X10Y134_SLICE_X12Y134_BQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C2 = CLBLM_R_X11Y139_SLICE_X14Y139_BO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C3 = 1'b1;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C4 = CLBLM_L_X8Y136_SLICE_X11Y136_CO5;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C5 = CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_C6 = CLBLM_L_X10Y138_SLICE_X13Y138_AQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A1 = CLBLM_R_X5Y142_SLICE_X6Y142_B5Q;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A2 = CLBLL_L_X4Y141_SLICE_X4Y141_BQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A3 = CLBLM_R_X3Y139_SLICE_X3Y139_AQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A4 = CLBLL_L_X4Y141_SLICE_X4Y141_CQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_A6 = CLBLL_L_X4Y141_SLICE_X4Y141_AQ;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C5 = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_C6 = CLBLM_R_X5Y140_SLICE_X7Y140_A5Q;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B1 = CLBLM_R_X5Y142_SLICE_X6Y142_B5Q;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B2 = CLBLL_L_X4Y141_SLICE_X4Y141_BQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B3 = CLBLL_L_X4Y141_SLICE_X4Y141_CQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B4 = CLBLL_L_X4Y141_SLICE_X4Y141_AQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_B6 = CLBLL_L_X4Y136_SLICE_X4Y136_CQ;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D2 = CLBLM_R_X7Y135_SLICE_X8Y135_CO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D3 = CLBLM_L_X10Y137_SLICE_X13Y137_CO6;
  assign CLBLM_R_X11Y138_SLICE_X14Y138_D5 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C1 = CLBLL_L_X4Y141_SLICE_X4Y141_BQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C2 = CLBLL_L_X4Y141_SLICE_X4Y141_CQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C4 = CLBLL_L_X4Y138_SLICE_X5Y138_A5Q;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C5 = CLBLM_R_X5Y142_SLICE_X6Y142_B5Q;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_C6 = CLBLL_L_X4Y141_SLICE_X4Y141_AQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D1 = CLBLM_R_X5Y141_SLICE_X7Y141_AO6;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D2 = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D3 = CLBLL_L_X4Y141_SLICE_X4Y141_DQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D4 = CLBLM_R_X3Y140_SLICE_X3Y140_DQ;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y141_SLICE_X4Y141_D6 = CLBLL_L_X4Y130_SLICE_X4Y130_D5Q;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A2 = CLBLM_R_X5Y141_SLICE_X7Y141_AO5;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A3 = CLBLL_L_X4Y141_SLICE_X5Y141_AQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A4 = CLBLM_R_X5Y141_SLICE_X7Y141_BO6;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A5 = CLBLM_R_X5Y136_SLICE_X6Y136_AQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_A6 = CLBLM_L_X10Y130_SLICE_X12Y130_B5Q;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D3 = CLBLM_L_X8Y138_SLICE_X10Y138_DQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B2 = CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B3 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B4 = CLBLM_R_X3Y135_SLICE_X2Y135_AQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B5 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_B6 = 1'b1;
  assign CLBLM_L_X10Y140_SLICE_X12Y140_D5 = CLBLM_L_X10Y140_SLICE_X13Y140_BQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C1 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C2 = CLBLL_L_X4Y139_SLICE_X4Y139_AQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C3 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C5 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_C6 = CLBLM_L_X8Y140_SLICE_X10Y140_DQ;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D1 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D2 = CLBLM_L_X8Y140_SLICE_X10Y140_C5Q;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D3 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D4 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D5 = 1'b1;
  assign CLBLL_L_X4Y141_SLICE_X5Y141_D6 = CLBLM_R_X7Y137_SLICE_X8Y137_C5Q;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A1 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A2 = CLBLM_L_X8Y137_SLICE_X11Y137_BQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A4 = CLBLM_R_X3Y135_SLICE_X3Y135_A5Q;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A5 = CLBLM_R_X3Y136_SLICE_X3Y136_AQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_A6 = CLBLM_L_X8Y134_SLICE_X11Y134_CO6;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B1 = CLBLM_R_X7Y136_SLICE_X9Y136_CQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B2 = CLBLM_L_X8Y136_SLICE_X11Y136_AQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B3 = CLBLL_L_X4Y136_SLICE_X5Y136_AQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B4 = CLBLM_L_X8Y139_SLICE_X11Y139_BQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B5 = CLBLM_R_X3Y136_SLICE_X3Y136_AQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_B6 = CLBLM_L_X8Y137_SLICE_X11Y137_BQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C1 = CLBLM_L_X8Y132_SLICE_X10Y132_A5Q;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C2 = CLBLM_L_X8Y136_SLICE_X11Y136_AQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C3 = CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C4 = CLBLM_L_X8Y137_SLICE_X11Y137_BQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C5 = CLBLM_R_X7Y136_SLICE_X9Y136_CQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_C6 = CLBLM_L_X8Y137_SLICE_X11Y137_DQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D1 = CLBLL_L_X4Y136_SLICE_X5Y136_AQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D2 = CLBLM_L_X8Y137_SLICE_X10Y137_BQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D3 = CLBLM_L_X10Y140_SLICE_X13Y140_DQ;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D4 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D5 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X11Y135_D6 = CLBLM_L_X8Y139_SLICE_X11Y139_BQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A1 = CLBLM_R_X7Y135_SLICE_X9Y135_CQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A2 = CLBLM_L_X8Y132_SLICE_X10Y132_A5Q;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A3 = CLBLM_L_X8Y135_SLICE_X10Y135_AQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_A6 = CLBLM_R_X7Y135_SLICE_X9Y135_B5Q;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B1 = CLBLM_L_X12Y136_SLICE_X16Y136_A5Q;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B2 = CLBLM_R_X7Y133_SLICE_X8Y133_BQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B3 = CLBLM_L_X8Y135_SLICE_X10Y135_AQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B4 = CLBLM_R_X7Y132_SLICE_X9Y132_A5Q;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_B6 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C2 = CLBLM_R_X7Y136_SLICE_X8Y136_CQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C3 = CLBLM_R_X5Y135_SLICE_X7Y135_CQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C4 = CLBLM_L_X12Y136_SLICE_X16Y136_A5Q;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C5 = CLBLM_L_X8Y136_SLICE_X11Y136_AQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_C6 = 1'b1;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D2 = CLBLM_L_X8Y131_SLICE_X11Y131_DQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D3 = CLBLM_R_X7Y135_SLICE_X9Y135_CQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D4 = CLBLM_R_X3Y133_SLICE_X3Y133_B5Q;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D5 = CLBLM_R_X5Y132_SLICE_X6Y132_BQ;
  assign CLBLM_L_X8Y135_SLICE_X10Y135_D6 = 1'b1;
  assign LIOB33_X0Y125_IOB_X0Y126_O = CLBLM_R_X5Y133_SLICE_X7Y133_AQ;
  assign LIOB33_X0Y125_IOB_X0Y125_O = CLBLM_L_X8Y138_SLICE_X10Y138_CQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C2 = CLBLM_R_X3Y138_SLICE_X2Y138_CQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C3 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A1 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A2 = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A3 = CLBLM_L_X12Y135_SLICE_X17Y135_AO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A4 = CLBLM_L_X10Y137_SLICE_X12Y137_AO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C4 = CLBLM_R_X7Y138_SLICE_X9Y138_A5Q;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A5 = CLBLM_R_X11Y139_SLICE_X14Y139_AQ;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_A6 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B1 = CLBLM_R_X7Y139_SLICE_X9Y139_DO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B2 = CLBLM_R_X11Y138_SLICE_X15Y138_DO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B3 = CLBLM_R_X11Y139_SLICE_X14Y139_AO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B4 = CLBLM_R_X11Y136_SLICE_X15Y136_DO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C6 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_B6 = CLBLM_R_X11Y139_SLICE_X15Y139_CO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A2 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A3 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A4 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A5 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_A6 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C1 = CLBLM_R_X11Y138_SLICE_X14Y138_CO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C2 = CLBLM_L_X10Y139_SLICE_X13Y139_DO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_C3 = CLBLM_L_X12Y136_SLICE_X17Y136_CO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B2 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B3 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B4 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B5 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_B6 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D1 = CLBLM_L_X12Y133_SLICE_X17Y133_AO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D2 = CLBLM_L_X10Y133_SLICE_X13Y133_BO6;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C2 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C3 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C4 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C5 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_C6 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D3 = CLBLM_R_X3Y139_SLICE_X3Y139_BO6;
  assign CLBLM_R_X11Y139_SLICE_X15Y139_D4 = CLBLM_L_X12Y139_SLICE_X16Y139_CO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A1 = CLBLM_R_X11Y137_SLICE_X14Y137_DO6;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A3 = CLBLM_R_X11Y140_SLICE_X15Y140_B5Q;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A4 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_A6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D2 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D3 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D4 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D5 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X9Y129_D6 = 1'b1;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_AX = CLBLM_R_X11Y140_SLICE_X14Y140_CQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B1 = CLBLM_L_X12Y140_SLICE_X16Y140_AO5;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D1 = CLBLM_R_X5Y135_SLICE_X6Y135_CO5;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B2 = CLBLM_L_X10Y131_SLICE_X12Y131_BQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B3 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_R_X11Y139_SLICE_X14Y139_B4 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A2 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A3 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A4 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A5 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_A6 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D2 = CLBLM_R_X11Y138_SLICE_X15Y138_CO6;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A2 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A3 = CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A4 = CLBLL_L_X4Y143_SLICE_X5Y143_BO5;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A5 = CLBLL_L_X4Y139_SLICE_X5Y139_BQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_A6 = CLBLM_R_X5Y141_SLICE_X7Y141_AO6;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_AX = CLBLM_R_X7Y134_SLICE_X8Y134_AQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B1 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_AX = CLBLL_L_X4Y142_SLICE_X4Y142_BO5;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B2 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B2 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B4 = CLBLM_L_X12Y141_SLICE_X16Y141_AQ;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B5 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_B6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B4 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B5 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C1 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C2 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C3 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C4 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C5 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_C6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C3 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C4 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A3 = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D3 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D4 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D5 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D6 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_A6 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D1 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X4Y142_D2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B3 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_B6 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C3 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_C6 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_D1 = CLBLM_L_X12Y142_SLICE_X16Y142_BO5;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D3 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X0Y75_D6 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A1 = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A3 = CLBLL_L_X4Y141_SLICE_X4Y141_AQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A4 = CLBLL_L_X4Y141_SLICE_X4Y141_BQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A5 = CLBLM_R_X5Y135_SLICE_X6Y135_B5Q;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_A6 = CLBLM_R_X5Y142_SLICE_X6Y142_B5Q;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_AX = CLBLL_L_X4Y142_SLICE_X5Y142_CO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B1 = CLBLL_L_X4Y142_SLICE_X5Y142_DO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B2 = CLBLL_L_X4Y142_SLICE_X5Y142_BQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B4 = CLBLM_R_X5Y141_SLICE_X7Y141_AO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B5 = CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_B6 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C1 = CLBLL_L_X4Y141_SLICE_X5Y141_AQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C2 = CLBLM_R_X5Y141_SLICE_X7Y141_AO6;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C3 = CLBLL_L_X4Y140_SLICE_X4Y140_BO5;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C4 = CLBLL_L_X4Y142_SLICE_X5Y142_A5Q;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_C6 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A3 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D3 = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D4 = CLBLL_L_X4Y142_SLICE_X5Y142_A5Q;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D5 = CLBLM_R_X5Y141_SLICE_X6Y141_DQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D6 = CLBLM_R_X5Y142_SLICE_X6Y142_CQ;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_A6 = 1'b1;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D1 = CLBLM_R_X5Y142_SLICE_X7Y142_AQ;
  assign CLBLL_L_X4Y142_SLICE_X5Y142_D2 = CLBLL_L_X4Y140_SLICE_X4Y140_CO5;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A3 = CLBLM_L_X8Y136_SLICE_X11Y136_AQ;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A4 = CLBLM_L_X8Y137_SLICE_X11Y137_BQ;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A5 = CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_A6 = CLBLM_L_X10Y140_SLICE_X12Y140_CQ;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B3 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_B6 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B6 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C3 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_C6 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_B5 = CLBLM_L_X8Y137_SLICE_X11Y137_AQ;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C5 = CLBLM_R_X7Y134_SLICE_X8Y134_A5Q;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C1 = CLBLM_L_X12Y132_SLICE_X16Y132_BO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_C2 = CLBLM_R_X3Y135_SLICE_X3Y135_A5Q;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D1 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D2 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D3 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D4 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D5 = 1'b1;
  assign CLBLL_L_X2Y75_SLICE_X1Y75_D6 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D1 = CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D2 = CLBLM_L_X8Y135_SLICE_X10Y135_BQ;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D3 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D4 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D5 = CLBLM_R_X11Y133_SLICE_X15Y133_AO6;
  assign CLBLM_L_X8Y136_SLICE_X11Y136_D6 = CLBLM_L_X12Y132_SLICE_X16Y132_BO6;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_D1 = CLBLM_R_X103Y178_SLICE_X163Y178_AO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A1 = CLBLM_R_X3Y136_SLICE_X3Y136_AQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A2 = CLBLM_L_X8Y137_SLICE_X11Y137_BQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A3 = CLBLL_L_X4Y136_SLICE_X5Y136_AQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A4 = CLBLM_L_X8Y139_SLICE_X11Y139_BQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A5 = CLBLM_L_X8Y136_SLICE_X11Y136_AQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_A6 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_T1 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D2 = CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_AX = CLBLM_L_X10Y135_SLICE_X12Y135_BQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B1 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B2 = CLBLM_R_X11Y132_SLICE_X15Y132_AO5;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B3 = CLBLM_R_X3Y136_SLICE_X3Y136_BQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B4 = CLBLM_R_X7Y136_SLICE_X8Y136_B5Q;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B5 = CLBLL_L_X4Y139_SLICE_X5Y139_BQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_B6 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C3 = CLBLM_R_X7Y140_SLICE_X8Y140_CQ;
  assign LIOB33_X0Y127_IOB_X0Y128_O = CLBLM_L_X10Y130_SLICE_X12Y130_CQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C4 = CLBLM_R_X5Y133_SLICE_X6Y133_A5Q;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_BX = CLBLM_L_X10Y132_SLICE_X12Y132_CQ;
  assign LIOB33_X0Y127_IOB_X0Y127_O = CLBLM_L_X10Y140_SLICE_X13Y140_D5Q;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C1 = CLBLM_L_X8Y131_SLICE_X11Y131_CQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C2 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C3 = CLBLM_R_X11Y133_SLICE_X15Y133_AO6;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C4 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C5 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_C6 = CLBLM_R_X7Y137_SLICE_X8Y137_BQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D5 = CLBLM_R_X5Y138_SLICE_X7Y138_BO5;
  assign CLBLM_R_X5Y140_SLICE_X7Y140_D6 = CLBLM_R_X5Y134_SLICE_X6Y134_DQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C6 = CLBLM_L_X10Y138_SLICE_X13Y138_BQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D1 = CLBLM_L_X8Y136_SLICE_X11Y136_AQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D2 = CLBLM_L_X10Y136_SLICE_X12Y136_C5Q;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D3 = CLBLM_L_X8Y137_SLICE_X11Y137_BQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D4 = CLBLM_R_X7Y133_SLICE_X9Y133_CQ;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D5 = 1'b1;
  assign CLBLM_L_X8Y136_SLICE_X10Y136_D6 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A1 = CLBLM_R_X11Y139_SLICE_X14Y139_AO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A2 = CLBLM_R_X7Y133_SLICE_X9Y133_B5Q;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A3 = CLBLM_R_X11Y140_SLICE_X15Y140_AQ;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A5 = CLBLM_R_X11Y140_SLICE_X14Y140_BO5;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_A6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D1 = CLBLM_R_X5Y136_SLICE_X7Y136_AQ;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B1 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B2 = CLBLM_R_X11Y139_SLICE_X15Y139_BO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B3 = CLBLL_L_X4Y130_SLICE_X5Y130_BQ;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B5 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_B6 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A1 = CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A2 = CLBLM_R_X7Y135_SLICE_X9Y135_C5Q;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A3 = CLBLM_R_X7Y130_SLICE_X9Y130_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A5 = CLBLM_R_X7Y133_SLICE_X8Y133_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_A6 = CLBLM_L_X10Y130_SLICE_X12Y130_C5Q;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D5 = CLBLL_L_X4Y138_SLICE_X5Y138_A5Q;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C1 = CLBLM_R_X11Y139_SLICE_X14Y139_AQ;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_C2 = CLBLM_R_X7Y135_SLICE_X8Y135_BQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B1 = CLBLL_L_X4Y137_SLICE_X5Y137_C5Q;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B2 = CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B3 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B4 = CLBLM_R_X5Y130_SLICE_X7Y130_DQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_B6 = CLBLM_R_X7Y131_SLICE_X8Y131_CQ;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D1 = CLBLM_R_X11Y140_SLICE_X14Y140_AQ;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C1 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C2 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C3 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C4 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C5 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_C6 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D3 = CLBLM_L_X12Y140_SLICE_X16Y140_AO6;
  assign CLBLM_R_X11Y140_SLICE_X15Y140_D4 = CLBLM_L_X12Y136_SLICE_X17Y136_BO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A1 = CLBLM_L_X8Y137_SLICE_X11Y137_DQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A2 = CLBLM_L_X10Y139_SLICE_X13Y139_A5Q;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A4 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A5 = CLBLM_R_X11Y139_SLICE_X14Y139_CO6;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D1 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D2 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D3 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D4 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D5 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X9Y130_D6 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_A6 = 1'b1;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_AX = CLBLM_L_X10Y137_SLICE_X12Y137_AQ;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B1 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B3 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X11Y140_SLICE_X14Y140_B4 = CLBLM_L_X10Y138_SLICE_X13Y138_BQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A1 = CLBLL_L_X4Y136_SLICE_X4Y136_A5Q;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A2 = CLBLM_L_X10Y135_SLICE_X12Y135_A5Q;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A1 = CLBLM_R_X5Y141_SLICE_X6Y141_CQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A2 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A3 = CLBLL_L_X4Y136_SLICE_X5Y136_CQ;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A4 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A5 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_A6 = 1'b1;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_B6 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A3 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B1 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B2 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B3 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B4 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B5 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_B6 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B2 = CLBLM_R_X7Y130_SLICE_X8Y130_BQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B3 = CLBLM_R_X5Y131_SLICE_X7Y131_CQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_B4 = CLBLM_R_X7Y130_SLICE_X8Y130_DO6;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C1 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C2 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C3 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C4 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C5 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_C6 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C1 = CLBLM_R_X7Y134_SLICE_X9Y134_BQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C2 = CLBLM_R_X7Y138_SLICE_X8Y138_CQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C3 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C4 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C5 = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_C6 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D1 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D2 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D3 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D4 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D5 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X4Y143_D6 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D1 = CLBLM_R_X7Y134_SLICE_X9Y134_BQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D2 = CLBLM_R_X7Y130_SLICE_X8Y130_AQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C4 = 1'b1;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D3 = CLBLM_R_X5Y131_SLICE_X7Y131_BQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D4 = CLBLM_R_X7Y138_SLICE_X8Y138_CQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D5 = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign CLBLM_R_X7Y130_SLICE_X8Y130_D6 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_D = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_R_X5Y140_SLICE_X6Y140_C6 = CLBLM_R_X5Y141_SLICE_X6Y141_BQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A2 = CLBLM_R_X5Y141_SLICE_X7Y141_AO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A3 = CLBLL_L_X4Y143_SLICE_X5Y143_AQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A4 = CLBLL_L_X4Y143_SLICE_X5Y143_BO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A5 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_A6 = CLBLM_R_X7Y140_SLICE_X9Y140_CQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B1 = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B2 = CLBLM_R_X5Y142_SLICE_X6Y142_CQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B3 = CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B4 = CLBLL_L_X4Y142_SLICE_X5Y142_BQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B5 = CLBLM_R_X5Y142_SLICE_X7Y142_BO6;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C1 = CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C2 = CLBLM_R_X5Y142_SLICE_X6Y142_CQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C3 = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C4 = CLBLL_L_X4Y142_SLICE_X5Y142_BQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C5 = CLBLL_L_X4Y143_SLICE_X5Y143_AQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_C6 = CLBLM_R_X5Y142_SLICE_X7Y142_BO6;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D1 = CLBLL_L_X4Y142_SLICE_X4Y142_AQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D2 = CLBLM_R_X5Y142_SLICE_X6Y142_CQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D3 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D4 = 1'b1;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D5 = CLBLL_L_X4Y143_SLICE_X5Y143_AQ;
  assign CLBLL_L_X4Y143_SLICE_X5Y143_D6 = CLBLL_L_X4Y142_SLICE_X5Y142_BQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A2 = CLBLM_L_X8Y138_SLICE_X10Y138_C5Q;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A3 = CLBLM_L_X8Y137_SLICE_X11Y137_AQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A4 = CLBLM_L_X8Y138_SLICE_X11Y138_CQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A5 = CLBLM_R_X7Y135_SLICE_X9Y135_B5Q;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_D1 = 1'b1;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B1 = CLBLM_R_X7Y138_SLICE_X8Y138_DQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B2 = CLBLM_L_X8Y137_SLICE_X11Y137_BQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B3 = CLBLM_L_X8Y136_SLICE_X10Y136_AO5;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B4 = CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B5 = 1'b1;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C1 = 1'b1;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C2 = CLBLM_L_X8Y137_SLICE_X11Y137_CQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C3 = CLBLM_R_X7Y140_SLICE_X9Y140_AQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C4 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C5 = CLBLM_R_X3Y136_SLICE_X2Y136_DQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D1 = CLBLM_R_X5Y134_SLICE_X7Y134_AQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D3 = CLBLM_R_X7Y142_SLICE_X9Y142_AQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D4 = CLBLL_L_X4Y131_SLICE_X5Y131_B5Q;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D5 = CLBLM_R_X5Y131_SLICE_X6Y131_AQ;
  assign CLBLM_L_X8Y137_SLICE_X11Y137_D6 = 1'b1;
  assign LIOB33_X0Y129_IOB_X0Y129_O = CLBLM_R_X3Y132_SLICE_X3Y132_BQ;
  assign LIOB33_X0Y129_IOB_X0Y130_O = CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A2 = CLBLM_L_X8Y135_SLICE_X10Y135_D5Q;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A3 = CLBLM_L_X8Y137_SLICE_X10Y137_AQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A4 = CLBLM_L_X10Y140_SLICE_X13Y140_D5Q;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A5 = CLBLM_R_X7Y131_SLICE_X9Y131_D5Q;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_A6 = CLBLM_R_X5Y139_SLICE_X7Y139_CQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B1 = CLBLM_R_X3Y135_SLICE_X3Y135_DQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B2 = CLBLM_L_X10Y140_SLICE_X13Y140_BQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B3 = CLBLM_R_X7Y140_SLICE_X8Y140_AQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B5 = CLBLM_R_X7Y132_SLICE_X9Y132_AQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_B6 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_T1 = 1'b1;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C1 = CLBLM_R_X3Y135_SLICE_X2Y135_AQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C2 = CLBLM_R_X7Y137_SLICE_X8Y137_BQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C3 = CLBLM_R_X11Y140_SLICE_X15Y140_B5Q;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C5 = CLBLM_L_X8Y137_SLICE_X11Y137_D5Q;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_C6 = 1'b1;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D1 = CLBLM_L_X8Y132_SLICE_X10Y132_BQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D2 = CLBLL_L_X4Y139_SLICE_X5Y139_CQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D3 = CLBLM_R_X5Y126_SLICE_X6Y126_A5Q;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D4 = CLBLM_L_X10Y137_SLICE_X12Y137_BQ;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y137_SLICE_X10Y137_D6 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A1 = CLBLM_R_X11Y140_SLICE_X14Y140_BO5;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A2 = CLBLM_R_X11Y140_SLICE_X14Y140_BQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A4 = CLBLM_L_X10Y138_SLICE_X13Y138_BQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A5 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_A6 = CLBLM_R_X11Y141_SLICE_X15Y141_AQ;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_D1 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B1 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B2 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B3 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B4 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B5 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_B6 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A1 = CLBLM_R_X7Y135_SLICE_X9Y135_B5Q;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A2 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A3 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A4 = CLBLM_L_X8Y133_SLICE_X11Y133_AQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_A6 = CLBLM_R_X5Y133_SLICE_X6Y133_A5Q;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C2 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C3 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_C4 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B1 = CLBLL_L_X4Y138_SLICE_X4Y138_BQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B2 = CLBLM_L_X10Y140_SLICE_X13Y140_D5Q;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B3 = CLBLL_L_X4Y129_SLICE_X4Y129_AQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B4 = CLBLM_R_X7Y131_SLICE_X9Y131_D5Q;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_B6 = CLBLM_R_X7Y131_SLICE_X9Y131_BQ;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D1 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C1 = CLBLM_R_X7Y129_SLICE_X8Y129_AQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C3 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C4 = CLBLM_R_X5Y130_SLICE_X7Y130_BQ;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_C6 = CLBLL_L_X4Y138_SLICE_X5Y138_D5Q;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D3 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X15Y141_D4 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A1 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A2 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A3 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A4 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A5 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D2 = CLBLM_L_X10Y140_SLICE_X13Y140_D5Q;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D3 = CLBLM_R_X5Y131_SLICE_X7Y131_D5Q;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D4 = CLBLL_L_X4Y137_SLICE_X5Y137_C5Q;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D5 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X9Y131_D6 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_A6 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_AX = CLBLM_R_X11Y140_SLICE_X14Y140_AO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B1 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B2 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B3 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_B4 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A1 = CLBLM_R_X7Y131_SLICE_X8Y131_BO5;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A3 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A4 = CLBLM_R_X5Y130_SLICE_X6Y130_B5Q;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A5 = CLBLM_L_X8Y130_SLICE_X10Y130_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_A6 = CLBLM_R_X5Y130_SLICE_X7Y130_BQ;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C1 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C2 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_AX = CLBLM_R_X7Y131_SLICE_X8Y131_BO6;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_C3 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B1 = CLBLL_L_X4Y134_SLICE_X4Y134_CQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B2 = CLBLM_R_X7Y136_SLICE_X8Y136_BQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B4 = CLBLM_R_X5Y130_SLICE_X6Y130_B5Q;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B5 = CLBLM_R_X7Y131_SLICE_X8Y131_A5Q;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_B6 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D1 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D2 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C2 = CLBLM_R_X7Y131_SLICE_X8Y131_CQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C3 = CLBLM_R_X7Y132_SLICE_X8Y132_D5Q;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C5 = CLBLM_L_X8Y131_SLICE_X10Y131_AQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_C6 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D3 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D4 = 1'b1;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D5 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y141_SLICE_X14Y141_D6 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D2 = 1'b1;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D3 = CLBLM_R_X7Y131_SLICE_X8Y131_DQ;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D4 = CLBLM_R_X13Y134_SLICE_X18Y134_AO6;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D5 = CLBLM_R_X7Y134_SLICE_X8Y134_A5Q;
  assign CLBLM_R_X7Y131_SLICE_X8Y131_D6 = CLBLM_R_X5Y142_SLICE_X6Y142_AQ;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A2 = CLBLM_L_X8Y138_SLICE_X10Y138_D5Q;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A3 = CLBLM_L_X8Y138_SLICE_X11Y138_AQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A4 = CLBLM_L_X8Y141_SLICE_X11Y141_BQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A5 = CLBLM_L_X8Y130_SLICE_X11Y130_AO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_A6 = CLBLM_R_X5Y133_SLICE_X6Y133_A5Q;
  assign LIOB33_X0Y131_IOB_X0Y131_O = CLBLL_L_X2Y75_SLICE_X0Y75_AO6;
  assign LIOB33_X0Y131_IOB_X0Y132_O = CLBLM_R_X3Y131_SLICE_X2Y131_AO6;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B2 = CLBLM_L_X8Y138_SLICE_X10Y138_D5Q;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B3 = CLBLM_R_X7Y132_SLICE_X8Y132_BQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B4 = CLBLM_L_X8Y138_SLICE_X11Y138_BQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B5 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_B6 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C1 = CLBLM_L_X8Y137_SLICE_X11Y137_AQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C2 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C3 = CLBLM_R_X5Y137_SLICE_X7Y137_BQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C5 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_C6 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D1 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D2 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D3 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D4 = CLBLM_R_X3Y137_SLICE_X3Y137_B5Q;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D5 = CLBLM_L_X8Y138_SLICE_X11Y138_B5Q;
  assign CLBLM_L_X8Y138_SLICE_X11Y138_D6 = CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A2 = CLBLM_L_X8Y137_SLICE_X10Y137_D5Q;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A3 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A4 = CLBLM_R_X7Y137_SLICE_X9Y137_BQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A5 = CLBLM_R_X11Y142_SLICE_X14Y142_AQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_A6 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B2 = CLBLL_L_X4Y138_SLICE_X5Y138_D5Q;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B3 = CLBLM_L_X12Y136_SLICE_X16Y136_AQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B4 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B5 = CLBLM_L_X8Y139_SLICE_X10Y139_AQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_B6 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C1 = CLBLL_L_X4Y138_SLICE_X5Y138_C5Q;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C2 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C4 = CLBLM_L_X10Y140_SLICE_X13Y140_BQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_C6 = 1'b1;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D1 = CLBLM_L_X10Y140_SLICE_X12Y140_DQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D2 = CLBLL_L_X4Y135_SLICE_X5Y135_BQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D4 = CLBLM_L_X8Y137_SLICE_X10Y137_D5Q;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D5 = CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  assign CLBLM_L_X8Y138_SLICE_X10Y138_D6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_D1 = CLBLL_L_X4Y141_SLICE_X5Y141_DO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A2 = CLBLL_L_X4Y138_SLICE_X4Y138_AQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A3 = CLBLM_R_X11Y136_SLICE_X15Y136_BO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A4 = CLBLM_L_X10Y139_SLICE_X13Y139_A5Q;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A5 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_A6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_T1 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_D1 = CLBLM_L_X12Y142_SLICE_X16Y142_AO6;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B1 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B2 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B3 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B4 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B5 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_B6 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_D1 = CLBLL_L_X4Y139_SLICE_X5Y139_DO5;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_T1 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A1 = CLBLM_L_X8Y133_SLICE_X11Y133_A5Q;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A2 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A4 = CLBLM_R_X5Y133_SLICE_X6Y133_AQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A5 = CLBLM_R_X11Y142_SLICE_X14Y142_AQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_A6 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C1 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C2 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_C3 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B1 = CLBLM_R_X7Y135_SLICE_X9Y135_D5Q;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B2 = CLBLM_R_X7Y132_SLICE_X9Y132_BQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B4 = CLBLM_L_X10Y140_SLICE_X13Y140_D5Q;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B5 = CLBLM_R_X7Y131_SLICE_X9Y131_D5Q;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_B6 = CLBLM_R_X7Y134_SLICE_X8Y134_BQ;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D1 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D2 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C2 = CLBLM_R_X7Y133_SLICE_X9Y133_AQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C3 = CLBLM_R_X7Y132_SLICE_X9Y132_BQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C4 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C5 = CLBLM_R_X7Y132_SLICE_X9Y132_CQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_C6 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D3 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X15Y142_D4 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A1 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A2 = CLBLM_R_X11Y137_SLICE_X14Y137_AO6;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A5 = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D1 = CLBLM_R_X7Y133_SLICE_X8Y133_C5Q;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D2 = CLBLL_L_X4Y134_SLICE_X4Y134_C5Q;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D3 = CLBLM_R_X7Y131_SLICE_X9Y131_DQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_A6 = CLBLM_R_X7Y138_SLICE_X9Y138_CQ;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D5 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X9Y132_D6 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_A6 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B1 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B2 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_B3 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A1 = CLBLM_R_X7Y133_SLICE_X9Y133_B5Q;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A2 = CLBLM_R_X7Y135_SLICE_X9Y135_C5Q;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A3 = CLBLM_R_X7Y132_SLICE_X8Y132_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A4 = CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_A6 = CLBLM_L_X8Y138_SLICE_X10Y138_CQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C1 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_C2 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B2 = CLBLL_L_X4Y132_SLICE_X4Y132_CQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B4 = CLBLM_R_X7Y135_SLICE_X9Y135_B5Q;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B5 = CLBLM_R_X7Y133_SLICE_X8Y133_C5Q;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_B6 = CLBLM_R_X7Y132_SLICE_X8Y132_BQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D1 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D2 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C2 = CLBLM_R_X7Y132_SLICE_X8Y132_CQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C3 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C4 = 1'b1;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C5 = CLBLM_L_X8Y133_SLICE_X10Y133_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_C6 = CLBLM_R_X3Y132_SLICE_X2Y132_BQ;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D5 = 1'b1;
  assign CLBLM_R_X11Y142_SLICE_X14Y142_D6 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B4 = CLBLM_L_X10Y140_SLICE_X13Y140_CQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D1 = CLBLM_R_X3Y131_SLICE_X2Y131_AQ;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D3 = CLBLM_R_X7Y131_SLICE_X9Y131_BQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_B6 = CLBLM_L_X10Y139_SLICE_X13Y139_A5Q;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D4 = CLBLM_R_X7Y137_SLICE_X9Y137_D5Q;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D5 = CLBLM_R_X7Y132_SLICE_X9Y132_D5Q;
  assign CLBLM_R_X7Y132_SLICE_X8Y132_D6 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C1 = CLBLM_R_X5Y140_SLICE_X7Y140_A5Q;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C2 = CLBLM_L_X10Y141_SLICE_X13Y141_CQ;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C3 = CLBLM_L_X10Y136_SLICE_X12Y136_C5Q;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C5 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_C6 = CLBLM_R_X7Y142_SLICE_X9Y142_DO5;
  assign LIOB33_X0Y133_IOB_X0Y134_O = CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  assign LIOB33_X0Y133_IOB_X0Y133_O = CLBLL_L_X4Y133_SLICE_X4Y133_BO5;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A2 = CLBLM_R_X11Y131_SLICE_X14Y131_BO6;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A3 = CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A4 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A5 = CLBLM_R_X5Y140_SLICE_X6Y140_AQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_A6 = CLBLM_L_X10Y140_SLICE_X13Y140_B5Q;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B1 = CLBLM_L_X8Y140_SLICE_X11Y140_B5Q;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B2 = CLBLM_L_X8Y139_SLICE_X11Y139_BQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B3 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B4 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B5 = CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C1 = CLBLM_L_X8Y138_SLICE_X11Y138_C5Q;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C2 = CLBLM_L_X8Y139_SLICE_X11Y139_CQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C3 = CLBLM_L_X10Y140_SLICE_X13Y140_BQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C4 = CLBLM_R_X5Y137_SLICE_X7Y137_BQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_C6 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D1 = CLBLM_R_X5Y140_SLICE_X7Y140_A5Q;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D3 = CLBLM_L_X10Y141_SLICE_X12Y141_DO6;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_D = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D1 = CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D2 = CLBLM_R_X11Y141_SLICE_X14Y141_AQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D3 = CLBLM_L_X10Y140_SLICE_X13Y140_C5Q;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D4 = CLBLM_L_X10Y140_SLICE_X13Y140_B5Q;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D5 = CLBLL_L_X4Y133_SLICE_X4Y133_AQ;
  assign CLBLM_L_X8Y139_SLICE_X11Y139_D6 = CLBLM_L_X10Y139_SLICE_X12Y139_AO5;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D4 = CLBLM_L_X10Y141_SLICE_X12Y141_DO5;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D5 = CLBLM_L_X8Y140_SLICE_X10Y140_CQ;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_D = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_L_X10Y141_SLICE_X13Y141_D6 = CLBLM_L_X10Y141_SLICE_X13Y141_DQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A1 = CLBLM_L_X8Y140_SLICE_X11Y140_B5Q;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A2 = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A3 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A4 = CLBLM_L_X8Y141_SLICE_X11Y141_BQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A5 = CLBLM_R_X5Y137_SLICE_X7Y137_B5Q;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_A6 = CLBLM_R_X7Y133_SLICE_X8Y133_A5Q;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_AX = CLBLM_R_X7Y133_SLICE_X9Y133_BQ;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B1 = CLBLM_R_X3Y133_SLICE_X3Y133_DO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B2 = CLBLM_L_X8Y144_SLICE_X10Y144_BO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B3 = CLBLM_R_X7Y134_SLICE_X8Y134_DO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B4 = CLBLM_R_X7Y139_SLICE_X8Y139_DO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B5 = CLBLM_R_X7Y139_SLICE_X8Y139_AO5;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_B6 = CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C1 = CLBLM_L_X12Y134_SLICE_X17Y134_AO5;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C2 = CLBLL_L_X4Y130_SLICE_X5Y130_DO5;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C3 = CLBLM_L_X8Y139_SLICE_X11Y139_DO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C4 = CLBLM_R_X7Y139_SLICE_X8Y139_DO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C5 = CLBLM_R_X7Y139_SLICE_X9Y139_CO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_C6 = CLBLM_L_X8Y144_SLICE_X10Y144_BO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A2 = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A4 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_A6 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D1 = CLBLM_L_X10Y133_SLICE_X12Y133_CO6;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D2 = CLBLM_R_X5Y136_SLICE_X6Y136_B5Q;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D3 = CLBLM_L_X8Y137_SLICE_X10Y137_D5Q;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D4 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D5 = 1'b1;
  assign CLBLM_L_X8Y139_SLICE_X10Y139_D6 = CLBLL_L_X4Y134_SLICE_X4Y134_D5Q;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A2 = CLBLM_R_X7Y142_SLICE_X9Y142_DO5;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B3 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A3 = CLBLM_L_X10Y141_SLICE_X12Y141_AQ;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_B6 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C2 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A4 = CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_C6 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_A5 = CLBLM_R_X5Y140_SLICE_X7Y140_A5Q;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X163Y178_D6 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_A6 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B3 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_B6 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C1 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C2 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C3 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A1 = CLBLM_R_X5Y133_SLICE_X7Y133_DQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A2 = CLBLM_R_X7Y138_SLICE_X8Y138_AQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A4 = CLBLM_L_X8Y135_SLICE_X10Y135_BQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A5 = CLBLM_L_X10Y140_SLICE_X13Y140_B5Q;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_A6 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C4 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C5 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_C6 = 1'b1;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B4 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B2 = CLBLM_R_X3Y131_SLICE_X3Y131_AQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B4 = CLBLM_L_X8Y135_SLICE_X10Y135_BQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B5 = CLBLL_L_X4Y131_SLICE_X5Y131_B5Q;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B5 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B6 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_B1 = CLBLM_R_X5Y134_SLICE_X6Y134_CQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_B6 = CLBLM_L_X10Y140_SLICE_X12Y140_CQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C2 = CLBLM_R_X3Y134_SLICE_X3Y134_A5Q;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C3 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C4 = CLBLM_R_X7Y134_SLICE_X8Y134_BQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C5 = CLBLM_L_X10Y140_SLICE_X13Y140_BQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_C6 = 1'b1;
  assign CLBLM_R_X103Y178_SLICE_X162Y178_D6 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D2 = CLBLM_R_X5Y133_SLICE_X7Y133_CQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D3 = CLBLM_L_X8Y136_SLICE_X11Y136_B5Q;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D4 = CLBLM_R_X7Y136_SLICE_X9Y136_AQ;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D5 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X9Y133_D6 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A1 = CLBLM_R_X7Y134_SLICE_X9Y134_DQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A2 = CLBLM_R_X7Y141_SLICE_X8Y141_AQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A4 = CLBLL_L_X4Y133_SLICE_X4Y133_A5Q;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A5 = CLBLM_R_X5Y130_SLICE_X7Y130_BQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_A6 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B1 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B2 = CLBLM_R_X7Y133_SLICE_X8Y133_BQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B3 = CLBLM_R_X7Y141_SLICE_X8Y141_AQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B4 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_B6 = CLBLM_R_X7Y132_SLICE_X8Y132_DQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C1 = CLBLM_L_X8Y141_SLICE_X11Y141_AQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C5 = CLBLM_L_X10Y140_SLICE_X13Y140_C5Q;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C2 = CLBLL_L_X4Y137_SLICE_X5Y137_C5Q;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C5 = CLBLM_R_X7Y136_SLICE_X8Y136_DQ;
  assign CLBLM_L_X10Y141_SLICE_X12Y141_C6 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_C6 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D1 = CLBLM_R_X7Y132_SLICE_X9Y132_D5Q;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D2 = CLBLM_L_X12Y136_SLICE_X16Y136_AQ;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D4 = CLBLM_R_X5Y132_SLICE_X7Y132_C5Q;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D5 = 1'b1;
  assign CLBLM_R_X7Y133_SLICE_X8Y133_D6 = 1'b1;
  assign LIOB33_X0Y135_IOB_X0Y136_O = CLBLM_L_X8Y141_SLICE_X11Y141_BQ;
  assign LIOB33_X0Y135_IOB_X0Y135_O = CLBLM_R_X3Y132_SLICE_X3Y132_AQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A1 = CLBLM_L_X8Y141_SLICE_X10Y141_BQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A2 = CLBLM_R_X5Y133_SLICE_X7Y133_AQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A3 = CLBLM_L_X8Y140_SLICE_X11Y140_AQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A5 = CLBLL_L_X4Y135_SLICE_X4Y135_D5Q;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_A6 = CLBLM_L_X8Y139_SLICE_X11Y139_CQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B1 = CLBLM_R_X3Y134_SLICE_X2Y134_CO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B2 = CLBLM_L_X10Y140_SLICE_X12Y140_BQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B3 = CLBLM_R_X7Y137_SLICE_X8Y137_CQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B5 = CLBLM_L_X8Y141_SLICE_X11Y141_CO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_B6 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C2 = CLBLM_L_X8Y140_SLICE_X11Y140_CQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C3 = CLBLM_R_X13Y134_SLICE_X18Y134_AO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C4 = CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C5 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_C6 = CLBLM_R_X7Y140_SLICE_X9Y140_CQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D1 = CLBLM_L_X10Y141_SLICE_X12Y141_BQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D2 = CLBLM_R_X7Y140_SLICE_X9Y140_D5Q;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D3 = CLBLM_L_X8Y141_SLICE_X10Y141_DO6;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D4 = CLBLM_L_X8Y134_SLICE_X11Y134_BQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D5 = CLBLM_L_X10Y140_SLICE_X12Y140_CQ;
  assign CLBLM_L_X8Y140_SLICE_X11Y140_D6 = CLBLM_R_X7Y136_SLICE_X8Y136_D5Q;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_T1 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A1 = CLBLM_R_X5Y140_SLICE_X6Y140_CQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A3 = CLBLM_L_X8Y140_SLICE_X10Y140_AQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A4 = CLBLL_L_X4Y136_SLICE_X4Y136_D5Q;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A5 = CLBLM_R_X7Y140_SLICE_X8Y140_BQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_A6 = CLBLM_L_X8Y138_SLICE_X10Y138_CQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B1 = CLBLL_L_X4Y136_SLICE_X4Y136_D5Q;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B2 = CLBLM_L_X8Y140_SLICE_X10Y140_BQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B3 = CLBLM_L_X8Y138_SLICE_X10Y138_AQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B4 = CLBLM_L_X8Y140_SLICE_X10Y140_D5Q;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_B6 = CLBLM_L_X8Y138_SLICE_X10Y138_CQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C6 = CLBLL_L_X4Y140_SLICE_X4Y140_CO5;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C1 = CLBLM_R_X7Y140_SLICE_X8Y140_BQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C2 = CLBLM_L_X8Y142_SLICE_X10Y142_A5Q;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C3 = CLBLM_L_X10Y141_SLICE_X13Y141_DQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C5 = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_C6 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D1 = CLBLM_L_X10Y139_SLICE_X12Y139_AQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D2 = CLBLM_R_X5Y140_SLICE_X6Y140_CQ;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D3 = CLBLM_R_X5Y140_SLICE_X6Y140_A5Q;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D5 = 1'b1;
  assign CLBLM_L_X8Y140_SLICE_X10Y140_D6 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_D1 = CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C4 = CLBLM_R_X7Y140_SLICE_X9Y140_DQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C5 = CLBLM_R_X3Y133_SLICE_X3Y133_DO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A1 = CLBLM_R_X7Y133_SLICE_X8Y133_AQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A2 = CLBLL_L_X4Y135_SLICE_X4Y135_D5Q;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A4 = CLBLM_R_X7Y134_SLICE_X9Y134_AQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A5 = CLBLM_R_X5Y133_SLICE_X7Y133_AQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_A6 = CLBLM_R_X7Y138_SLICE_X9Y138_CQ;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_C6 = CLBLM_R_X7Y135_SLICE_X9Y135_DQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B1 = CLBLM_L_X8Y134_SLICE_X11Y134_B5Q;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B2 = CLBLM_R_X7Y134_SLICE_X8Y134_DO5;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B4 = CLBLM_R_X5Y133_SLICE_X6Y133_A5Q;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B5 = CLBLM_R_X7Y140_SLICE_X9Y140_D5Q;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_B6 = CLBLM_R_X7Y134_SLICE_X9Y134_BQ;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_T1 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C1 = CLBLM_R_X7Y138_SLICE_X8Y138_AQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C2 = CLBLM_R_X7Y134_SLICE_X9Y134_CQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C4 = CLBLM_L_X8Y138_SLICE_X10Y138_CQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C5 = CLBLM_R_X7Y138_SLICE_X9Y138_A5Q;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_C6 = CLBLL_L_X4Y136_SLICE_X4Y136_D5Q;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D2 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D3 = CLBLM_R_X7Y134_SLICE_X9Y134_DQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D4 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D5 = CLBLL_L_X4Y134_SLICE_X4Y134_AQ;
  assign CLBLM_R_X7Y134_SLICE_X9Y134_D6 = CLBLM_R_X7Y134_SLICE_X9Y134_AQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A1 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A2 = CLBLL_L_X4Y135_SLICE_X4Y135_BQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A3 = CLBLM_L_X8Y136_SLICE_X10Y136_BQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A4 = CLBLM_L_X12Y136_SLICE_X16Y136_AQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_A6 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B1 = CLBLM_R_X7Y136_SLICE_X8Y136_B5Q;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B2 = CLBLM_R_X5Y134_SLICE_X7Y134_BQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B4 = CLBLM_R_X7Y134_SLICE_X9Y134_BQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B5 = CLBLM_R_X5Y134_SLICE_X6Y134_CQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_B6 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D2 = CLBLM_R_X7Y138_SLICE_X9Y138_DO6;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D3 = CLBLL_L_X4Y138_SLICE_X4Y138_CO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C1 = CLBLM_R_X7Y133_SLICE_X9Y133_D5Q;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C2 = CLBLL_L_X2Y138_SLICE_X1Y138_BO6;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C3 = CLBLL_L_X4Y135_SLICE_X4Y135_DQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C4 = CLBLM_R_X7Y140_SLICE_X9Y140_BQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_C6 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D5 = CLBLM_L_X10Y141_SLICE_X13Y141_BQ;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_D = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B5 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X9Y139_D6 = 1'b1;
  assign LIOB33_X0Y137_IOB_X0Y137_O = CLBLM_R_X7Y137_SLICE_X9Y137_D5Q;
  assign LIOB33_X0Y137_IOB_X0Y138_O = CLBLM_R_X3Y139_SLICE_X3Y139_A5Q;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_D1 = CLBLM_R_X5Y133_SLICE_X7Y133_A5Q;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D1 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D2 = CLBLM_R_X7Y134_SLICE_X9Y134_BQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D3 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D4 = CLBLM_R_X7Y138_SLICE_X8Y138_CQ;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D5 = 1'b1;
  assign CLBLM_R_X7Y134_SLICE_X8Y134_D6 = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_T1 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_D1 = CLBLM_L_X12Y142_SLICE_X16Y142_AO5;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_B6 = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_D1 = CLBLM_R_X3Y132_SLICE_X3Y132_BQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_T1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A2 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A3 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A4 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A5 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_A6 = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_T1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B2 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B3 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B4 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B5 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_B6 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_D1 = CLBLM_L_X12Y143_SLICE_X16Y143_AO6;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C2 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C3 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C4 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C5 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_C6 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D1 = CLBLM_R_X11Y141_SLICE_X14Y141_AQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_T1 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D2 = CLBLL_L_X4Y134_SLICE_X4Y134_C5Q;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_T1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D2 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D3 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D4 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D5 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X0Y133_D6 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D3 = CLBLM_L_X10Y140_SLICE_X13Y140_BQ;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D4 = CLBLM_L_X12Y136_SLICE_X16Y136_A5Q;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D5 = 1'b1;
  assign CLBLM_R_X11Y137_SLICE_X14Y137_D6 = CLBLM_L_X10Y136_SLICE_X13Y136_CO6;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1 = 1'b1;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B5 = CLBLM_L_X10Y136_SLICE_X12Y136_BQ;
  assign CLBLM_L_X8Y133_SLICE_X11Y133_B6 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A1 = CLBLM_L_X8Y141_SLICE_X11Y141_AQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A3 = CLBLM_R_X5Y140_SLICE_X7Y140_A5Q;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A5 = CLBLM_R_X11Y140_SLICE_X14Y140_AQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A6 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_A2 = CLBLM_L_X10Y134_SLICE_X12Y134_AQ;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C4 = CLBLL_L_X4Y142_SLICE_X5Y142_A5Q;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_C5 = CLBLM_R_X5Y141_SLICE_X6Y141_DQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B1 = CLBLM_L_X8Y141_SLICE_X11Y141_DO6;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B5 = CLBLM_L_X8Y141_SLICE_X11Y141_CO5;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B6 = CLBLM_L_X10Y141_SLICE_X12Y141_CQ;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A4 = CLBLM_R_X3Y133_SLICE_X2Y133_AQ;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_A6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B2 = CLBLM_L_X8Y141_SLICE_X11Y141_BQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_B3 = CLBLM_R_X5Y132_SLICE_X6Y132_AQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C3 = CLBLM_L_X8Y140_SLICE_X11Y140_B5Q;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C4 = CLBLM_L_X8Y141_SLICE_X11Y141_BQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C5 = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_C6 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B2 = CLBLM_R_X7Y134_SLICE_X8Y134_CQ;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B3 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B4 = CLBLM_R_X3Y141_SLICE_X2Y141_CO6;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B5 = CLBLL_L_X4Y138_SLICE_X4Y138_BQ;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_B6 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C2 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C3 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C4 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C5 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_C6 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D1 = CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D2 = CLBLM_L_X8Y141_SLICE_X10Y141_CO6;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D3 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D4 = CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D5 = CLBLM_L_X8Y143_SLICE_X11Y143_AQ;
  assign CLBLM_L_X8Y141_SLICE_X11Y141_D6 = CLBLM_L_X8Y143_SLICE_X10Y143_BO6;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D1 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D2 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D3 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D4 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D5 = 1'b1;
  assign CLBLL_L_X2Y133_SLICE_X1Y133_D6 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A1 = CLBLM_L_X8Y143_SLICE_X10Y143_BO5;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A3 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A4 = CLBLM_R_X5Y134_SLICE_X7Y134_AQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A5 = CLBLM_L_X8Y141_SLICE_X10Y141_CO5;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_A6 = CLBLM_L_X8Y141_SLICE_X10Y141_CO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B2 = CLBLM_L_X8Y141_SLICE_X10Y141_BQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B3 = CLBLM_L_X8Y144_SLICE_X10Y144_AO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B4 = CLBLM_R_X5Y137_SLICE_X7Y137_A5Q;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B5 = CLBLM_L_X8Y141_SLICE_X10Y141_CO5;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_B6 = CLBLM_L_X8Y141_SLICE_X10Y141_CO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C1 = CLBLM_L_X8Y144_SLICE_X10Y144_AO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C2 = CLBLM_L_X8Y141_SLICE_X11Y141_BQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C3 = CLBLM_R_X7Y133_SLICE_X8Y133_A5Q;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C4 = CLBLM_L_X8Y141_SLICE_X10Y141_BQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C5 = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_C6 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C4 = CLBLM_L_X8Y137_SLICE_X10Y137_B5Q;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D5 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C5 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X7Y141_D6 = CLBLL_L_X4Y142_SLICE_X5Y142_A5Q;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D1 = CLBLM_L_X10Y141_SLICE_X13Y141_CQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D2 = CLBLM_R_X7Y142_SLICE_X9Y142_AQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D3 = 1'b1;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D4 = CLBLM_L_X8Y142_SLICE_X10Y142_DO6;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D5 = CLBLM_L_X10Y141_SLICE_X13Y141_DQ;
  assign CLBLM_L_X8Y141_SLICE_X10Y141_D6 = CLBLM_L_X10Y141_SLICE_X12Y141_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_C6 = CLBLM_R_X7Y138_SLICE_X8Y138_BQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D1 = CLBLM_R_X7Y141_SLICE_X8Y141_AQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A1 = CLBLL_L_X4Y138_SLICE_X5Y138_DQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A2 = CLBLM_L_X10Y140_SLICE_X12Y140_D5Q;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A4 = CLBLM_R_X5Y134_SLICE_X6Y134_A5Q;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A5 = CLBLM_R_X3Y135_SLICE_X2Y135_CQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_A6 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D2 = CLBLM_R_X5Y139_SLICE_X6Y139_CQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D3 = CLBLM_R_X7Y135_SLICE_X9Y135_C5Q;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_D = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B1 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B2 = CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B3 = CLBLM_R_X3Y134_SLICE_X2Y134_AQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B4 = CLBLM_R_X7Y130_SLICE_X9Y130_AQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B5 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_B6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D4 = CLBLM_R_X7Y141_SLICE_X9Y141_AQ;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D5 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_BX = CLBLL_L_X4Y135_SLICE_X5Y135_DO5;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C1 = CLBLM_R_X7Y130_SLICE_X9Y130_AQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C4 = CLBLM_R_X7Y140_SLICE_X8Y140_C5Q;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C5 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_C6 = 1'b1;
  assign CLBLM_R_X7Y139_SLICE_X8Y139_D6 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D2 = CLBLM_L_X10Y135_SLICE_X13Y135_AQ;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D3 = CLBLM_R_X5Y142_SLICE_X6Y142_B5Q;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D4 = CLBLL_L_X4Y137_SLICE_X5Y137_C5Q;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D5 = CLBLM_L_X8Y139_SLICE_X11Y139_C5Q;
  assign CLBLM_R_X7Y135_SLICE_X9Y135_D6 = 1'b1;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A1 = CLBLM_R_X7Y136_SLICE_X8Y136_DQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A2 = CLBLL_L_X4Y133_SLICE_X5Y133_DQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A3 = CLBLM_R_X7Y135_SLICE_X9Y135_A5Q;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A4 = CLBLL_L_X4Y135_SLICE_X4Y135_C5Q;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A5 = CLBLM_L_X8Y135_SLICE_X10Y135_DQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_A6 = CLBLM_R_X7Y134_SLICE_X8Y134_B5Q;
  assign LIOB33_X0Y139_IOB_X0Y139_O = CLBLM_R_X3Y139_SLICE_X2Y139_C5Q;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B5 = 1'b1;
  assign LIOB33_X0Y139_IOB_X0Y140_O = CLBLM_R_X3Y137_SLICE_X3Y137_D5Q;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_AX = CLBLM_R_X3Y135_SLICE_X3Y135_BQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B1 = CLBLM_L_X10Y137_SLICE_X13Y137_BO6;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_B6 = CLBLM_R_X5Y142_SLICE_X6Y142_BQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B2 = CLBLM_L_X12Y135_SLICE_X16Y135_AO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B3 = CLBLM_R_X11Y133_SLICE_X14Y133_CO5;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B4 = CLBLL_L_X4Y132_SLICE_X5Y132_D5Q;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B5 = CLBLL_L_X4Y132_SLICE_X5Y132_AQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_B6 = CLBLL_L_X4Y135_SLICE_X4Y135_BQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_BX = CLBLM_R_X7Y134_SLICE_X8Y134_B5Q;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C1 = CLBLM_R_X3Y135_SLICE_X3Y135_AQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C2 = CLBLM_R_X11Y133_SLICE_X14Y133_CO5;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C3 = CLBLM_L_X10Y137_SLICE_X13Y137_BO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C4 = CLBLL_L_X4Y138_SLICE_X5Y138_A5Q;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C5 = CLBLM_L_X12Y135_SLICE_X16Y135_AO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_C6 = CLBLM_R_X7Y135_SLICE_X9Y135_BQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_CE = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D1 = CLBLM_L_X12Y134_SLICE_X17Y134_AO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D2 = CLBLM_R_X7Y132_SLICE_X8Y132_CQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D3 = CLBLM_R_X3Y135_SLICE_X2Y135_BQ;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D4 = CLBLM_R_X11Y131_SLICE_X14Y131_CO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D5 = CLBLM_L_X10Y137_SLICE_X13Y137_BO6;
  assign CLBLM_R_X7Y135_SLICE_X8Y135_D6 = CLBLM_R_X5Y135_SLICE_X7Y135_BQ;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_A1 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_A2 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_A3 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_A4 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_A5 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_A6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C4 = CLBLM_L_X8Y142_SLICE_X10Y142_A5Q;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C5 = CLBLM_R_X5Y141_SLICE_X6Y141_CQ;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_B1 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_B2 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_B3 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_B4 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_B5 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_B6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_C6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_C1 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_C2 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_C3 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_C4 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_C5 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_C6 = 1'b1;
  assign CLBLM_R_X5Y141_SLICE_X6Y141_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_D1 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_D2 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_D3 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_D4 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_D5 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X0Y134_D6 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A1 = CLBLM_L_X8Y138_SLICE_X11Y138_B5Q;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A3 = CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A4 = CLBLM_L_X8Y142_SLICE_X11Y142_AQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A5 = CLBLM_L_X8Y141_SLICE_X10Y141_CO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_A6 = CLBLM_L_X8Y142_SLICE_X11Y142_CO6;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_A2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_A3 = CLBLL_L_X4Y138_SLICE_X4Y138_BQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B1 = CLBLM_L_X8Y143_SLICE_X11Y143_BO6;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B2 = CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B3 = CLBLM_L_X8Y143_SLICE_X11Y143_AQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B4 = CLBLM_L_X10Y135_SLICE_X12Y135_B5Q;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_B1 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_B6 = CLBLM_L_X8Y143_SLICE_X11Y143_CO6;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_A4 = CLBLM_R_X3Y135_SLICE_X2Y135_AQ;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_B4 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C1 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C2 = CLBLM_L_X8Y142_SLICE_X11Y142_AQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C3 = CLBLM_L_X8Y140_SLICE_X11Y140_B5Q;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C4 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C5 = CLBLM_R_X5Y137_SLICE_X7Y137_B5Q;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_C6 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_B3 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_C3 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_C4 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_C5 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_C6 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_C1 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_C2 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D1 = CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D2 = CLBLM_L_X8Y143_SLICE_X11Y143_AQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D3 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D4 = CLBLM_L_X8Y143_SLICE_X10Y143_BO5;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D5 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_L_X8Y142_SLICE_X11Y142_D6 = CLBLM_R_X7Y143_SLICE_X8Y143_A5Q;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_D1 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_D2 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_D3 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_D4 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_D5 = 1'b1;
  assign CLBLL_L_X2Y134_SLICE_X1Y134_D6 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A1 = CLBLM_R_X7Y142_SLICE_X9Y142_CQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A2 = CLBLM_L_X8Y141_SLICE_X11Y141_AO5;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A3 = CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A4 = CLBLM_R_X5Y140_SLICE_X7Y140_A5Q;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_A6 = CLBLM_L_X10Y141_SLICE_X12Y141_C5Q;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_AX = CLBLM_L_X8Y142_SLICE_X10Y142_BO6;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B1 = CLBLM_L_X8Y134_SLICE_X10Y134_A5Q;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B2 = CLBLM_L_X8Y141_SLICE_X11Y141_BQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B3 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B4 = CLBLM_R_X7Y133_SLICE_X8Y133_A5Q;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_B6 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C1 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C2 = CLBLM_L_X10Y134_SLICE_X12Y134_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C3 = CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C4 = CLBLM_L_X8Y141_SLICE_X11Y141_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C5 = CLBLM_R_X7Y142_SLICE_X9Y142_CQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_C6 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D1 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D2 = CLBLM_L_X8Y142_SLICE_X10Y142_AQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D3 = CLBLM_R_X7Y142_SLICE_X9Y142_CQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D4 = CLBLM_R_X7Y142_SLICE_X9Y142_BQ;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D5 = 1'b1;
  assign CLBLM_L_X8Y142_SLICE_X10Y142_D6 = CLBLM_L_X8Y141_SLICE_X11Y141_AQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B5 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A2 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A3 = CLBLM_L_X8Y136_SLICE_X10Y136_AQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A4 = CLBLM_R_X7Y136_SLICE_X9Y136_D5Q;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A5 = CLBLM_R_X11Y142_SLICE_X14Y142_AQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_A6 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B2 = CLBLM_R_X7Y136_SLICE_X9Y136_BQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B3 = CLBLM_R_X7Y134_SLICE_X9Y134_AQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B4 = CLBLM_R_X11Y131_SLICE_X14Y131_BO6;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B5 = CLBLM_R_X7Y136_SLICE_X9Y136_DQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_B6 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B6 = 1'b1;
  assign LIOB33_X0Y141_IOB_X0Y141_O = CLBLL_L_X4Y134_SLICE_X5Y134_DQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A1 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A2 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A3 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A4 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A5 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_A6 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C1 = CLBLM_R_X5Y141_SLICE_X6Y141_AQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C2 = CLBLM_R_X7Y136_SLICE_X9Y136_CQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_C3 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B1 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B2 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B3 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B4 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B5 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_B6 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D1 = CLBLM_R_X7Y138_SLICE_X9Y138_AQ;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C1 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C2 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C3 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C4 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C5 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_C6 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D3 = CLBLM_R_X5Y134_SLICE_X6Y134_DQ;
  assign CLBLM_R_X7Y136_SLICE_X9Y136_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A1 = CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A2 = CLBLM_R_X7Y135_SLICE_X9Y135_A5Q;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A3 = CLBLM_R_X7Y136_SLICE_X8Y136_AQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A4 = CLBLM_R_X7Y133_SLICE_X8Y133_DQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_A6 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D1 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D2 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D3 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D4 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D5 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X7Y126_D6 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B2 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B3 = CLBLM_R_X3Y138_SLICE_X2Y138_AQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B4 = CLBLM_L_X12Y136_SLICE_X16Y136_A5Q;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_B5 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A1 = CLBLM_R_X5Y126_SLICE_X6Y126_BO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A2 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A3 = CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A4 = CLBLM_R_X5Y137_SLICE_X6Y137_BQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A5 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C1 = CLBLM_R_X5Y140_SLICE_X7Y140_A5Q;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C2 = CLBLM_R_X7Y131_SLICE_X8Y131_A5Q;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_AX = CLBLM_R_X5Y127_SLICE_X6Y127_DO6;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B1 = CLBLM_R_X5Y128_SLICE_X6Y128_DO6;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B2 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B3 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B4 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B5 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_B6 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D1 = CLBLM_R_X3Y135_SLICE_X3Y135_CQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D2 = CLBLM_L_X10Y141_SLICE_X12Y141_BQ;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C1 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C2 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C3 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C4 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C5 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_C6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B3 = 1'b1;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D5 = CLBLM_R_X3Y135_SLICE_X2Y135_DQ;
  assign CLBLM_R_X7Y136_SLICE_X8Y136_D6 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D1 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D2 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D3 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D4 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D5 = 1'b1;
  assign CLBLM_R_X5Y126_SLICE_X6Y126_D6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_B6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C2 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_C5 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A1 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A3 = CLBLM_L_X8Y143_SLICE_X11Y143_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A4 = CLBLM_L_X8Y143_SLICE_X11Y143_BO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A5 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_A6 = CLBLM_L_X8Y143_SLICE_X11Y143_CO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B1 = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B2 = CLBLM_L_X8Y143_SLICE_X10Y143_BO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B3 = CLBLM_L_X8Y143_SLICE_X11Y143_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B4 = CLBLM_L_X8Y141_SLICE_X11Y141_BQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B5 = CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_B6 = CLBLM_R_X7Y133_SLICE_X8Y133_A5Q;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C2 = CLBLL_L_X4Y137_SLICE_X5Y137_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C1 = CLBLM_R_X7Y143_SLICE_X8Y143_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C2 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C3 = CLBLM_L_X8Y143_SLICE_X10Y143_BO5;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C4 = CLBLM_L_X8Y141_SLICE_X10Y141_CO6;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C5 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_C6 = CLBLM_R_X7Y143_SLICE_X8Y143_A5Q;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_D1 = CLBLM_L_X10Y137_SLICE_X13Y137_AQ;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D1 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D2 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D3 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D4 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D5 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X11Y143_D6 = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_T1 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_D1 = CLBLM_L_X12Y143_SLICE_X16Y143_AO5;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C3 = CLBLM_L_X12Y136_SLICE_X16Y136_A5Q;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D1 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A1 = CLBLM_R_X7Y131_SLICE_X8Y131_AQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A2 = CLBLM_L_X8Y142_SLICE_X10Y142_CO5;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A3 = CLBLM_L_X8Y143_SLICE_X10Y143_AQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A5 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_A6 = CLBLM_R_X5Y140_SLICE_X7Y140_A5Q;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D2 = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_D1 = CLBLM_L_X10Y140_SLICE_X12Y140_AQ;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_T1 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D3 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B1 = CLBLM_R_X7Y143_SLICE_X8Y143_A5Q;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B2 = CLBLM_L_X8Y141_SLICE_X10Y141_BQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B3 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B4 = CLBLM_L_X8Y144_SLICE_X10Y144_AO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B5 = CLBLM_R_X7Y143_SLICE_X9Y143_AQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_B6 = 1'b1;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D4 = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_T1 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_D1 = CLBLM_R_X11Y140_SLICE_X14Y140_AO5;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D5 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C1 = CLBLM_R_X7Y133_SLICE_X8Y133_A5Q;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C2 = CLBLM_L_X8Y141_SLICE_X10Y141_AQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C3 = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C4 = CLBLM_L_X8Y144_SLICE_X10Y144_AO6;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C5 = CLBLM_L_X8Y141_SLICE_X10Y141_BQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_C6 = CLBLM_L_X8Y141_SLICE_X11Y141_BQ;
  assign CLBLM_R_X7Y129_SLICE_X8Y129_D6 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C4 = CLBLM_L_X8Y135_SLICE_X10Y135_B5Q;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_T1 = 1'b1;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D1 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D2 = CLBLM_R_X5Y137_SLICE_X7Y137_B5Q;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D3 = CLBLM_L_X8Y140_SLICE_X11Y140_B5Q;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D4 = CLBLM_L_X8Y142_SLICE_X10Y142_BO5;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D5 = CLBLM_L_X8Y142_SLICE_X11Y142_AQ;
  assign CLBLM_L_X8Y143_SLICE_X10Y143_D6 = CLBLM_R_X7Y143_SLICE_X9Y143_BO5;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1 = CLBLM_R_X3Y140_SLICE_X3Y140_AQ;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_C4 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_C5 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C6 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X17Y140_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1 = CLBLL_L_X4Y142_SLICE_X5Y142_AQ;
  assign LIOB33_X0Y143_IOB_X0Y143_O = CLBLL_L_X4Y138_SLICE_X4Y138_AO5;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A1 = CLBLM_R_X7Y137_SLICE_X9Y137_CQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A2 = CLBLM_R_X5Y133_SLICE_X7Y133_AQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A3 = CLBLM_R_X7Y137_SLICE_X9Y137_AQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A4 = CLBLL_L_X4Y135_SLICE_X4Y135_D5Q;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A5 = CLBLM_R_X5Y135_SLICE_X6Y135_AQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_A6 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B1 = CLBLM_R_X7Y137_SLICE_X9Y137_CQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B2 = CLBLM_R_X7Y137_SLICE_X9Y137_BQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B4 = CLBLM_R_X7Y137_SLICE_X9Y137_D5Q;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B5 = CLBLM_L_X12Y132_SLICE_X16Y132_AO6;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_B6 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A1 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A2 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A3 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A4 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A5 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_A6 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C1 = CLBLL_L_X4Y136_SLICE_X4Y136_D5Q;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C2 = CLBLM_R_X7Y137_SLICE_X9Y137_CQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_C3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B1 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B2 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B3 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B4 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B5 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_B6 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D2 = CLBLM_R_X7Y131_SLICE_X9Y131_CQ;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C1 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C2 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C3 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C4 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C5 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_C6 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D3 = CLBLM_L_X8Y139_SLICE_X11Y139_AQ;
  assign CLBLM_R_X7Y137_SLICE_X9Y137_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_A6 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A1 = CLBLM_R_X7Y133_SLICE_X8Y133_DQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A2 = CLBLM_R_X7Y131_SLICE_X9Y131_D5Q;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A3 = CLBLM_R_X7Y137_SLICE_X8Y137_AQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A5 = CLBLM_R_X7Y138_SLICE_X8Y138_B5Q;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D1 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D2 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D3 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D4 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D5 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X7Y127_D6 = 1'b1;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_A6 = CLBLM_L_X10Y140_SLICE_X13Y140_D5Q;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B1 = CLBLM_R_X7Y140_SLICE_X8Y140_B5Q;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B2 = CLBLM_L_X8Y137_SLICE_X10Y137_CQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B3 = CLBLL_L_X4Y131_SLICE_X5Y131_B5Q;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_B4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A1 = CLBLM_R_X5Y135_SLICE_X7Y135_DQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A3 = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A4 = CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A5 = CLBLM_R_X5Y126_SLICE_X6Y126_BO6;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B1 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_A6 = CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_C1 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B2 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B1 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B2 = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B4 = CLBLM_R_X5Y127_SLICE_X6Y127_DO5;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B3 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B5 = CLBLM_R_X5Y126_SLICE_X6Y126_BO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_B6 = CLBLM_L_X8Y131_SLICE_X10Y131_CQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B4 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C1 = CLBLM_R_X5Y126_SLICE_X6Y126_BO6;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C2 = CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C3 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B5 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C5 = CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_C6 = CLBLM_L_X8Y132_SLICE_X10Y132_AQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D3 = CLBLM_R_X7Y138_SLICE_X8Y138_BQ;
  assign CLBLM_R_X7Y137_SLICE_X8Y137_D4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_B6 = 1'b1;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_X105Y177_IOB_X1Y177_O = CLBLM_L_X8Y140_SLICE_X11Y140_BQ;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_A4 = CLBLM_R_X11Y140_SLICE_X14Y140_DQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D1 = CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D2 = CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D3 = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D4 = CLBLL_L_X4Y130_SLICE_X4Y130_BQ;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y127_SLICE_X6Y127_D6 = 1'b1;
  assign RIOB33_X105Y179_IOB_X1Y180_O = CLBLM_R_X3Y135_SLICE_X2Y135_AQ;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOB33_X105Y179_IOB_X1Y179_O = CLBLM_R_X5Y139_SLICE_X6Y139_BQ;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_D = RIOB33_X105Y135_IOB_X1Y136_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_D = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C1 = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C2 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C3 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C4 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C5 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_C6 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_B3 = CLBLM_R_X11Y140_SLICE_X14Y140_BQ;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_B4 = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_B5 = CLBLM_L_X12Y135_SLICE_X17Y135_CO6;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A1 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A2 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A3 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A4 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A5 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_A6 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B1 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B2 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B3 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B4 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B5 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_B6 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C1 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C2 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C3 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C4 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C5 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_C6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D1 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D1 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D2 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D3 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D4 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D5 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X11Y144_D6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D2 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D3 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D4 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_C4 = CLBLM_R_X11Y140_SLICE_X14Y140_DQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A1 = CLBLM_R_X5Y137_SLICE_X7Y137_B5Q;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A2 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A3 = CLBLM_L_X8Y142_SLICE_X11Y142_AQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A4 = CLBLM_L_X8Y140_SLICE_X11Y140_B5Q;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_C5 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A5 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_A6 = CLBLM_L_X10Y141_SLICE_X12Y141_C5Q;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D5 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X13Y142_D6 = 1'b1;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_C6 = CLBLM_R_X11Y140_SLICE_X14Y140_CQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B1 = CLBLM_R_X5Y137_SLICE_X7Y137_B5Q;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B2 = CLBLM_L_X10Y141_SLICE_X13Y141_AQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B3 = CLBLM_L_X8Y142_SLICE_X11Y142_AQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B4 = CLBLM_L_X8Y140_SLICE_X11Y140_B5Q;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B5 = CLBLM_L_X10Y142_SLICE_X12Y142_AQ;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_B6 = CLBLM_L_X8Y141_SLICE_X10Y141_CO6;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C1 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C2 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C3 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C4 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C5 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_C6 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D1 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D2 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D3 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D4 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D5 = 1'b1;
  assign CLBLM_L_X8Y144_SLICE_X10Y144_D6 = 1'b1;
  assign LIOB33_X0Y145_IOB_X0Y146_O = CLBLM_R_X3Y141_SLICE_X3Y141_BO6;
  assign LIOB33_X0Y145_IOB_X0Y145_O = CLBLM_R_X3Y137_SLICE_X2Y137_DO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_A4 = CLBLM_L_X8Y143_SLICE_X10Y143_DO6;
  assign CLBLM_L_X12Y140_SLICE_X16Y140_D5 = CLBLM_L_X8Y138_SLICE_X10Y138_B5Q;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A1 = CLBLM_R_X3Y140_SLICE_X3Y140_C5Q;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A2 = CLBLM_R_X3Y133_SLICE_X3Y133_B5Q;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A3 = CLBLM_L_X10Y139_SLICE_X13Y139_CQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A4 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A5 = CLBLM_R_X7Y138_SLICE_X9Y138_B5Q;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_A6 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B1 = CLBLM_R_X7Y138_SLICE_X9Y138_B5Q;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B2 = CLBLM_L_X10Y141_SLICE_X12Y141_AQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B3 = CLBLM_R_X5Y138_SLICE_X7Y138_CO6;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B4 = CLBLM_R_X5Y130_SLICE_X7Y130_DQ;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_B6 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B4 = CLBLM_R_X7Y133_SLICE_X8Y133_A5Q;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A1 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A2 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A3 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A4 = 1'b1;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B5 = CLBLM_L_X8Y142_SLICE_X11Y142_CO5;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A5 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_A6 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_C1 = CLBLM_R_X5Y134_SLICE_X6Y134_CQ;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_B6 = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B1 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B2 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B3 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B4 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B5 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_B6 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C1 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C2 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C3 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C4 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C5 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_C6 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X9Y138_D3 = CLBLL_L_X4Y138_SLICE_X4Y138_BO5;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B3 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A1 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A2 = CLBLM_R_X5Y138_SLICE_X7Y138_BO6;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A4 = CLBLM_R_X7Y139_SLICE_X8Y139_BO6;
  assign CLBLL_L_X4Y129_SLICE_X5Y129_B4 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A5 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D1 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D2 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D3 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D4 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D5 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X7Y128_D6 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_A6 = CLBLM_L_X8Y131_SLICE_X11Y131_CQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B1 = CLBLM_R_X5Y140_SLICE_X6Y140_CQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B2 = CLBLM_R_X7Y135_SLICE_X8Y135_BQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_B4 = CLBLM_R_X5Y139_SLICE_X7Y139_B5Q;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A1 = CLBLM_R_X5Y142_SLICE_X6Y142_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A2 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A3 = CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A4 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A5 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_A6 = CLBLM_R_X5Y128_SLICE_X6Y128_CO6;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C4 = CLBLM_R_X7Y133_SLICE_X8Y133_A5Q;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C1 = CLBLM_R_X7Y131_SLICE_X9Y131_AQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_C2 = CLBLM_R_X7Y138_SLICE_X8Y138_CQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C5 = CLBLM_R_X5Y138_SLICE_X6Y138_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B2 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B3 = CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B4 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B5 = CLBLM_R_X5Y128_SLICE_X6Y128_CO5;
  assign CLBLM_L_X10Y142_SLICE_X12Y142_C6 = CLBLM_L_X8Y142_SLICE_X11Y142_BQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_B6 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C1 = CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C2 = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C3 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C4 = CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C5 = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_C6 = 1'b1;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D2 = CLBLM_R_X7Y130_SLICE_X9Y130_BQ;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D3 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D4 = CLBLM_R_X5Y139_SLICE_X6Y139_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y138_SLICE_X8Y138_D6 = 1'b1;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D1 = CLBLM_R_X5Y126_SLICE_X6Y126_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D2 = CLBLM_R_X5Y128_SLICE_X6Y128_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D3 = CLBLM_R_X5Y128_SLICE_X6Y128_BQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D4 = CLBLM_R_X5Y127_SLICE_X6Y127_CQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D5 = CLBLM_R_X5Y127_SLICE_X6Y127_AQ;
  assign CLBLM_R_X5Y128_SLICE_X6Y128_D6 = CLBLM_R_X5Y127_SLICE_X6Y127_BQ;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1 = CLBLM_R_X3Y134_SLICE_X2Y134_AO5;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1 = 1'b1;
endmodule
