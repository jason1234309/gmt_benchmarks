module top(
  input LIOB33_SING_X0Y50_IOB_X0Y50_IPAD,
  input LIOB33_X0Y51_IOB_X0Y51_IPAD,
  input LIOB33_X0Y51_IOB_X0Y52_IPAD,
  input LIOB33_X0Y53_IOB_X0Y53_IPAD,
  input LIOB33_X0Y53_IOB_X0Y54_IPAD,
  input LIOB33_X0Y55_IOB_X0Y55_IPAD,
  input LIOB33_X0Y55_IOB_X0Y56_IPAD,
  input LIOB33_X0Y57_IOB_X0Y57_IPAD,
  input LIOB33_X0Y57_IOB_X0Y58_IPAD,
  input LIOB33_X0Y59_IOB_X0Y59_IPAD,
  input LIOB33_X0Y59_IOB_X0Y60_IPAD,
  input LIOB33_X0Y61_IOB_X0Y61_IPAD,
  input LIOB33_X0Y61_IOB_X0Y62_IPAD,
  input LIOB33_X0Y63_IOB_X0Y63_IPAD,
  input LIOB33_X0Y63_IOB_X0Y64_IPAD,
  input LIOB33_X0Y65_IOB_X0Y65_IPAD,
  input LIOB33_X0Y65_IOB_X0Y66_IPAD,
  input LIOB33_X0Y67_IOB_X0Y67_IPAD,
  input LIOB33_X0Y67_IOB_X0Y68_IPAD,
  input LIOB33_X0Y69_IOB_X0Y69_IPAD,
  input LIOB33_X0Y69_IOB_X0Y70_IPAD,
  input LIOB33_X0Y71_IOB_X0Y71_IPAD,
  input LIOB33_X0Y71_IOB_X0Y72_IPAD,
  input LIOB33_X0Y73_IOB_X0Y73_IPAD,
  input LIOB33_X0Y73_IOB_X0Y74_IPAD,
  input LIOB33_X0Y75_IOB_X0Y75_IPAD,
  input LIOB33_X0Y75_IOB_X0Y76_IPAD,
  input LIOB33_X0Y77_IOB_X0Y77_IPAD,
  input LIOB33_X0Y77_IOB_X0Y78_IPAD,
  input LIOB33_X0Y79_IOB_X0Y79_IPAD,
  input RIOB33_SING_X105Y100_IOB_X1Y100_IPAD,
  input RIOB33_SING_X105Y149_IOB_X1Y149_IPAD,
  input RIOB33_X105Y101_IOB_X1Y101_IPAD,
  input RIOB33_X105Y101_IOB_X1Y102_IPAD,
  input RIOB33_X105Y103_IOB_X1Y103_IPAD,
  input RIOB33_X105Y103_IOB_X1Y104_IPAD,
  input RIOB33_X105Y105_IOB_X1Y105_IPAD,
  input RIOB33_X105Y105_IOB_X1Y106_IPAD,
  input RIOB33_X105Y107_IOB_X1Y107_IPAD,
  input RIOB33_X105Y107_IOB_X1Y108_IPAD,
  input RIOB33_X105Y109_IOB_X1Y109_IPAD,
  input RIOB33_X105Y109_IOB_X1Y110_IPAD,
  input RIOB33_X105Y111_IOB_X1Y111_IPAD,
  input RIOB33_X105Y111_IOB_X1Y112_IPAD,
  input RIOB33_X105Y113_IOB_X1Y113_IPAD,
  input RIOB33_X105Y113_IOB_X1Y114_IPAD,
  input RIOB33_X105Y115_IOB_X1Y115_IPAD,
  input RIOB33_X105Y115_IOB_X1Y116_IPAD,
  input RIOB33_X105Y117_IOB_X1Y117_IPAD,
  input RIOB33_X105Y117_IOB_X1Y118_IPAD,
  input RIOB33_X105Y119_IOB_X1Y119_IPAD,
  input RIOB33_X105Y119_IOB_X1Y120_IPAD,
  input RIOB33_X105Y121_IOB_X1Y121_IPAD,
  input RIOB33_X105Y121_IOB_X1Y122_IPAD,
  input RIOB33_X105Y123_IOB_X1Y123_IPAD,
  input RIOB33_X105Y123_IOB_X1Y124_IPAD,
  input RIOB33_X105Y125_IOB_X1Y125_IPAD,
  input RIOB33_X105Y125_IOB_X1Y126_IPAD,
  input RIOB33_X105Y127_IOB_X1Y127_IPAD,
  input RIOB33_X105Y127_IOB_X1Y128_IPAD,
  input RIOB33_X105Y129_IOB_X1Y129_IPAD,
  input RIOB33_X105Y129_IOB_X1Y130_IPAD,
  input RIOB33_X105Y131_IOB_X1Y131_IPAD,
  input RIOB33_X105Y131_IOB_X1Y132_IPAD,
  input RIOB33_X105Y133_IOB_X1Y133_IPAD,
  input RIOB33_X105Y133_IOB_X1Y134_IPAD,
  input RIOB33_X105Y135_IOB_X1Y135_IPAD,
  input RIOB33_X105Y135_IOB_X1Y136_IPAD,
  input RIOB33_X105Y137_IOB_X1Y137_IPAD,
  input RIOB33_X105Y137_IOB_X1Y138_IPAD,
  input RIOB33_X105Y139_IOB_X1Y139_IPAD,
  input RIOB33_X105Y139_IOB_X1Y140_IPAD,
  input RIOB33_X105Y141_IOB_X1Y141_IPAD,
  input RIOB33_X105Y141_IOB_X1Y142_IPAD,
  input RIOB33_X105Y143_IOB_X1Y143_IPAD,
  input RIOB33_X105Y143_IOB_X1Y144_IPAD,
  input RIOB33_X105Y145_IOB_X1Y145_IPAD,
  input RIOB33_X105Y145_IOB_X1Y146_IPAD,
  input RIOB33_X105Y147_IOB_X1Y147_IPAD,
  input RIOB33_X105Y147_IOB_X1Y148_IPAD,
  output LIOB33_SING_X0Y100_IOB_X0Y100_OPAD,
  output LIOB33_SING_X0Y149_IOB_X0Y149_OPAD,
  output LIOB33_SING_X0Y150_IOB_X0Y150_OPAD,
  output LIOB33_SING_X0Y199_IOB_X0Y199_OPAD,
  output LIOB33_X0Y101_IOB_X0Y101_OPAD,
  output LIOB33_X0Y101_IOB_X0Y102_OPAD,
  output LIOB33_X0Y103_IOB_X0Y103_OPAD,
  output LIOB33_X0Y103_IOB_X0Y104_OPAD,
  output LIOB33_X0Y105_IOB_X0Y105_OPAD,
  output LIOB33_X0Y105_IOB_X0Y106_OPAD,
  output LIOB33_X0Y107_IOB_X0Y107_OPAD,
  output LIOB33_X0Y107_IOB_X0Y108_OPAD,
  output LIOB33_X0Y109_IOB_X0Y109_OPAD,
  output LIOB33_X0Y109_IOB_X0Y110_OPAD,
  output LIOB33_X0Y111_IOB_X0Y111_OPAD,
  output LIOB33_X0Y111_IOB_X0Y112_OPAD,
  output LIOB33_X0Y113_IOB_X0Y113_OPAD,
  output LIOB33_X0Y113_IOB_X0Y114_OPAD,
  output LIOB33_X0Y115_IOB_X0Y115_OPAD,
  output LIOB33_X0Y115_IOB_X0Y116_OPAD,
  output LIOB33_X0Y117_IOB_X0Y117_OPAD,
  output LIOB33_X0Y117_IOB_X0Y118_OPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD,
  output LIOB33_X0Y125_IOB_X0Y125_OPAD,
  output LIOB33_X0Y125_IOB_X0Y126_OPAD,
  output LIOB33_X0Y127_IOB_X0Y127_OPAD,
  output LIOB33_X0Y127_IOB_X0Y128_OPAD,
  output LIOB33_X0Y129_IOB_X0Y129_OPAD,
  output LIOB33_X0Y129_IOB_X0Y130_OPAD,
  output LIOB33_X0Y131_IOB_X0Y131_OPAD,
  output LIOB33_X0Y131_IOB_X0Y132_OPAD,
  output LIOB33_X0Y133_IOB_X0Y133_OPAD,
  output LIOB33_X0Y133_IOB_X0Y134_OPAD,
  output LIOB33_X0Y135_IOB_X0Y135_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output LIOB33_X0Y141_IOB_X0Y141_OPAD,
  output LIOB33_X0Y141_IOB_X0Y142_OPAD,
  output LIOB33_X0Y143_IOB_X0Y143_OPAD,
  output LIOB33_X0Y145_IOB_X0Y145_OPAD,
  output LIOB33_X0Y145_IOB_X0Y146_OPAD,
  output LIOB33_X0Y147_IOB_X0Y147_OPAD,
  output LIOB33_X0Y147_IOB_X0Y148_OPAD,
  output LIOB33_X0Y151_IOB_X0Y151_OPAD,
  output LIOB33_X0Y151_IOB_X0Y152_OPAD,
  output LIOB33_X0Y153_IOB_X0Y153_OPAD,
  output LIOB33_X0Y153_IOB_X0Y154_OPAD,
  output LIOB33_X0Y155_IOB_X0Y155_OPAD,
  output LIOB33_X0Y155_IOB_X0Y156_OPAD,
  output LIOB33_X0Y157_IOB_X0Y157_OPAD,
  output LIOB33_X0Y157_IOB_X0Y158_OPAD,
  output LIOB33_X0Y159_IOB_X0Y159_OPAD,
  output LIOB33_X0Y159_IOB_X0Y160_OPAD,
  output LIOB33_X0Y161_IOB_X0Y161_OPAD,
  output LIOB33_X0Y161_IOB_X0Y162_OPAD,
  output LIOB33_X0Y163_IOB_X0Y163_OPAD,
  output LIOB33_X0Y163_IOB_X0Y164_OPAD,
  output LIOB33_X0Y165_IOB_X0Y165_OPAD,
  output LIOB33_X0Y165_IOB_X0Y166_OPAD,
  output LIOB33_X0Y167_IOB_X0Y167_OPAD,
  output LIOB33_X0Y167_IOB_X0Y168_OPAD,
  output LIOB33_X0Y169_IOB_X0Y169_OPAD,
  output LIOB33_X0Y169_IOB_X0Y170_OPAD,
  output LIOB33_X0Y171_IOB_X0Y171_OPAD,
  output LIOB33_X0Y171_IOB_X0Y172_OPAD,
  output LIOB33_X0Y173_IOB_X0Y173_OPAD,
  output LIOB33_X0Y173_IOB_X0Y174_OPAD,
  output LIOB33_X0Y175_IOB_X0Y175_OPAD,
  output LIOB33_X0Y175_IOB_X0Y176_OPAD,
  output LIOB33_X0Y177_IOB_X0Y177_OPAD,
  output LIOB33_X0Y177_IOB_X0Y178_OPAD,
  output LIOB33_X0Y179_IOB_X0Y179_OPAD,
  output LIOB33_X0Y179_IOB_X0Y180_OPAD,
  output LIOB33_X0Y181_IOB_X0Y181_OPAD,
  output LIOB33_X0Y181_IOB_X0Y182_OPAD,
  output LIOB33_X0Y183_IOB_X0Y183_OPAD,
  output LIOB33_X0Y183_IOB_X0Y184_OPAD,
  output LIOB33_X0Y185_IOB_X0Y185_OPAD,
  output LIOB33_X0Y185_IOB_X0Y186_OPAD,
  output LIOB33_X0Y187_IOB_X0Y187_OPAD,
  output LIOB33_X0Y187_IOB_X0Y188_OPAD,
  output LIOB33_X0Y189_IOB_X0Y189_OPAD,
  output LIOB33_X0Y189_IOB_X0Y190_OPAD,
  output LIOB33_X0Y191_IOB_X0Y191_OPAD,
  output LIOB33_X0Y191_IOB_X0Y192_OPAD,
  output LIOB33_X0Y193_IOB_X0Y193_OPAD,
  output LIOB33_X0Y193_IOB_X0Y194_OPAD,
  output LIOB33_X0Y195_IOB_X0Y195_OPAD,
  output LIOB33_X0Y195_IOB_X0Y196_OPAD,
  output LIOB33_X0Y197_IOB_X0Y197_OPAD,
  output LIOB33_X0Y197_IOB_X0Y198_OPAD,
  output LIOB33_X0Y79_IOB_X0Y80_OPAD,
  output RIOB33_SING_X105Y150_IOB_X1Y150_OPAD,
  output RIOB33_SING_X105Y199_IOB_X1Y199_OPAD,
  output RIOB33_X105Y151_IOB_X1Y151_OPAD,
  output RIOB33_X105Y151_IOB_X1Y152_OPAD,
  output RIOB33_X105Y153_IOB_X1Y153_OPAD,
  output RIOB33_X105Y153_IOB_X1Y154_OPAD,
  output RIOB33_X105Y155_IOB_X1Y155_OPAD,
  output RIOB33_X105Y155_IOB_X1Y156_OPAD,
  output RIOB33_X105Y157_IOB_X1Y157_OPAD,
  output RIOB33_X105Y157_IOB_X1Y158_OPAD,
  output RIOB33_X105Y159_IOB_X1Y159_OPAD,
  output RIOB33_X105Y159_IOB_X1Y160_OPAD,
  output RIOB33_X105Y161_IOB_X1Y161_OPAD,
  output RIOB33_X105Y161_IOB_X1Y162_OPAD,
  output RIOB33_X105Y163_IOB_X1Y163_OPAD,
  output RIOB33_X105Y163_IOB_X1Y164_OPAD,
  output RIOB33_X105Y165_IOB_X1Y165_OPAD,
  output RIOB33_X105Y165_IOB_X1Y166_OPAD,
  output RIOB33_X105Y167_IOB_X1Y167_OPAD,
  output RIOB33_X105Y167_IOB_X1Y168_OPAD,
  output RIOB33_X105Y169_IOB_X1Y169_OPAD,
  output RIOB33_X105Y169_IOB_X1Y170_OPAD,
  output RIOB33_X105Y171_IOB_X1Y171_OPAD,
  output RIOB33_X105Y171_IOB_X1Y172_OPAD,
  output RIOB33_X105Y173_IOB_X1Y173_OPAD,
  output RIOB33_X105Y173_IOB_X1Y174_OPAD,
  output RIOB33_X105Y175_IOB_X1Y175_OPAD,
  output RIOB33_X105Y175_IOB_X1Y176_OPAD,
  output RIOB33_X105Y177_IOB_X1Y177_OPAD,
  output RIOB33_X105Y177_IOB_X1Y178_OPAD,
  output RIOB33_X105Y179_IOB_X1Y179_OPAD,
  output RIOB33_X105Y179_IOB_X1Y180_OPAD,
  output RIOB33_X105Y181_IOB_X1Y181_OPAD,
  output RIOB33_X105Y181_IOB_X1Y182_OPAD,
  output RIOB33_X105Y183_IOB_X1Y183_OPAD,
  output RIOB33_X105Y183_IOB_X1Y184_OPAD,
  output RIOB33_X105Y185_IOB_X1Y185_OPAD,
  output RIOB33_X105Y185_IOB_X1Y186_OPAD,
  output RIOB33_X105Y187_IOB_X1Y187_OPAD,
  output RIOB33_X105Y187_IOB_X1Y188_OPAD,
  output RIOB33_X105Y189_IOB_X1Y189_OPAD,
  output RIOB33_X105Y189_IOB_X1Y190_OPAD,
  output RIOB33_X105Y191_IOB_X1Y191_OPAD,
  output RIOB33_X105Y191_IOB_X1Y192_OPAD,
  output RIOB33_X105Y193_IOB_X1Y193_OPAD,
  output RIOB33_X105Y193_IOB_X1Y194_OPAD,
  output RIOB33_X105Y195_IOB_X1Y195_OPAD,
  output RIOB33_X105Y195_IOB_X1Y196_OPAD,
  output RIOB33_X105Y197_IOB_X1Y197_OPAD,
  output RIOB33_X105Y197_IOB_X1Y198_OPAD
  );
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_A;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_A1;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_A2;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_A3;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_A4;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_A5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_A6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_AMUX;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_AO5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_AO6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_A_CY;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_A_XOR;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_B;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_B1;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_B2;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_B3;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_B4;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_B5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_B6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_BMUX;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_BO5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_BO6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_B_CY;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_B_XOR;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_C;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_C1;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_C2;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_C3;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_C4;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_C5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_C6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_CO5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_CO6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_C_CY;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_C_XOR;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_D;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_D1;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_D2;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_D3;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_D4;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_D5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_D6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_DO5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_DO6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_D_CY;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X0Y139_D_XOR;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_A;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_A1;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_A2;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_A3;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_A4;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_A5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_A6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_AO5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_AO6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_A_CY;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_A_XOR;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_B;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_B1;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_B2;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_B3;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_B4;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_B5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_B6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_BO5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_BO6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_B_CY;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_B_XOR;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_C;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_C1;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_C2;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_C3;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_C4;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_C5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_C6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_CO5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_CO6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_C_CY;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_C_XOR;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_D;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_D1;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_D2;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_D3;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_D4;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_D5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_D6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_DO5;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_DO6;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_D_CY;
  wire [0:0] CLBLL_L_X2Y139_SLICE_X1Y139_D_XOR;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_A;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_A1;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_A2;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_A3;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_A4;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_A5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_A6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_AMUX;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_AO5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_AO6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_A_CY;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_A_XOR;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_B;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_B1;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_B2;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_B3;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_B4;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_B5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_B6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_BMUX;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_BO5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_BO6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_B_CY;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_B_XOR;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_C;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_C1;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_C2;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_C3;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_C4;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_C5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_C6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_CO5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_CO6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_C_CY;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_C_XOR;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_D;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_D1;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_D2;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_D3;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_D4;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_D5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_D6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_DO5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_DO6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_D_CY;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X0Y140_D_XOR;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_A;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_A1;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_A2;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_A3;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_A4;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_A5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_A6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_AO5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_AO6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_A_CY;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_A_XOR;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_B;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_B1;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_B2;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_B3;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_B4;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_B5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_B6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_BO5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_BO6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_B_CY;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_B_XOR;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_C;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_C1;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_C2;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_C3;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_C4;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_C5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_C6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_CO5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_CO6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_C_CY;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_C_XOR;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_D;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_D1;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_D2;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_D3;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_D4;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_D5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_D6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_DO5;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_DO6;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_D_CY;
  wire [0:0] CLBLL_L_X2Y140_SLICE_X1Y140_D_XOR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A1;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A2;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A3;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A4;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_AO5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_AO6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A_CY;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_A_XOR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B1;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B2;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B3;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B4;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_BO5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_BO6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B_CY;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_B_XOR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C1;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C2;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C3;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C4;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_CO5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_CO6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C_CY;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_C_XOR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D1;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D2;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D3;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D4;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_DO5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_DO6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D_CY;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X0Y153_D_XOR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A1;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A2;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A3;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A4;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_AMUX;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_AO5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_AO6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A_CY;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_A_XOR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B1;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B2;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B3;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B4;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_BO5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B_CY;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_B_XOR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C1;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C2;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C3;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C4;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_CO5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_CO6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C_CY;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_C_XOR;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D1;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D2;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D3;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D4;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_DO5;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_DO6;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D_CY;
  wire [0:0] CLBLL_L_X2Y153_SLICE_X1Y153_D_XOR;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_A;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_A1;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_A2;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_A3;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_A4;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_A5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_A6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_AO5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_AO6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_A_CY;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_A_XOR;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_B;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_B1;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_B2;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_B3;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_B4;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_B5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_B6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_BO5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_BO6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_B_CY;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_B_XOR;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_C;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_C1;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_C2;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_C3;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_C4;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_C5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_C6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_CO5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_CO6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_C_CY;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_C_XOR;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_D;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_D1;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_D2;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_D3;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_D4;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_D5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_D6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_DO5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_DO6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_D_CY;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X0Y154_D_XOR;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_A;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_A1;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_A2;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_A3;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_A4;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_A5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_A6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_AMUX;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_AO5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_AO6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_A_CY;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_A_XOR;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_B;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_B1;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_B2;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_B3;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_B4;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_B5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_B6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_BO5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_BO6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_B_CY;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_B_XOR;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_C;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_C1;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_C2;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_C3;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_C4;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_C5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_C6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_CO5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_CO6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_C_CY;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_C_XOR;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_D;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_D1;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_D2;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_D3;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_D4;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_D5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_D6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_DO5;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_DO6;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_D_CY;
  wire [0:0] CLBLL_L_X2Y154_SLICE_X1Y154_D_XOR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A1;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A2;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A3;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A4;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_AO5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_AO6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A_CY;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_A_XOR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B1;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B2;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B3;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B4;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_BO5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_BO6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B_CY;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_B_XOR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C1;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C2;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C3;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C4;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_CO5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_CO6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C_CY;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_C_XOR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D1;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D2;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D3;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D4;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_DO5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_DO6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D_CY;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X0Y155_D_XOR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A1;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A2;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A3;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A4;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_AMUX;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_AO5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_AO6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A_CY;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_A_XOR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B1;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B2;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B3;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B4;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_BMUX;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_BO5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_BO6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B_CY;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_B_XOR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C1;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C2;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C3;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C4;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_CMUX;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_CO5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_CO6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C_CY;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_C_XOR;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D1;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D2;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D3;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D4;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_DO5;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D_CY;
  wire [0:0] CLBLL_L_X2Y155_SLICE_X1Y155_D_XOR;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_A;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_A1;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_A2;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_A3;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_A4;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_A5;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_A6;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_AO5;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_AO6;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_A_CY;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_A_XOR;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_B;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_B1;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_B2;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_B3;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_B4;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_B5;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_B6;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_BO5;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_BO6;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_B_CY;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_B_XOR;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_C;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_C1;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_C2;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_C3;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_C4;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_C5;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_C6;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_CO5;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_CO6;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_C_CY;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_C_XOR;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_D;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_D1;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_D2;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_D3;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_D4;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_D5;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_D6;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_DO5;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_DO6;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_D_CY;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X54Y150_D_XOR;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_A;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_A1;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_A2;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_A3;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_A4;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_A5;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_A6;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_AO5;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_AO6;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_A_CY;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_A_XOR;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_B;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_B1;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_B2;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_B3;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_B4;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_B5;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_B6;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_BO5;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_BO6;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_B_CY;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_B_XOR;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_C;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_C1;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_C2;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_C3;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_C4;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_C5;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_C6;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_CO5;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_CO6;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_C_CY;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_C_XOR;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_D;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_D1;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_D2;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_D3;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_D4;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_D5;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_D6;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_DO5;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_DO6;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_D_CY;
  wire [0:0] CLBLL_L_X36Y150_SLICE_X55Y150_D_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_AO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_AO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_A_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_BO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_BO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_B_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_CO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_CO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_C_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_DO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_DO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X4Y146_D_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_AMUX;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_AO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_AQ;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_A_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_BO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_BO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_B_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_CLK;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_CO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_CO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_C_XOR;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D1;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D2;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D3;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D4;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_DO5;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_DO6;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D_CY;
  wire [0:0] CLBLL_L_X4Y146_SLICE_X5Y146_D_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_AO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_AO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_A_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_BO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_BO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_B_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_CO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_CO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_C_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_DO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_DO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X4Y147_D_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_AO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_AO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_AQ;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_A_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_BO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_BO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_B_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_CLK;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_CO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_CO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_C_XOR;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D1;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D2;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D3;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D4;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_DO5;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_DO6;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D_CY;
  wire [0:0] CLBLL_L_X4Y147_SLICE_X5Y147_D_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_AO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_AO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_AQ;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_A_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_BMUX;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_BO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_BO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_B_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_CLK;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_CO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_CO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_C_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_DO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_DO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X4Y148_D_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_AO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_AO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_AQ;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_A_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_BO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_BO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_B_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_CLK;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_CO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_CO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_CQ;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_C_XOR;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D1;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D2;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D3;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D4;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_DO5;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_DO6;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_DQ;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D_CY;
  wire [0:0] CLBLL_L_X4Y148_SLICE_X5Y148_D_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A5Q;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_AMUX;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_AO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_AO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_AQ;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_AX;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_A_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_BO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_BO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_BQ;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_B_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_CLK;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_CO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_CO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_C_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_DO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_DO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X4Y149_D_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A5Q;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_AMUX;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_AO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_AO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_AQ;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_AX;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_A_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_BMUX;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_BO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_BO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_B_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_CLK;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_CMUX;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_CO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_CO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_C_XOR;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D1;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D2;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D3;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D4;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_DMUX;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_DO5;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_DO6;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D_CY;
  wire [0:0] CLBLL_L_X4Y149_SLICE_X5Y149_D_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_AO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_AO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_AQ;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_A_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_BO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_BO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_BQ;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_B_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_CLK;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_CO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_CO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_CQ;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_C_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_DO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X4Y150_D_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_AO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_AO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_AQ;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_A_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_BO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_BO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_BQ;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_B_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C5Q;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_CLK;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_CMUX;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_CO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_CO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_CQ;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_C_XOR;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D1;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D2;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D3;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D4;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D5Q;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_DMUX;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_DO5;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_DO6;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_DQ;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D_CY;
  wire [0:0] CLBLL_L_X4Y150_SLICE_X5Y150_D_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_AO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_AO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_A_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_BO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_BO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_BQ;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_B_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C5Q;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_CLK;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_CMUX;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_CO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_CO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_CQ;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_C_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D5Q;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_DMUX;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_DO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_DO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_DQ;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X4Y151_D_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_AO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_AO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_AQ;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_A_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_BO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_BO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_BQ;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_B_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_CLK;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_CO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_CO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_CQ;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_C_XOR;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D1;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D2;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D3;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D4;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_DO5;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_DO6;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D_CY;
  wire [0:0] CLBLL_L_X4Y151_SLICE_X5Y151_D_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_AO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_AO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_AQ;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_A_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_BO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_BO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_B_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_CLK;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_CO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_CO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_C_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_DO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_DO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X4Y152_D_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_AO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_AO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_AQ;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_A_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_BO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_BO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_BQ;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_B_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_CLK;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_CO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_CO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_CQ;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_C_XOR;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D1;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D2;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D3;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D4;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_DMUX;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_DO5;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_DO6;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D_CY;
  wire [0:0] CLBLL_L_X4Y152_SLICE_X5Y152_D_XOR;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A1;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A2;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A3;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A4;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_AO5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_AO6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A_CY;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_A_XOR;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B1;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B2;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B3;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B4;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_BO5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_BO6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B_CY;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_B_XOR;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C1;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C2;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C3;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C4;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_CO5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_CO6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C_CY;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_C_XOR;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D1;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D2;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D3;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D4;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_DO5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_DO6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D_CY;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X4Y153_D_XOR;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A1;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A2;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A3;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A4;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_AO5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_AO6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_AQ;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A_CY;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_A_XOR;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B1;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B2;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B3;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B4;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_BO5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_BO6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B_CY;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_B_XOR;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C1;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C2;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C3;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C4;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_CLK;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_CO5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_CO6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C_CY;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_C_XOR;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D1;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D2;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D3;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D4;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_DMUX;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_DO5;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_DO6;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D_CY;
  wire [0:0] CLBLL_L_X4Y153_SLICE_X5Y153_D_XOR;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_A;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_A1;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_A2;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_A3;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_A4;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_A5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_A6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_AO5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_AO6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_A_CY;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_A_XOR;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_B;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_B1;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_B2;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_B3;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_B4;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_B5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_B6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_BO5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_BO6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_B_CY;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_B_XOR;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_C;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_C1;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_C2;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_C3;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_C4;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_C5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_C6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_CO5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_CO6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_C_CY;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_C_XOR;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_D;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_D1;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_D2;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_D3;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_D4;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_D5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_D6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_DMUX;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_DO5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_DO6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_D_CY;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X4Y154_D_XOR;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_A;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_A1;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_A2;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_A3;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_A4;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_A5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_A6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_AO5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_AO6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_AQ;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_A_CY;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_A_XOR;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_B;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_B1;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_B2;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_B3;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_B4;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_B5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_B6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_BO5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_BO6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_B_CY;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_B_XOR;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_C;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_C1;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_C2;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_C3;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_C4;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_C5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_C6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_CLK;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_CO5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_CO6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_C_CY;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_C_XOR;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_D;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_D1;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_D2;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_D3;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_D4;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_D5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_D6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_DO5;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_DO6;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_D_CY;
  wire [0:0] CLBLL_L_X4Y154_SLICE_X5Y154_D_XOR;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A1;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A2;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A3;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A4;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_AO5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_AO6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_AQ;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A_CY;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_A_XOR;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B1;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B2;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B3;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B4;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_BO5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_BO6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_BQ;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B_CY;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_B_XOR;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C1;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C2;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C3;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C4;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_CLK;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_CO5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_CO6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C_CY;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_C_XOR;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D1;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D2;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D3;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D4;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_DO5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_DO6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D_CY;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X4Y155_D_XOR;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A1;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A2;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A3;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A4;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A5Q;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_AMUX;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_AO5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_AO6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_AQ;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A_CY;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_A_XOR;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B1;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B2;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B3;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B4;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_BO5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_BO6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_BQ;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B_CY;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_B_XOR;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C1;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C2;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C3;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C4;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_CLK;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_CO5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_CO6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C_CY;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_C_XOR;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D1;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D2;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D3;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D4;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_DO5;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_DO6;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D_CY;
  wire [0:0] CLBLL_L_X4Y155_SLICE_X5Y155_D_XOR;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_A;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_A1;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_A2;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_A3;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_A4;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_A5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_A6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_AMUX;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_AO5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_AO6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_AQ;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_A_CY;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_A_XOR;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_B;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_B1;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_B2;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_B3;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_B4;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_B5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_B6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_BMUX;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_BO5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_BO6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_B_CY;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_B_XOR;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_C;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_C1;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_C2;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_C3;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_C4;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_C5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_C6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_CLK;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_CMUX;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_CO5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_CO6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_C_CY;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_C_XOR;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_D;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_D1;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_D2;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_D3;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_D4;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_D5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_D6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_DO5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_DO6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_D_CY;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X4Y156_D_XOR;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_A;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_A1;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_A2;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_A3;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_A4;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_A5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_A6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_AO5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_AO6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_A_CY;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_A_XOR;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_B;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_B1;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_B2;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_B3;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_B4;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_B5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_B6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_BO5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_BO6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_B_CY;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_B_XOR;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_C;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_C1;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_C2;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_C3;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_C4;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_C5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_C6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_CMUX;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_CO5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_CO6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_C_CY;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_C_XOR;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_D;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_D1;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_D2;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_D3;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_D4;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_D5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_D6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_DMUX;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_DO5;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_DO6;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_D_CY;
  wire [0:0] CLBLL_L_X4Y156_SLICE_X5Y156_D_XOR;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_A;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_A1;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_A2;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_A3;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_A4;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_A5;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_A6;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_AMUX;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_AO5;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_AO6;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_A_CY;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_A_XOR;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_B;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_B1;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_B2;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_B3;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_B4;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_B5;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_B6;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_BMUX;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_BO5;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_BO6;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_B_CY;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_B_XOR;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_C;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_C1;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_C2;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_C3;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_C4;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_C5;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_C6;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_CMUX;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_CO5;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_CO6;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_C_CY;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_C_XOR;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_D;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_D1;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_D2;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_D3;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_D4;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_D5;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_D6;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_DO5;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_DO6;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_D_CY;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X4Y157_D_XOR;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_A;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_A1;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_A2;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_A3;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_A4;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_A5;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_A6;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_AMUX;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_AO5;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_AO6;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_A_CY;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_A_XOR;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_B;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_B1;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_B2;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_B3;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_B4;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_B5;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_B6;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_BO5;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_BO6;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_B_CY;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_B_XOR;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_C;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_C1;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_C2;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_C3;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_C4;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_C5;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_C6;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_CO5;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_CO6;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_C_CY;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_C_XOR;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_D;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_D1;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_D2;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_D3;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_D4;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_D5;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_D6;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_DO5;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_DO6;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_D_CY;
  wire [0:0] CLBLL_L_X4Y157_SLICE_X5Y157_D_XOR;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_A;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_A1;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_A2;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_A3;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_A4;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_A5;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_A6;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_AO5;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_AO6;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_A_CY;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_A_XOR;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_B;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_B1;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_B2;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_B3;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_B4;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_B5;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_B6;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_BO5;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_BO6;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_B_CY;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_B_XOR;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_C;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_C1;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_C2;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_C3;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_C4;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_C5;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_C6;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_CO5;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_CO6;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_C_CY;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_C_XOR;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_D;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_D1;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_D2;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_D3;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_D4;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_D5;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_D6;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_DO5;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_DO6;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_D_CY;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X4Y158_D_XOR;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_A;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_A1;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_A2;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_A3;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_A4;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_A5;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_A6;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_AO5;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_AO6;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_AQ;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_AX;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_A_CY;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_A_XOR;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_B;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_B1;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_B2;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_B3;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_B4;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_B5;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_B6;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_BO5;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_BO6;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_B_CY;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_B_XOR;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_C;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_C1;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_C2;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_C3;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_C4;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_C5;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_C6;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_CLK;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_CO5;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_CO6;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_C_CY;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_C_XOR;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_D;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_D1;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_D2;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_D3;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_D4;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_D5;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_D6;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_DO5;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_DO6;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_D_CY;
  wire [0:0] CLBLL_L_X4Y158_SLICE_X5Y158_D_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_AO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_A_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_BO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_BO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_B_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_CO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_CO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_C_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_DO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_DO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X78Y126_D_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_AO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_AO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_A_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_BO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_BO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_B_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_CO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_CO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_C_XOR;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D1;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D2;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D3;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D4;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_DO5;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_DO6;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D_CY;
  wire [0:0] CLBLL_L_X52Y126_SLICE_X79Y126_D_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_AMUX;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_AO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_A_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_BO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_BO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_B_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_CLK;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_CO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_CO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_C_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_DO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_DO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X12Y144_D_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_AO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_AO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_A_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_BO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_BO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_B_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_CO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_C_XOR;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D1;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D2;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D3;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D4;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_DO5;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_DO6;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D_CY;
  wire [0:0] CLBLM_L_X10Y144_SLICE_X13Y144_D_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_AO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_AO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_A_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_BO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_BO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_BQ;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_B_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_CLK;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_CO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_CO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_CQ;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_C_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_DO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_DO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X12Y145_D_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_AO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_AQ;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_A_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_BO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_BQ;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_B_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_CLK;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_CO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_CQ;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_C_XOR;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D1;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D2;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D3;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D4;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_DMUX;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_DO5;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_DO6;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D_CY;
  wire [0:0] CLBLM_L_X10Y145_SLICE_X13Y145_D_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_AO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_AO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_AQ;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_A_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_BO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_BO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_BQ;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_B_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C5Q;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_CLK;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_CMUX;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_CO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_CO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_CQ;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_C_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_DO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_DO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X12Y146_D_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_AO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_AO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_A_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_BMUX;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_BO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_BO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_B_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_CO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_CO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_C_XOR;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D1;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D2;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D3;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D4;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_DO5;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D_CY;
  wire [0:0] CLBLM_L_X10Y146_SLICE_X13Y146_D_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_AO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_AO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_AQ;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_A_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_BO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_BO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_BQ;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_B_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_CLK;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_CO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_CO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_CQ;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_C_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_DO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_DO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_DQ;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X12Y147_D_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_AO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_AO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_AQ;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_A_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_BO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_BO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_BQ;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_B_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_CLK;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_CO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_CO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_CQ;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_C_XOR;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D1;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D2;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D3;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D4;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_DMUX;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_DO5;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_DO6;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D_CY;
  wire [0:0] CLBLM_L_X10Y147_SLICE_X13Y147_D_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_AO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_AO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_AQ;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_A_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_BMUX;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_BO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_BO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_B_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_CLK;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_CMUX;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_CO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_CO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_C_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_DO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_DO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X12Y148_D_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_AO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_AO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_AQ;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_A_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_BO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_BO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_BQ;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_B_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_CLK;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_CO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_CO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_CQ;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_C_XOR;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D1;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D2;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D3;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D4;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_DO5;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_DO6;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D_CY;
  wire [0:0] CLBLM_L_X10Y148_SLICE_X13Y148_D_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_AO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_AO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_AQ;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_A_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_BO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_BO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_BQ;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_B_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C5Q;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_CLK;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_CMUX;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_CO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_CO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_CQ;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_C_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_DMUX;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_DO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_DO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X12Y149_D_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A5Q;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_AMUX;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_AO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_AO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_AX;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_A_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_BMUX;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_BO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_BO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_BQ;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_BX;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_B_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_CLK;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_CMUX;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_CO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_CO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_C_XOR;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D1;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D2;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D3;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D4;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_DO5;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_DO6;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D_CY;
  wire [0:0] CLBLM_L_X10Y149_SLICE_X13Y149_D_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A5Q;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_AMUX;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_AO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_AO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_AQ;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_A_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_BMUX;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_BO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_BO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_BQ;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_BX;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_B_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_CLK;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_CO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_CO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_CQ;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_CX;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_C_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_DO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_DO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X12Y150_D_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_AO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_AO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_AQ;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_A_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B5Q;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_BMUX;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_BO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_BO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_BQ;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_B_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C5Q;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_CLK;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_CMUX;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_CO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_CO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_CQ;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_C_XOR;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D1;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D2;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D3;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D4;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_DO5;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_DO6;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D_CY;
  wire [0:0] CLBLM_L_X10Y150_SLICE_X13Y150_D_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_AO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_AO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_AQ;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_A_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_BO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_BO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_BQ;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_B_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_CLK;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_CO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_CO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_CQ;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_C_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_DO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_DO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_DQ;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X12Y151_D_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_AO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_AO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_AQ;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_A_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B5Q;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_BMUX;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_BO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_BO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_BQ;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_B_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_CLK;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_CO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_CO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_CQ;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_C_XOR;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D1;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D2;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D3;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D4;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_DO5;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_DO6;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D_CY;
  wire [0:0] CLBLM_L_X10Y151_SLICE_X13Y151_D_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_AO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_AO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_AQ;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_A_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_BO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_BO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_BQ;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_B_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_CLK;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_CMUX;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_CO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_CO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_C_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_DO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_DO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X12Y152_D_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_AO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_AO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_AQ;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_A_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_BMUX;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_BO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_BO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_B_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_CLK;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_CMUX;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_CO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_CO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_C_XOR;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D1;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D2;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D3;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D4;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_DO5;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_DO6;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D_CY;
  wire [0:0] CLBLM_L_X10Y152_SLICE_X13Y152_D_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_AO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_AO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_AQ;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_A_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_BO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_BO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_BQ;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_B_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_CLK;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_CO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_CO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_C_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_DO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_DO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X12Y153_D_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_AO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_AO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_AQ;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_A_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_BMUX;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_BO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_BO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_B_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_CLK;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_CO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_CO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_CQ;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_C_XOR;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D1;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D2;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D3;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D4;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_DO5;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_DO6;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_DQ;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D_CY;
  wire [0:0] CLBLM_L_X10Y153_SLICE_X13Y153_D_XOR;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_A;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_A1;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_A2;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_A3;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_A4;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_A5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_A5Q;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_A6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_AMUX;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_AO5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_AO6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_AQ;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_AX;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_A_CY;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_A_XOR;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_B;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_B1;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_B2;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_B3;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_B4;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_B5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_B6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_BMUX;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_BO5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_BO6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_B_CY;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_B_XOR;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_C;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_C1;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_C2;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_C3;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_C4;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_C5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_C6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_CLK;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_CO5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_CO6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_CQ;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_C_CY;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_C_XOR;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_D;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_D1;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_D2;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_D3;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_D4;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_D5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_D6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_DO5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_DO6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_DQ;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_D_CY;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X12Y154_D_XOR;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_A;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_A1;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_A2;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_A3;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_A4;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_A5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_A6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_AMUX;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_AO5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_AO6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_AQ;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_A_CY;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_A_XOR;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_B;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_B1;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_B2;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_B3;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_B4;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_B5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_B6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_BO5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_BO6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_BQ;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_B_CY;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_B_XOR;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_C;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_C1;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_C2;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_C3;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_C4;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_C5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_C5Q;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_C6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_CLK;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_CMUX;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_CO5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_CO6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_CQ;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_C_CY;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_C_XOR;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_D;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_D1;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_D2;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_D3;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_D4;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_D5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_D6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_DO5;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_DO6;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_DQ;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_D_CY;
  wire [0:0] CLBLM_L_X10Y154_SLICE_X13Y154_D_XOR;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_A;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_A1;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_A2;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_A3;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_A4;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_A5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_A6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_AO5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_AO6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_AQ;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_A_CY;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_A_XOR;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_B;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_B1;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_B2;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_B3;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_B4;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_B5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_B6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_BO5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_BO6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_BQ;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_B_CY;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_B_XOR;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_C;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_C1;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_C2;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_C3;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_C4;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_C5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_C6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_CLK;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_CO5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_CO6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_CQ;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_C_CY;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_C_XOR;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_D;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_D1;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_D2;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_D3;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_D4;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_D5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_D6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_DO5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_DO6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_D_CY;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X12Y155_D_XOR;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_A;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_A1;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_A2;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_A3;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_A4;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_A5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_A5Q;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_A6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_AMUX;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_AO5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_AO6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_AQ;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_A_CY;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_A_XOR;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_B;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_B1;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_B2;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_B3;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_B4;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_B5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_B6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_BO5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_BO6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_BQ;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_B_CY;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_B_XOR;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_C;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_C1;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_C2;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_C3;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_C4;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_C5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_C6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_CLK;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_CO5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_CO6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_C_CY;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_C_XOR;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_D;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_D1;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_D2;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_D3;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_D4;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_D5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_D6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_DMUX;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_DO5;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_DO6;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_D_CY;
  wire [0:0] CLBLM_L_X10Y155_SLICE_X13Y155_D_XOR;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_A;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_A1;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_A2;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_A3;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_A4;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_A5;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_A6;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_AO5;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_AO6;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_AQ;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_A_CY;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_A_XOR;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_B;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_B1;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_B2;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_B3;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_B4;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_B5;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_B6;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_BO5;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_BO6;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_B_CY;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_B_XOR;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_C;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_C1;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_C2;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_C3;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_C4;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_C5;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_C6;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_CLK;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_CMUX;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_CO5;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_CO6;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_C_CY;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_C_XOR;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_D;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_D1;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_D2;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_D3;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_D4;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_D5;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_D6;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_DO5;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_DO6;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_D_CY;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X12Y156_D_XOR;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_A;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_A1;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_A2;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_A3;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_A4;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_A5;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_A6;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_AMUX;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_AO5;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_AO6;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_A_CY;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_A_XOR;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_B;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_B1;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_B2;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_B3;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_B4;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_B5;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_B6;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_BO5;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_BO6;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_BQ;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_B_CY;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_B_XOR;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_C;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_C1;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_C2;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_C3;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_C4;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_C5;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_C6;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_CLK;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_CO5;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_CO6;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_C_CY;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_C_XOR;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_D;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_D1;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_D2;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_D3;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_D4;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_D5;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_D6;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_DO5;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_DO6;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_D_CY;
  wire [0:0] CLBLM_L_X10Y156_SLICE_X13Y156_D_XOR;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_A;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_A1;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_A2;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_A3;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_A4;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_A5;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_A6;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_AO5;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_AO6;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_AQ;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_A_CY;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_A_XOR;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_B;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_B1;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_B2;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_B3;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_B4;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_B5;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_B6;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_BO5;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_BO6;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_BQ;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_B_CY;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_B_XOR;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_C;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_C1;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_C2;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_C3;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_C4;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_C5;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_C6;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_CLK;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_CMUX;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_CO5;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_CO6;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_C_CY;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_C_XOR;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_D;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_D1;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_D2;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_D3;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_D4;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_D5;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_D6;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_DO5;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_DO6;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_D_CY;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X12Y157_D_XOR;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_A;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_A1;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_A2;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_A3;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_A4;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_A5;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_A6;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_AMUX;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_AO5;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_AO6;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_A_CY;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_A_XOR;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_B;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_B1;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_B2;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_B3;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_B4;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_B5;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_B6;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_BO5;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_BO6;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_B_CY;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_B_XOR;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_C;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_C1;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_C2;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_C3;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_C4;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_C5;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_C6;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_CO5;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_CO6;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_C_CY;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_C_XOR;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_D;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_D1;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_D2;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_D3;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_D4;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_D5;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_D6;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_DO5;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_DO6;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_D_CY;
  wire [0:0] CLBLM_L_X10Y157_SLICE_X13Y157_D_XOR;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_A;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_A1;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_A2;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_A3;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_A4;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_A5;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_A6;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_AO5;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_AO6;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_AQ;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_A_CY;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_A_XOR;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_B;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_B1;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_B2;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_B3;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_B4;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_B5;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_B6;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_BO5;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_BO6;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_BQ;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_B_CY;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_B_XOR;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_C;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_C1;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_C2;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_C3;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_C4;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_C5;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_C6;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_CLK;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_CO5;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_CO6;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_C_CY;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_C_XOR;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_D;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_D1;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_D2;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_D3;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_D4;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_D5;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_D6;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_DO5;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_DO6;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_D_CY;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X12Y158_D_XOR;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_A;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_A1;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_A2;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_A3;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_A4;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_A5;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_A6;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_AO5;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_AO6;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_AQ;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_A_CY;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_A_XOR;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_B;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_B1;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_B2;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_B3;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_B4;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_B5;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_B6;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_BO5;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_BO6;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_BQ;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_B_CY;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_B_XOR;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_C;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_C1;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_C2;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_C3;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_C4;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_C5;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_C6;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_CLK;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_CO5;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_CO6;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_C_CY;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_C_XOR;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_D;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_D1;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_D2;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_D3;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_D4;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_D5;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_D6;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_DO5;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_DO6;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_D_CY;
  wire [0:0] CLBLM_L_X10Y158_SLICE_X13Y158_D_XOR;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_A;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_A1;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_A2;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_A3;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_A4;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_A5;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_A6;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_AO5;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_AO6;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_A_CY;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_A_XOR;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_B;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_B1;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_B2;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_B3;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_B4;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_B5;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_B6;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_BO5;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_BO6;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_B_CY;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_B_XOR;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_C;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_C1;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_C2;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_C3;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_C4;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_C5;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_C6;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_CO5;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_CO6;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_C_CY;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_C_XOR;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_D;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_D1;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_D2;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_D3;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_D4;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_D5;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_D6;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_DO5;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_DO6;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_D_CY;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X12Y159_D_XOR;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_A;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_A1;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_A2;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_A3;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_A4;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_A5;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_A6;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_AMUX;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_AO5;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_AO6;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_A_CY;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_A_XOR;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_B;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_B1;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_B2;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_B3;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_B4;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_B5;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_B6;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_BMUX;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_BO5;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_BO6;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_B_CY;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_B_XOR;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_C;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_C1;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_C2;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_C3;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_C4;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_C5;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_C6;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_CO5;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_CO6;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_C_CY;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_C_XOR;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_D;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_D1;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_D2;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_D3;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_D4;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_D5;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_D6;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_DO5;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_DO6;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_D_CY;
  wire [0:0] CLBLM_L_X10Y159_SLICE_X13Y159_D_XOR;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_A;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_A1;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_A2;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_A3;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_A4;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_A5;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_A6;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_AO5;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_AO6;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_A_CY;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_A_XOR;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_B;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_B1;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_B2;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_B3;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_B4;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_B5;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_B6;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_BO5;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_BO6;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_B_CY;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_B_XOR;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_C;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_C1;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_C2;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_C3;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_C4;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_C5;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_C6;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_CO5;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_CO6;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_C_CY;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_C_XOR;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_D;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_D1;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_D2;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_D3;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_D4;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_D5;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_D6;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_DO5;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_DO6;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_D_CY;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X12Y163_D_XOR;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_A;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_A1;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_A2;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_A3;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_A4;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_A5;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_A6;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_AO5;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_AO6;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_A_CY;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_A_XOR;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_B;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_B1;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_B2;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_B3;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_B4;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_B5;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_B6;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_BO5;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_BO6;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_B_CY;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_B_XOR;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_C;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_C1;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_C2;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_C3;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_C4;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_C5;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_C6;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_CO5;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_CO6;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_C_CY;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_C_XOR;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_D;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_D1;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_D2;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_D3;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_D4;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_D5;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_D6;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_DO5;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_DO6;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_D_CY;
  wire [0:0] CLBLM_L_X10Y163_SLICE_X13Y163_D_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_AO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_AO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_AQ;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_A_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_BO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_BO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_BQ;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_B_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_CLK;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_CO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_CQ;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_C_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_DO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_DO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_DQ;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X16Y146_D_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_AO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_AO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_A_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_BO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_BO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_B_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_CO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_CO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_C_XOR;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D1;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D2;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D3;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D4;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_DO5;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_DO6;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D_CY;
  wire [0:0] CLBLM_L_X12Y146_SLICE_X17Y146_D_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_AO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_AO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_AQ;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_A_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_BMUX;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_BO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_BO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_B_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_CLK;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_CO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_CO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_C_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_DO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X16Y147_D_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_AO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_AO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_A_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_BO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_BO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_B_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_CO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_CO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_C_XOR;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D1;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D2;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D3;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D4;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_DO5;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_DO6;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D_CY;
  wire [0:0] CLBLM_L_X12Y147_SLICE_X17Y147_D_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_AMUX;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_AO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_AO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_A_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_BO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_BO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_B_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_CO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_CO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_C_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_DO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_DO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X16Y148_D_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_AO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_AO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_A_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_BO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_BO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_B_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_CO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_CO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_C_XOR;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D1;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D2;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D3;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D4;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_DMUX;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_DO5;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_DO6;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D_CY;
  wire [0:0] CLBLM_L_X12Y148_SLICE_X17Y148_D_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_AO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_AO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_AQ;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_A_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B5Q;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_BMUX;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_BO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_BO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_BQ;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_B_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_CLK;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_CO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_CO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_CQ;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_C_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_DO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_DO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_DQ;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X16Y149_D_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A5Q;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_AMUX;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_AO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_AO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_AQ;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_AX;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_A_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_BMUX;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_BO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_BO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_B_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_CLK;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_CMUX;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_CO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_CO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_C_XOR;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D1;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D2;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D3;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D4;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_DMUX;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_DO5;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_DO6;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D_CY;
  wire [0:0] CLBLM_L_X12Y149_SLICE_X17Y149_D_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A5Q;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_AMUX;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_AO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_AO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_AQ;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_AX;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_A_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_BO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_BO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_BQ;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_B_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_CLK;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_CO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_CO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_CQ;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_C_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_DO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_DO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X16Y150_D_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_AO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_AO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_AQ;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_A_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_BO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_BO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_BQ;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_B_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_CLK;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_CO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_CO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_C_XOR;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D1;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D2;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D3;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D4;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_DO5;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_DO6;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D_CY;
  wire [0:0] CLBLM_L_X12Y150_SLICE_X17Y150_D_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_AO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_AO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_A_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_BO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_BO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_BQ;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_B_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C5Q;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_CLK;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_CMUX;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_CO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_CO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_CQ;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_C_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_DO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X16Y151_D_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A5Q;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_AMUX;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_AO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_AO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_AQ;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_A_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_BO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_BO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_BQ;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_B_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_CLK;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_CO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_CO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_C_XOR;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D1;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D2;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D3;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D4;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_DO5;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_DO6;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D_CY;
  wire [0:0] CLBLM_L_X12Y151_SLICE_X17Y151_D_XOR;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A1;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A2;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A3;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A4;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_AMUX;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_AO5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_AO6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_AQ;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A_CY;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_A_XOR;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B1;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B2;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B3;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B4;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B5Q;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_BMUX;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_BO5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_BO6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_BQ;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_BX;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B_CY;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_B_XOR;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C1;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C2;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C3;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C4;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_CLK;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_CO5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_CO6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_CQ;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C_CY;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_C_XOR;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D1;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D2;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D3;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D4;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_DO5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_DO6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D_CY;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X16Y152_D_XOR;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A1;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A2;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A3;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A4;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A5Q;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_AMUX;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_AO5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_AO6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_AQ;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_AX;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A_CY;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_A_XOR;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B1;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B2;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B3;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B4;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_BMUX;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_BO5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_BO6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B_CY;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_B_XOR;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C1;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C2;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C3;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C4;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_CLK;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_CO5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_CO6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C_CY;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_C_XOR;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D1;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D2;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D3;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D4;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_DO5;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_DO6;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D_CY;
  wire [0:0] CLBLM_L_X12Y152_SLICE_X17Y152_D_XOR;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A1;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A2;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A3;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A4;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_AO5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_AO6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_AQ;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A_CY;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_A_XOR;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B1;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B2;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B3;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B4;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_BMUX;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_BO5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_BO6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B_CY;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_B_XOR;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C1;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C2;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C3;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C4;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_CLK;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_CO5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_CO6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C_CY;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_C_XOR;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D1;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D2;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D3;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D4;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_DO5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_DO6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D_CY;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X16Y153_D_XOR;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A1;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A2;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A3;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A4;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_AO5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_AO6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_AQ;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A_CY;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_A_XOR;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B1;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B2;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B3;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B4;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_BO5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_BO6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_BQ;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B_CY;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_B_XOR;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C1;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C2;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C3;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C4;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_CLK;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_CO5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_CO6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_CQ;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C_CY;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_C_XOR;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D1;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D2;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D3;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D4;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_DMUX;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_DO5;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_DO6;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D_CY;
  wire [0:0] CLBLM_L_X12Y153_SLICE_X17Y153_D_XOR;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_A;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_A1;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_A2;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_A3;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_A4;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_A5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_A5Q;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_A6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_AMUX;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_AO5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_AO6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_AQ;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_AX;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_A_CY;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_A_XOR;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_B;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_B1;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_B2;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_B3;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_B4;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_B5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_B6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_BO5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_BO6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_BQ;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_B_CY;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_B_XOR;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_C;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_C1;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_C2;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_C3;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_C4;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_C5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_C6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_CLK;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_CMUX;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_CO5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_CO6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_C_CY;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_C_XOR;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_D;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_D1;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_D2;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_D3;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_D4;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_D5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_D6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_DMUX;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_DO5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_DO6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_D_CY;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X16Y154_D_XOR;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_A;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_A1;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_A2;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_A3;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_A4;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_A5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_A5Q;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_A6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_AMUX;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_AO5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_AO6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_AQ;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_AX;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_A_CY;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_A_XOR;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_B;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_B1;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_B2;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_B3;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_B4;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_B5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_B6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_BO5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_BO6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_BQ;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_B_CY;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_B_XOR;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_C;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_C1;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_C2;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_C3;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_C4;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_C5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_C6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_CLK;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_CMUX;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_CO5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_CO6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_C_CY;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_C_XOR;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_D;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_D1;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_D2;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_D3;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_D4;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_D5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_D6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_DO5;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_DO6;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_DQ;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_D_CY;
  wire [0:0] CLBLM_L_X12Y154_SLICE_X17Y154_D_XOR;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_A;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_A1;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_A2;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_A3;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_A4;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_A5;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_A6;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_AMUX;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_AO5;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_AO6;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_AQ;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_AX;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_A_CY;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_A_XOR;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_B;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_B1;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_B2;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_B3;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_B4;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_B5;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_B6;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_BMUX;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_BO5;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_BO6;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_B_CY;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_B_XOR;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_C;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_C1;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_C2;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_C3;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_C4;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_C5;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_C6;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_CE;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_CLK;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_CO5;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_CO6;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_C_CY;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_C_XOR;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_D;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_D1;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_D2;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_D3;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_D4;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_D5;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_D6;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_DO5;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_DO6;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_D_CY;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_D_XOR;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X16Y155_SR;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_A;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_A1;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_A2;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_A3;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_A4;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_A5;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_A6;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_AO5;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_AO6;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_AQ;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_A_CY;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_A_XOR;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_B;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_B1;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_B2;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_B3;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_B4;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_B5;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_B6;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_BO5;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_BO6;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_BQ;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_B_CY;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_B_XOR;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_C;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_C1;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_C2;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_C3;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_C4;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_C5;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_C6;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_CLK;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_CO5;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_CO6;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_CQ;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_C_CY;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_C_XOR;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_D;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_D1;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_D2;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_D3;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_D4;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_D5;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_D6;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_DMUX;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_DO5;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_DO6;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_D_CY;
  wire [0:0] CLBLM_L_X12Y155_SLICE_X17Y155_D_XOR;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_A;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_A1;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_A2;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_A3;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_A4;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_A5;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_A6;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_AO5;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_AO6;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_AQ;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_AX;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_A_CY;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_A_XOR;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_B;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_B1;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_B2;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_B3;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_B4;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_B5;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_B6;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_BO5;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_BO6;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_BQ;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_BX;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_B_CY;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_B_XOR;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_C;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_C1;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_C2;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_C3;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_C4;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_C5;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_C6;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_CE;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_CLK;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_CO5;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_CO6;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_C_CY;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_C_XOR;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_D;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_D1;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_D2;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_D3;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_D4;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_D5;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_D6;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_DO5;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_DO6;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_D_CY;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_D_XOR;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X16Y156_SR;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_A;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_A1;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_A2;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_A3;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_A4;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_A5;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_A6;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_AO5;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_AO6;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_AQ;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_A_CY;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_A_XOR;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_B;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_B1;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_B2;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_B3;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_B4;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_B5;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_B6;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_BO5;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_BO6;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_BQ;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_B_CY;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_B_XOR;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_C;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_C1;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_C2;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_C3;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_C4;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_C5;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_C6;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_CLK;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_CO5;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_CO6;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_C_CY;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_C_XOR;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_D;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_D1;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_D2;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_D3;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_D4;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_D5;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_D6;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_DO5;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_DO6;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_D_CY;
  wire [0:0] CLBLM_L_X12Y156_SLICE_X17Y156_D_XOR;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_A;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_A1;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_A2;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_A3;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_A4;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_A5;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_A5Q;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_A6;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_AMUX;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_AO5;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_AO6;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_AQ;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_AX;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_A_CY;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_A_XOR;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_B;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_B1;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_B2;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_B3;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_B4;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_B5;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_B6;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_BO5;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_BO6;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_BQ;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_B_CY;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_B_XOR;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_C;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_C1;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_C2;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_C3;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_C4;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_C5;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_C6;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_CLK;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_CO5;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_CO6;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_CQ;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_C_CY;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_C_XOR;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_D;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_D1;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_D2;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_D3;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_D4;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_D5;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_D6;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_DMUX;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_DO5;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_DO6;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_D_CY;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X16Y157_D_XOR;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_A;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_A1;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_A2;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_A3;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_A4;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_A5;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_A5Q;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_A6;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_AMUX;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_AO5;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_AO6;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_AQ;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_AX;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_A_CY;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_A_XOR;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_B;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_B1;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_B2;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_B3;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_B4;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_B5;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_B6;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_BO5;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_BO6;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_BQ;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_B_CY;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_B_XOR;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_C;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_C1;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_C2;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_C3;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_C4;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_C5;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_C6;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_CLK;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_CO5;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_CO6;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_CQ;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_C_CY;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_C_XOR;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_D;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_D1;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_D2;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_D3;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_D4;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_D5;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_D6;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_DO5;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_DO6;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_D_CY;
  wire [0:0] CLBLM_L_X12Y157_SLICE_X17Y157_D_XOR;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_A;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_A1;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_A2;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_A3;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_A4;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_A5;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_A5Q;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_A6;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_AMUX;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_AO5;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_AO6;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_AQ;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_AX;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_A_CY;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_A_XOR;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_B;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_B1;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_B2;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_B3;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_B4;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_B5;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_B6;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_BMUX;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_BO5;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_BO6;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_B_CY;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_B_XOR;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_C;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_C1;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_C2;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_C3;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_C4;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_C5;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_C6;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_CLK;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_CMUX;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_CO5;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_CO6;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_C_CY;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_C_XOR;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_D;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_D1;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_D2;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_D3;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_D4;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_D5;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_D6;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_DMUX;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_DO5;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_DO6;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_D_CY;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X16Y158_D_XOR;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_A;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_A1;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_A2;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_A3;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_A4;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_A5;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_A6;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_AO5;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_AO6;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_AQ;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_A_CY;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_A_XOR;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_B;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_B1;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_B2;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_B3;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_B4;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_B5;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_B6;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_BO5;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_BO6;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_BQ;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_B_CY;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_B_XOR;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_C;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_C1;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_C2;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_C3;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_C4;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_C5;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_C6;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_CLK;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_CO5;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_CO6;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_C_CY;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_C_XOR;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_D;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_D1;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_D2;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_D3;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_D4;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_D5;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_D6;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_DO5;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_DO6;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_D_CY;
  wire [0:0] CLBLM_L_X12Y158_SLICE_X17Y158_D_XOR;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_A;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_A1;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_A2;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_A3;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_A4;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_A5;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_A6;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_AMUX;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_AO5;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_AO6;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_AQ;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_AX;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_A_CY;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_A_XOR;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_B;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_B1;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_B2;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_B3;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_B4;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_B5;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_B6;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_BMUX;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_BO5;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_BO6;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_BQ;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_BX;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_B_CY;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_B_XOR;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_C;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_C1;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_C2;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_C3;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_C4;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_C5;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_C6;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_CE;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_CLK;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_CMUX;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_CO5;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_CO6;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_C_CY;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_C_XOR;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_D;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_D1;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_D2;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_D3;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_D4;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_D5;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_D6;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_DO5;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_DO6;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_D_CY;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_D_XOR;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X16Y159_SR;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_A;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_A1;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_A2;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_A3;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_A4;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_A5;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_A6;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_AMUX;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_AO5;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_AO6;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_A_CY;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_A_XOR;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_B;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_B1;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_B2;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_B3;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_B4;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_B5;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_B6;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_BO5;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_BO6;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_B_CY;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_B_XOR;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_C;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_C1;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_C2;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_C3;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_C4;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_C5;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_C6;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_CO5;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_CO6;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_C_CY;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_C_XOR;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_D;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_D1;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_D2;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_D3;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_D4;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_D5;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_D6;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_DO5;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_DO6;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_D_CY;
  wire [0:0] CLBLM_L_X12Y159_SLICE_X17Y159_D_XOR;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_A;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_A1;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_A2;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_A3;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_A4;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_A5;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_A6;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_AMUX;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_AO5;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_AO6;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_A_CY;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_A_XOR;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_B;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_B1;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_B2;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_B3;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_B4;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_B5;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_B6;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_BO5;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_BO6;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_B_CY;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_B_XOR;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_C;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_C1;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_C2;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_C3;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_C4;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_C5;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_C6;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_CO5;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_CO6;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_C_CY;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_C_XOR;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_D;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_D1;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_D2;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_D3;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_D4;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_D5;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_D6;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_DO5;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_DO6;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_D_CY;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X22Y156_D_XOR;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_A;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_A1;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_A2;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_A3;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_A4;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_A5;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_A6;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_AO5;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_AO6;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_A_CY;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_A_XOR;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_B;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_B1;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_B2;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_B3;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_B4;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_B5;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_B6;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_BO5;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_BO6;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_B_CY;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_B_XOR;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_C;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_C1;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_C2;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_C3;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_C4;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_C5;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_C6;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_CO5;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_CO6;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_C_CY;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_C_XOR;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_D;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_D1;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_D2;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_D3;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_D4;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_D5;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_D6;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_DO5;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_DO6;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_D_CY;
  wire [0:0] CLBLM_L_X16Y156_SLICE_X23Y156_D_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_AO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_A_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B5Q;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_BMUX;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_BO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_BO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_BQ;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_B_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_CLK;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_CO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_CO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_C_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_DO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_DO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X10Y146_D_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_AO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_AO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_AQ;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_A_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_BO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_BO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_BQ;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_B_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_CLK;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_CO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_CO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_CQ;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_C_XOR;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D1;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D2;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D3;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D4;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_DO5;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D_CY;
  wire [0:0] CLBLM_L_X8Y146_SLICE_X11Y146_D_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_AMUX;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_AO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_AO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_A_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_BO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_BO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_BQ;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_B_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_CLK;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_CO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_CO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_CQ;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_C_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_DMUX;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_DO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_DO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X10Y147_D_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_AO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_AO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_AQ;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_A_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_BO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_BQ;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_B_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_CLK;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_CO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_CO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_C_XOR;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D1;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D2;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D3;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D4;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_DO5;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_DO6;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D_CY;
  wire [0:0] CLBLM_L_X8Y147_SLICE_X11Y147_D_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_AO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_AO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_AQ;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_A_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_BO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_BO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_BQ;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_B_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_CLK;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_CO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_CO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_CQ;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_C_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_DO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_DO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X10Y148_D_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A5Q;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_AMUX;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_AO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_AO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_AQ;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_AX;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_A_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B5Q;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_BMUX;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_BO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_BO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_BQ;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_B_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_CLK;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_CMUX;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_CO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_CO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_C_XOR;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D1;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D2;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D3;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D4;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_DMUX;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_DO5;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_DO6;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D_CY;
  wire [0:0] CLBLM_L_X8Y148_SLICE_X11Y148_D_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_AO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_AO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_AQ;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_A_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_BMUX;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_BO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_BO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_B_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_CLK;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_CO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_CO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_C_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_DO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_DO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X10Y149_D_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_AO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_AO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_A_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_BO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_BO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_BQ;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_B_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_CLK;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_CO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_CO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_CQ;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_C_XOR;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D1;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D2;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D3;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D4;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_DO5;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_DO6;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D_CY;
  wire [0:0] CLBLM_L_X8Y149_SLICE_X11Y149_D_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_AMUX;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_AO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_AO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_AX;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_A_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_BO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_BO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_BQ;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_B_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_CLK;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_CMUX;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_CO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_CO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_C_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_DO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_DO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X10Y150_D_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_AO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_AO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_AQ;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_A_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_BO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_BO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_BQ;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_B_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_CLK;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_CO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_CO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_CQ;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_C_XOR;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D1;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D2;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D3;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D4;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_DO5;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_DO6;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D_CY;
  wire [0:0] CLBLM_L_X8Y150_SLICE_X11Y150_D_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_AO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_AO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_A_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_BO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_BO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_BQ;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_B_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_CLK;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_CO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_CO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_CQ;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_C_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_DO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_DO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X10Y151_D_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_AO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_AO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_AQ;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_A_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_BO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_BO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_B_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_CLK;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_CO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_CO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_C_XOR;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D1;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D2;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D3;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D4;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_DO5;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_DO6;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D_CY;
  wire [0:0] CLBLM_L_X8Y151_SLICE_X11Y151_D_XOR;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A1;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A2;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A3;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A4;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_AO5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_AO6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_AQ;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A_CY;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_A_XOR;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B1;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B2;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B3;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B4;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_BO5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_BO6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_BQ;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B_CY;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_B_XOR;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C1;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C2;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C3;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C4;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_CLK;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_CO5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_CO6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_CQ;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C_CY;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_C_XOR;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D1;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D2;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D3;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D4;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_DO5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_DO6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D_CY;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X10Y152_D_XOR;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A1;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A2;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A3;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A4;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_AMUX;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_AO5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_AO6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A_CY;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_A_XOR;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B1;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B2;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B3;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B4;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_BMUX;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_BO5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_BO6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B_CY;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_B_XOR;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C1;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C2;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C3;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C4;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_CO5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_CO6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C_CY;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_C_XOR;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D1;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D2;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D3;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D4;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_DO5;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_DO6;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D_CY;
  wire [0:0] CLBLM_L_X8Y152_SLICE_X11Y152_D_XOR;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A1;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A2;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A3;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A4;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A5Q;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_AMUX;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_AO5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_AO6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_AQ;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A_CY;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_A_XOR;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B1;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B2;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B3;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B4;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_BO5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_BO6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B_CY;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_B_XOR;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C1;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C2;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C3;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C4;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_CLK;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_CO5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_CO6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C_CY;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_C_XOR;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D1;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D2;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D3;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D4;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_DO5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_DO6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D_CY;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X10Y153_D_XOR;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A1;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A2;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A3;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A4;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_AO5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_AO6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_AQ;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A_CY;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_A_XOR;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B1;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B2;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B3;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B4;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_BO5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_BO6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_BQ;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B_CY;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_B_XOR;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C1;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C2;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C3;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C4;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C5Q;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_CLK;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_CMUX;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_CO5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_CO6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_CQ;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C_CY;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_C_XOR;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D1;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D2;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D3;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D4;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_DO5;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_DO6;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_DQ;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D_CY;
  wire [0:0] CLBLM_L_X8Y153_SLICE_X11Y153_D_XOR;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A1;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A2;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A3;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A4;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A5Q;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_AMUX;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_AO5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_AO6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_AQ;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A_CY;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_A_XOR;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B1;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B2;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B3;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B4;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B5Q;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_BMUX;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_BO5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_BO6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_BQ;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B_CY;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_B_XOR;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C1;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C2;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C3;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C4;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C5Q;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_CLK;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_CMUX;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_CO5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_CO6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_CQ;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C_CY;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_C_XOR;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D1;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D2;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D3;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D4;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_DO5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_DO6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_DQ;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D_CY;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X10Y154_D_XOR;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A1;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A2;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A3;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A4;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A5Q;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_AMUX;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_AO5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_AO6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_AQ;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_AX;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A_CY;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_A_XOR;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B1;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B2;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B3;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B4;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_BO5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_BO6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_BQ;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B_CY;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_B_XOR;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C1;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C2;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C3;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C4;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_CLK;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_CO5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_CO6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_CQ;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C_CY;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_C_XOR;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D1;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D2;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D3;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D4;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_DO5;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_DO6;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D_CY;
  wire [0:0] CLBLM_L_X8Y154_SLICE_X11Y154_D_XOR;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_A;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_A1;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_A2;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_A3;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_A4;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_A5;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_A6;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_AO5;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_AO6;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_AQ;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_A_CY;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_A_XOR;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_B;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_B1;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_B2;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_B3;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_B4;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_B5;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_B5Q;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_B6;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_BMUX;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_BO5;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_BO6;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_BQ;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_B_CY;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_B_XOR;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_C;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_C1;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_C2;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_C3;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_C4;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_C5;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_C6;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_CLK;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_CO5;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_CO6;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_CQ;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_C_CY;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_C_XOR;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_D;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_D1;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_D2;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_D3;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_D4;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_D5;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_D6;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_DO5;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_DO6;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_D_CY;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X10Y155_D_XOR;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_A;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_A1;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_A2;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_A3;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_A4;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_A5;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_A6;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_AO5;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_AO6;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_AQ;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_A_CY;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_A_XOR;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_B;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_B1;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_B2;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_B3;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_B4;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_B5;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_B6;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_BO5;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_BO6;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_BQ;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_B_CY;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_B_XOR;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_C;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_C1;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_C2;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_C3;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_C4;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_C5;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_C6;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_CLK;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_CO5;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_CO6;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_CQ;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_C_CY;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_C_XOR;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_D;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_D1;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_D2;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_D3;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_D4;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_D5;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_D6;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_DO5;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_DO6;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_D_CY;
  wire [0:0] CLBLM_L_X8Y155_SLICE_X11Y155_D_XOR;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_A;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_A1;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_A2;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_A3;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_A4;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_A5;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_A6;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_AO5;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_AO6;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_AQ;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_A_CY;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_A_XOR;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_B;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_B1;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_B2;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_B3;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_B4;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_B5;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_B6;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_BO5;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_BO6;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_BQ;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_B_CY;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_B_XOR;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_C;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_C1;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_C2;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_C3;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_C4;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_C5;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_C6;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_CLK;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_CO5;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_CO6;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_CQ;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_C_CY;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_C_XOR;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_D;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_D1;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_D2;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_D3;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_D4;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_D5;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_D6;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_DO5;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_DO6;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_D_CY;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X10Y156_D_XOR;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_A;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_A1;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_A2;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_A3;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_A4;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_A5;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_A6;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_AO5;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_AO6;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_AQ;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_A_CY;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_A_XOR;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_B;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_B1;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_B2;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_B3;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_B4;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_B5;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_B5Q;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_B6;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_BMUX;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_BO5;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_BO6;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_BQ;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_B_CY;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_B_XOR;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_C;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_C1;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_C2;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_C3;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_C4;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_C5;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_C6;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_CLK;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_CO5;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_CO6;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_C_CY;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_C_XOR;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_D;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_D1;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_D2;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_D3;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_D4;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_D5;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_D6;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_DO5;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_DO6;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_D_CY;
  wire [0:0] CLBLM_L_X8Y156_SLICE_X11Y156_D_XOR;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_A;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_A1;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_A2;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_A3;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_A4;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_A5;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_A6;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_AO5;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_AO6;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_AQ;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_A_CY;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_A_XOR;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_B;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_B1;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_B2;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_B3;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_B4;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_B5;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_B6;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_BO5;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_BO6;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_BQ;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_B_CY;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_B_XOR;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_C;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_C1;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_C2;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_C3;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_C4;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_C5;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_C6;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_CLK;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_CO5;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_CO6;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_CQ;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_C_CY;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_C_XOR;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_D;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_D1;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_D2;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_D3;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_D4;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_D5;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_D6;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_DO5;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_DO6;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_DQ;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_D_CY;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X10Y157_D_XOR;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_A;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_A1;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_A2;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_A3;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_A4;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_A5;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_A6;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_AO5;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_AO6;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_AQ;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_A_CY;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_A_XOR;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_B;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_B1;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_B2;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_B3;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_B4;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_B5;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_B6;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_BO5;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_BO6;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_BQ;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_B_CY;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_B_XOR;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_C;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_C1;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_C2;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_C3;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_C4;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_C5;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_C6;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_CLK;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_CO5;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_CO6;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_CQ;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_C_CY;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_C_XOR;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_D;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_D1;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_D2;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_D3;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_D4;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_D5;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_D6;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_DO5;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_DO6;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_D_CY;
  wire [0:0] CLBLM_L_X8Y157_SLICE_X11Y157_D_XOR;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_A;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_A1;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_A2;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_A3;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_A4;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_A5;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_A6;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_AO5;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_AO6;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_AQ;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_A_CY;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_A_XOR;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_B;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_B1;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_B2;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_B3;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_B4;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_B5;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_B6;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_BO5;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_BO6;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_BQ;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_B_CY;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_B_XOR;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_C;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_C1;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_C2;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_C3;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_C4;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_C5;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_C6;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_CLK;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_CO5;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_CO6;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_C_CY;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_C_XOR;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_D;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_D1;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_D2;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_D3;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_D4;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_D5;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_D6;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_DO5;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_DO6;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_D_CY;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X10Y158_D_XOR;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_A;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_A1;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_A2;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_A3;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_A4;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_A5;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_A6;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_AO5;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_AO6;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_AQ;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_A_CY;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_A_XOR;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_B;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_B1;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_B2;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_B3;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_B4;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_B5;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_B6;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_BO5;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_BO6;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_BQ;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_B_CY;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_B_XOR;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_C;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_C1;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_C2;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_C3;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_C4;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_C5;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_C6;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_CLK;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_CO5;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_CO6;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_C_CY;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_C_XOR;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_D;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_D1;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_D2;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_D3;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_D4;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_D5;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_D6;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_DO5;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_DO6;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_D_CY;
  wire [0:0] CLBLM_L_X8Y158_SLICE_X11Y158_D_XOR;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_A;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_A1;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_A2;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_A3;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_A4;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_A5;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_A6;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_AO5;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_AO6;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_AQ;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_A_CY;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_A_XOR;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_B;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_B1;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_B2;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_B3;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_B4;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_B5;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_B6;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_BMUX;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_BO5;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_BO6;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_B_CY;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_B_XOR;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_C;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_C1;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_C2;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_C3;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_C4;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_C5;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_C6;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_CLK;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_CO5;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_CO6;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_C_CY;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_C_XOR;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_D;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_D1;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_D2;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_D3;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_D4;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_D5;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_D6;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_DO5;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_DO6;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_D_CY;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X10Y159_D_XOR;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_A;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_A1;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_A2;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_A3;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_A4;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_A5;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_A6;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_AO5;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_AO6;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_A_CY;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_A_XOR;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_B;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_B1;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_B2;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_B3;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_B4;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_B5;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_B6;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_BO5;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_BO6;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_B_CY;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_B_XOR;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_C;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_C1;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_C2;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_C3;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_C4;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_C5;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_C6;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_CO5;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_CO6;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_C_CY;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_C_XOR;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_D;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_D1;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_D2;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_D3;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_D4;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_D5;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_D6;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_DO5;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_DO6;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_D_CY;
  wire [0:0] CLBLM_L_X8Y159_SLICE_X11Y159_D_XOR;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_A;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_A1;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_A2;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_A3;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_A4;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_A5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_A6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_AO5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_AO6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_A_CY;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_A_XOR;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_B;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_B1;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_B2;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_B3;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_B4;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_B5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_B6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_BO5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_BO6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_B_CY;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_B_XOR;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_C;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_C1;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_C2;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_C3;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_C4;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_C5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_C6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_CO5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_CO6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_C_CY;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_C_XOR;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_D;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_D1;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_D2;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_D3;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_D4;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_D5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_D6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_DO5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_DO6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_D_CY;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X162Y141_D_XOR;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_A;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_A1;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_A2;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_A3;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_A4;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_A5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_A6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_AMUX;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_AO5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_AO6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_A_CY;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_A_XOR;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_B;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_B1;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_B2;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_B3;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_B4;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_B5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_B6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_BO5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_BO6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_B_CY;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_B_XOR;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_C;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_C1;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_C2;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_C3;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_C4;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_C5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_C6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_CO5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_CO6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_C_CY;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_C_XOR;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_D;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_D1;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_D2;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_D3;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_D4;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_D5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_D6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_DO5;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_DO6;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_D_CY;
  wire [0:0] CLBLM_R_X103Y141_SLICE_X163Y141_D_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_AO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_AO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_A_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_BO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_BO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_B_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_CO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_CO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_C_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_DO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_DO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X162Y169_D_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_AMUX;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_A_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_BO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_BO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_B_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_CO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_CO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_C_XOR;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D1;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D2;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D3;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D4;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_DO5;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_DO6;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D_CY;
  wire [0:0] CLBLM_R_X103Y169_SLICE_X163Y169_D_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_AO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_AO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_A_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_BO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_BO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_B_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_CO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_CO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_C_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_DO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_DO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X162Y172_D_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_AMUX;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_A_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_BO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_BO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_B_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_CO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_CO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_C_XOR;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D1;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D2;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D3;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D4;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_DO5;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_DO6;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D_CY;
  wire [0:0] CLBLM_R_X103Y172_SLICE_X163Y172_D_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_AO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_AO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_A_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_BO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_BO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_B_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_CO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_CO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_C_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_DO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_DO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X162Y174_D_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_AMUX;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_A_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_BO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_BO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_B_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_CO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_CO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_C_XOR;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D1;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D2;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D3;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D4;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_DO5;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_DO6;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D_CY;
  wire [0:0] CLBLM_R_X103Y174_SLICE_X163Y174_D_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_AO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_AO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_A_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_BO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_BO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_B_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_CO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_CO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_C_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_DO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_DO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X162Y177_D_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AMUX;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_A_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_BO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_BO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_B_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_CO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_CO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_C_XOR;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D1;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D2;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D3;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D4;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_DO5;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_DO6;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D_CY;
  wire [0:0] CLBLM_R_X103Y177_SLICE_X163Y177_D_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_AO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_AO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_A_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_BO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_BO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_B_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_CO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_C_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_DO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X14Y144_D_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A5Q;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_AMUX;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_AO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_AO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_AQ;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_A_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_BO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_BO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_B_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_CLK;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_CO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_CO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_C_XOR;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D1;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D2;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D3;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D4;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_DO5;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_DO6;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D_CY;
  wire [0:0] CLBLM_R_X11Y144_SLICE_X15Y144_D_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_AO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_AO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_A_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_BO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_BO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_BQ;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_B_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_CLK;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_CO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_CO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_CQ;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_C_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_DO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_DO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_DQ;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X14Y146_D_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_AO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_AO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_AQ;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_A_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_BO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_BO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_BQ;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_B_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_CLK;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_CO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_CO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_CQ;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_C_XOR;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D1;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D2;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D3;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D4;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_DMUX;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_DO5;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_DO6;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D_CY;
  wire [0:0] CLBLM_R_X11Y146_SLICE_X15Y146_D_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_AMUX;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_AO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_AO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_A_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_BO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_BO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_B_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_CO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_C_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_DO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_DO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X14Y147_D_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_AO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_AO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_A_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_BMUX;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_BO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_BO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_B_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_CO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_CO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_C_XOR;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D1;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D2;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D3;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D4;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_DO5;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_DO6;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D_CY;
  wire [0:0] CLBLM_R_X11Y147_SLICE_X15Y147_D_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_AO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_AQ;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_A_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_BO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_BO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_BQ;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_B_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_CLK;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_CO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_CO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_CQ;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_C_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_DO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_DO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X14Y148_D_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_AO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_AO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_AQ;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_A_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_BO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_BO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_B_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_CLK;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_CO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_CO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_C_XOR;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D1;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D2;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D3;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D4;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_DO5;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_DO6;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D_CY;
  wire [0:0] CLBLM_R_X11Y148_SLICE_X15Y148_D_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_AO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_AO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_A_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_BO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_BO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_BQ;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_B_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_CLK;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_CO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_CO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_C_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_DO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_DO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_DQ;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X14Y149_D_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A5Q;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_AMUX;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_AO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_AO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_AQ;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_A_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_BO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_BO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_B_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_CLK;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_CO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_CO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_C_XOR;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D1;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D2;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D3;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D4;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_DMUX;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_DO5;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D_CY;
  wire [0:0] CLBLM_R_X11Y149_SLICE_X15Y149_D_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_AO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_AO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_AQ;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_A_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_BMUX;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_BO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_BO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_B_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_CLK;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_CO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_CO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_C_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_DO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_DO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X14Y150_D_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_AMUX;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_AO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_AO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_A_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_BO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_BO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_B_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_CO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_CO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_C_XOR;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D1;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D2;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D3;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D4;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_DO5;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_DO6;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D_CY;
  wire [0:0] CLBLM_R_X11Y150_SLICE_X15Y150_D_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_AO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_AO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_AQ;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_A_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_BO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_BO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_BQ;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_B_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_CLK;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_CO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_CO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_C_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_DO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_DO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X14Y151_D_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A5Q;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_AMUX;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_AO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_AO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_AQ;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_A_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_BO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_BO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_BQ;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_B_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_CLK;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_CO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_CO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_C_XOR;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D1;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D2;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D3;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D4;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_DMUX;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_DO5;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_DO6;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D_CY;
  wire [0:0] CLBLM_R_X11Y151_SLICE_X15Y151_D_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_AO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_AO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_AQ;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_A_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B5Q;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_BMUX;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_BO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_BO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_BQ;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_B_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_CLK;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_CO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_CO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_CQ;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_C_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_DMUX;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_DO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_DO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X14Y152_D_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_AO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_AO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_AQ;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_A_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_BO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_BO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_BQ;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_B_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_CLK;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_CO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_CO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_CQ;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_C_XOR;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D1;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D2;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D3;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D4;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_DO5;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_DO6;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_DQ;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D_CY;
  wire [0:0] CLBLM_R_X11Y152_SLICE_X15Y152_D_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_AO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_AO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_AQ;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_A_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_BO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_BO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_B_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_CLK;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_CO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_CO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_C_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_DO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_DO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X14Y153_D_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_AO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_AO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_AQ;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_A_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_BO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_BO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_BQ;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_B_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_CLK;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_CO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_CO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_CQ;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_C_XOR;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D1;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D2;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D3;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D4;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_DO5;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_DO6;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_DQ;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D_CY;
  wire [0:0] CLBLM_R_X11Y153_SLICE_X15Y153_D_XOR;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_A;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_A1;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_A2;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_A3;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_A4;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_A5;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_A6;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_AO5;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_AO6;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_AQ;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_A_CY;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_A_XOR;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_B;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_B1;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_B2;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_B3;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_B4;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_B5;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_B6;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_BMUX;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_BO5;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_BO6;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_B_CY;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_B_XOR;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_C;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_C1;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_C2;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_C3;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_C4;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_C5;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_C6;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_CLK;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_CO5;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_CO6;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_CQ;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_C_CY;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_C_XOR;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_D;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_D1;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_D2;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_D3;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_D4;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_D5;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_D5Q;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_D6;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_DMUX;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_DO5;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_DO6;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_DQ;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_D_CY;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X14Y154_D_XOR;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_A;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_A1;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_A2;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_A3;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_A4;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_A5;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_A6;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_AO5;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_AO6;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_AQ;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_A_CY;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_A_XOR;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_B;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_B1;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_B2;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_B3;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_B4;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_B5;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_B6;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_BO5;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_BO6;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_BQ;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_B_CY;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_B_XOR;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_C;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_C1;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_C2;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_C3;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_C4;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_C5;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_C6;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_CLK;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_CMUX;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_CO5;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_CO6;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_C_CY;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_C_XOR;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_D;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_D1;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_D2;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_D3;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_D4;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_D5;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_D6;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_DO5;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_DO6;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_D_CY;
  wire [0:0] CLBLM_R_X11Y154_SLICE_X15Y154_D_XOR;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_A;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_A1;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_A2;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_A3;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_A4;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_A5;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_A6;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_AO5;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_AO6;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_AQ;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_A_CY;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_A_XOR;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_B;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_B1;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_B2;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_B3;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_B4;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_B5;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_B6;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_BO5;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_BO6;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_BQ;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_B_CY;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_B_XOR;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_C;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_C1;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_C2;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_C3;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_C4;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_C5;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_C6;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_CLK;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_CO5;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_CO6;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_CQ;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_C_CY;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_C_XOR;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_D;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_D1;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_D2;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_D3;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_D4;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_D5;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_D6;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_DO5;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_DO6;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_DQ;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_D_CY;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X14Y155_D_XOR;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_A;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_A1;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_A2;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_A3;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_A4;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_A5;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_A6;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_AO5;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_AO6;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_AQ;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_A_CY;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_A_XOR;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_B;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_B1;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_B2;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_B3;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_B4;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_B5;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_B6;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_BO5;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_BO6;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_B_CY;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_B_XOR;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_C;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_C1;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_C2;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_C3;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_C4;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_C5;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_C6;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_CLK;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_CO5;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_CO6;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_C_CY;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_C_XOR;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_D;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_D1;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_D2;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_D3;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_D4;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_D5;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_D6;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_DMUX;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_DO5;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_DO6;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_D_CY;
  wire [0:0] CLBLM_R_X11Y155_SLICE_X15Y155_D_XOR;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_A;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_A1;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_A2;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_A3;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_A4;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_A5;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_A6;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_AO5;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_AO6;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_AQ;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_A_CY;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_A_XOR;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_B;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_B1;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_B2;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_B3;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_B4;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_B5;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_B6;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_BO5;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_BO6;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_BQ;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_B_CY;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_B_XOR;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_C;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_C1;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_C2;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_C3;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_C4;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_C5;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_C6;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_CLK;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_CO5;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_CO6;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_C_CY;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_C_XOR;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_D;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_D1;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_D2;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_D3;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_D4;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_D5;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_D6;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_DO5;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_DO6;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_D_CY;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X14Y156_D_XOR;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_A;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_A1;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_A2;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_A3;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_A4;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_A5;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_A6;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_AO5;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_AO6;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_AQ;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_A_CY;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_A_XOR;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_B;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_B1;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_B2;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_B3;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_B4;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_B5;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_B6;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_BO5;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_BO6;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_BQ;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_B_CY;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_B_XOR;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_C;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_C1;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_C2;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_C3;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_C4;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_C5;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_C6;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_CLK;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_CO5;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_CO6;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_C_CY;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_C_XOR;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_D;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_D1;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_D2;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_D3;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_D4;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_D5;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_D6;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_DO5;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_DO6;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_D_CY;
  wire [0:0] CLBLM_R_X11Y156_SLICE_X15Y156_D_XOR;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_A;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_A1;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_A2;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_A3;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_A4;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_A5;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_A6;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_AO5;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_AO6;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_AQ;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_A_CY;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_A_XOR;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_B;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_B1;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_B2;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_B3;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_B4;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_B5;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_B6;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_BO5;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_BO6;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_BQ;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_B_CY;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_B_XOR;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_C;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_C1;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_C2;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_C3;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_C4;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_C5;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_C6;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_CLK;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_CO5;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_CO6;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_CQ;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_C_CY;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_C_XOR;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_D;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_D1;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_D2;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_D3;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_D4;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_D5;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_D6;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_DO5;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_DO6;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_D_CY;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X14Y157_D_XOR;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_A;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_A1;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_A2;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_A3;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_A4;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_A5;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_A6;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_AO5;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_AO6;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_AQ;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_A_CY;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_A_XOR;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_B;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_B1;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_B2;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_B3;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_B4;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_B5;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_B6;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_BO5;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_BO6;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_BQ;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_B_CY;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_B_XOR;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_C;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_C1;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_C2;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_C3;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_C4;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_C5;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_C6;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_CLK;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_CO5;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_CO6;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_C_CY;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_C_XOR;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_D;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_D1;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_D2;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_D3;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_D4;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_D5;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_D6;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_DO5;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_DO6;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_D_CY;
  wire [0:0] CLBLM_R_X11Y157_SLICE_X15Y157_D_XOR;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_A;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_A1;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_A2;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_A3;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_A4;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_A5;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_A6;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_AO5;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_AO6;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_AQ;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_A_CY;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_A_XOR;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_B;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_B1;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_B2;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_B3;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_B4;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_B5;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_B6;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_BO5;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_BO6;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_BQ;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_B_CY;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_B_XOR;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_C;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_C1;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_C2;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_C3;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_C4;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_C5;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_C6;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_CLK;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_CO5;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_CO6;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_CQ;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_C_CY;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_C_XOR;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_D;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_D1;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_D2;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_D3;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_D4;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_D5;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_D6;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_DMUX;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_DO5;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_DO6;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_D_CY;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X14Y158_D_XOR;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_A;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_A1;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_A2;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_A3;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_A4;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_A5;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_A6;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_AO5;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_AO6;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_AQ;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_A_CY;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_A_XOR;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_B;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_B1;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_B2;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_B3;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_B4;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_B5;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_B6;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_BMUX;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_BO5;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_BO6;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_B_CY;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_B_XOR;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_C;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_C1;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_C2;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_C3;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_C4;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_C5;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_C6;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_CLK;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_CO5;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_CO6;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_C_CY;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_C_XOR;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_D;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_D1;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_D2;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_D3;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_D4;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_D5;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_D6;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_DO5;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_DO6;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_D_CY;
  wire [0:0] CLBLM_R_X11Y158_SLICE_X15Y158_D_XOR;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_A;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_A1;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_A2;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_A3;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_A4;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_A5;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_A6;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_AO5;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_AO6;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_AQ;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_A_CY;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_A_XOR;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_B;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_B1;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_B2;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_B3;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_B4;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_B5;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_B6;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_BO5;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_BO6;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_BQ;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_B_CY;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_B_XOR;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_C;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_C1;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_C2;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_C3;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_C4;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_C5;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_C6;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_CLK;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_CO5;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_CO6;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_CQ;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_C_CY;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_C_XOR;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_D;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_D1;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_D2;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_D3;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_D4;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_D5;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_D6;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_DO5;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_DO6;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_DQ;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_D_CY;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X14Y159_D_XOR;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_A;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_A1;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_A2;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_A3;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_A4;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_A5;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_A6;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_AO5;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_AO6;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_AQ;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_A_CY;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_A_XOR;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_B;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_B1;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_B2;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_B3;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_B4;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_B5;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_B6;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_BO5;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_BO6;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_BQ;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_B_CY;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_B_XOR;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_C;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_C1;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_C2;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_C3;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_C4;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_C5;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_C6;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_CLK;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_CMUX;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_CO5;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_CO6;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_C_CY;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_C_XOR;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_D;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_D1;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_D2;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_D3;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_D4;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_D5;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_D6;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_DMUX;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_DO5;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_DO6;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_D_CY;
  wire [0:0] CLBLM_R_X11Y159_SLICE_X15Y159_D_XOR;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_A;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_A1;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_A2;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_A3;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_A4;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_A5;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_A6;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_AO5;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_AO6;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_AQ;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_A_CY;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_A_XOR;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_B;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_B1;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_B2;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_B3;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_B4;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_B5;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_B6;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_BO5;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_BO6;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_B_CY;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_B_XOR;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_C;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_C1;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_C2;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_C3;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_C4;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_C5;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_C6;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_CLK;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_CO5;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_CO6;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_C_CY;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_C_XOR;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_D;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_D1;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_D2;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_D3;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_D4;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_D5;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_D6;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_DO5;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_DO6;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_D_CY;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X14Y160_D_XOR;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_A;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_A1;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_A2;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_A3;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_A4;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_A5;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_A6;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_AO5;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_AO6;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_A_CY;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_A_XOR;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_B;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_B1;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_B2;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_B3;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_B4;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_B5;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_B6;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_BO5;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_BO6;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_B_CY;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_B_XOR;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_C;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_C1;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_C2;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_C3;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_C4;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_C5;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_C6;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_CO5;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_CO6;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_C_CY;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_C_XOR;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_D;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_D1;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_D2;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_D3;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_D4;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_D5;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_D6;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_DO5;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_DO6;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_D_CY;
  wire [0:0] CLBLM_R_X11Y160_SLICE_X15Y160_D_XOR;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_A;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_A1;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_A2;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_A3;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_A4;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_A5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_A6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_AMUX;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_AO5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_AO6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_A_CY;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_A_XOR;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_B;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_B1;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_B2;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_B3;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_B4;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_B5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_B6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_BMUX;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_BO5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_BO6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_B_CY;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_B_XOR;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_C;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_C1;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_C2;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_C3;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_C4;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_C5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_C6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_CO5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_CO6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_C_CY;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_C_XOR;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_D;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_D1;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_D2;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_D3;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_D4;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_D5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_D6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_DO5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_DO6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_D_CY;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X18Y147_D_XOR;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_A;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_A1;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_A2;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_A3;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_A4;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_A5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_A6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_AO5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_AO6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_A_CY;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_A_XOR;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_B;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_B1;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_B2;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_B3;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_B4;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_B5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_B6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_BO5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_BO6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_B_CY;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_B_XOR;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_C;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_C1;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_C2;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_C3;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_C4;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_C5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_C6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_CO5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_CO6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_C_CY;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_C_XOR;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_D;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_D1;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_D2;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_D3;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_D4;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_D5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_D6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_DO5;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_DO6;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_D_CY;
  wire [0:0] CLBLM_R_X13Y147_SLICE_X19Y147_D_XOR;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_A;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_A1;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_A2;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_A3;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_A4;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_A5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_A6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_AMUX;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_AO5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_AO6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_AQ;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_A_CY;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_A_XOR;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_B;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_B1;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_B2;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_B3;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_B4;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_B5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_B6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_BMUX;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_BO5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_BO6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_B_CY;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_B_XOR;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_C;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_C1;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_C2;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_C3;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_C4;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_C5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_C6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_CLK;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_CMUX;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_CO5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_CO6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_C_CY;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_C_XOR;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_D;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_D1;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_D2;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_D3;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_D4;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_D5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_D6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_DO5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_DO6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_D_CY;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X18Y148_D_XOR;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_A;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_A1;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_A2;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_A3;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_A4;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_A5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_A6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_AO5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_AO6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_A_CY;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_A_XOR;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_B;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_B1;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_B2;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_B3;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_B4;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_B5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_B6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_BO5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_BO6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_B_CY;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_B_XOR;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_C;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_C1;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_C2;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_C3;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_C4;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_C5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_C6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_CO5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_CO6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_C_CY;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_C_XOR;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_D;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_D1;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_D2;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_D3;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_D4;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_D5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_D6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_DO5;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_DO6;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_D_CY;
  wire [0:0] CLBLM_R_X13Y148_SLICE_X19Y148_D_XOR;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A1;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A2;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A3;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A4;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A5Q;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_AMUX;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_AO5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_AO6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_AQ;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_AX;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A_CY;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_A_XOR;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B1;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B2;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B3;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B4;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_BO5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_BO6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_BQ;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B_CY;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_B_XOR;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C1;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C2;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C3;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C4;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_CLK;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_CO5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_CO6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_CQ;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C_CY;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_C_XOR;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D1;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D2;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D3;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D4;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_DO5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_DO6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D_CY;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X18Y149_D_XOR;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A1;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A2;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A3;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A4;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A5Q;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_AMUX;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_AO5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_AO6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_AQ;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A_CY;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_A_XOR;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B1;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B2;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B3;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B4;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_BMUX;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_BO5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_BO6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B_CY;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_B_XOR;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C1;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C2;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C3;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C4;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_CLK;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_CO5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_CO6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_CQ;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C_CY;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_C_XOR;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D1;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D2;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D3;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D4;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_DO5;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_DO6;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D_CY;
  wire [0:0] CLBLM_R_X13Y149_SLICE_X19Y149_D_XOR;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_A;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_A1;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_A2;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_A3;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_A4;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_A5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_A6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_AO5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_AO6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_AQ;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_A_CY;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_A_XOR;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_B;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_B1;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_B2;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_B3;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_B4;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_B5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_B6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_BO5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_BO6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_BQ;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_B_CY;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_B_XOR;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_C;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_C1;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_C2;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_C3;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_C4;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_C5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_C6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_CLK;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_CO5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_CO6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_CQ;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_C_CY;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_C_XOR;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_D;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_D1;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_D2;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_D3;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_D4;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_D5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_D6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_DMUX;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_DO5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_DO6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_D_CY;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X18Y150_D_XOR;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_A;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_A1;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_A2;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_A3;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_A4;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_A5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_A6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_AO5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_AO6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_AQ;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_A_CY;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_A_XOR;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_B;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_B1;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_B2;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_B3;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_B4;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_B5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_B6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_BO5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_BO6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_B_CY;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_B_XOR;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_C;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_C1;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_C2;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_C3;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_C4;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_C5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_C6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_CLK;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_CO5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_CO6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_C_CY;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_C_XOR;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_D;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_D1;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_D2;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_D3;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_D4;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_D5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_D6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_DO5;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_DO6;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_D_CY;
  wire [0:0] CLBLM_R_X13Y150_SLICE_X19Y150_D_XOR;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_A;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_A1;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_A2;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_A3;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_A4;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_A5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_A6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_AO5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_AO6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_AQ;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_A_CY;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_A_XOR;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_B;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_B1;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_B2;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_B3;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_B4;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_B5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_B6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_BO5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_BO6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_BQ;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_B_CY;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_B_XOR;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_C;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_C1;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_C2;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_C3;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_C4;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_C5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_C6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_CLK;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_CO5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_CO6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_CQ;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_C_CY;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_C_XOR;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_D;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_D1;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_D2;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_D3;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_D4;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_D5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_D6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_DO5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_DO6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_DQ;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_D_CY;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X18Y151_D_XOR;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_A;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_A1;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_A2;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_A3;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_A4;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_A5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_A6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_AO5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_AO6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_A_CY;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_A_XOR;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_B;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_B1;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_B2;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_B3;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_B4;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_B5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_B6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_BO5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_BO6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_B_CY;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_B_XOR;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_C;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_C1;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_C2;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_C3;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_C4;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_C5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_C6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_CO5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_CO6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_C_CY;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_C_XOR;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_D;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_D1;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_D2;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_D3;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_D4;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_D5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_D6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_DO5;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_DO6;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_D_CY;
  wire [0:0] CLBLM_R_X13Y151_SLICE_X19Y151_D_XOR;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_A;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_A1;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_A2;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_A3;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_A4;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_A5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_A5Q;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_A6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_AMUX;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_AO5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_AO6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_AQ;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_AX;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_A_CY;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_A_XOR;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_B;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_B1;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_B2;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_B3;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_B4;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_B5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_B6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_BMUX;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_BO5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_BO6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_B_CY;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_B_XOR;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_C;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_C1;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_C2;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_C3;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_C4;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_C5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_C6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_CLK;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_CO5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_CO6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_CQ;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_C_CY;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_C_XOR;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_D;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_D1;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_D2;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_D3;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_D4;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_D5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_D6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_DO5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_DO6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_D_CY;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X18Y152_D_XOR;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_A;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_A1;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_A2;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_A3;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_A4;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_A5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_A6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_AO5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_AO6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_AQ;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_A_CY;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_A_XOR;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_B;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_B1;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_B2;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_B3;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_B4;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_B5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_B6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_BO5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_BO6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_BQ;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_B_CY;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_B_XOR;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_C;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_C1;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_C2;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_C3;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_C4;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_C5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_C6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_CLK;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_CO5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_CO6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_C_CY;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_C_XOR;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_D;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_D1;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_D2;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_D3;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_D4;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_D5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_D6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_DO5;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_DO6;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_D_CY;
  wire [0:0] CLBLM_R_X13Y152_SLICE_X19Y152_D_XOR;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_A;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_A1;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_A2;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_A3;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_A4;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_A5;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_A6;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_AO5;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_AO6;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_AQ;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_A_CY;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_A_XOR;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_B;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_B1;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_B2;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_B3;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_B4;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_B5;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_B6;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_BO5;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_BO6;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_BQ;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_B_CY;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_B_XOR;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_C;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_C1;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_C2;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_C3;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_C4;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_C5;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_C5Q;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_C6;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_CLK;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_CMUX;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_CO5;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_CO6;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_CQ;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_C_CY;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_C_XOR;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_D;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_D1;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_D2;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_D3;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_D4;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_D5;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_D6;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_DO5;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_DO6;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_DQ;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_D_CY;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X18Y153_D_XOR;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_A;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_A1;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_A2;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_A3;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_A4;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_A5;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_A6;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_AO5;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_AO6;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_AQ;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_A_CY;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_A_XOR;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_B;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_B1;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_B2;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_B3;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_B4;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_B5;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_B6;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_BO5;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_BO6;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_BQ;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_B_CY;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_B_XOR;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_C;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_C1;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_C2;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_C3;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_C4;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_C5;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_C6;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_CLK;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_CO5;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_CO6;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_CQ;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_C_CY;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_C_XOR;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_D;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_D1;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_D2;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_D3;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_D4;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_D5;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_D6;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_DO5;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_DO6;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_D_CY;
  wire [0:0] CLBLM_R_X13Y153_SLICE_X19Y153_D_XOR;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_A;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_A1;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_A2;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_A3;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_A4;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_A5;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_A6;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_AO5;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_AO6;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_AQ;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_A_CY;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_A_XOR;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_B;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_B1;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_B2;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_B3;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_B4;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_B5;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_B6;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_BO5;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_BO6;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_BQ;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_B_CY;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_B_XOR;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_C;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_C1;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_C2;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_C3;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_C4;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_C5;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_C6;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_CLK;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_CO5;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_CO6;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_CQ;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_C_CY;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_C_XOR;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_D;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_D1;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_D2;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_D3;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_D4;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_D5;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_D6;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_DO5;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_DO6;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_D_CY;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X18Y154_D_XOR;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_A;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_A1;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_A2;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_A3;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_A4;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_A5;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_A6;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_AO5;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_AO6;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_AQ;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_A_CY;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_A_XOR;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_B;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_B1;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_B2;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_B3;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_B4;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_B5;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_B6;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_BO5;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_BO6;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_B_CY;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_B_XOR;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_C;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_C1;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_C2;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_C3;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_C4;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_C5;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_C6;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_CLK;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_CO5;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_CO6;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_C_CY;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_C_XOR;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_D;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_D1;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_D2;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_D3;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_D4;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_D5;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_D6;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_DO5;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_DO6;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_D_CY;
  wire [0:0] CLBLM_R_X13Y154_SLICE_X19Y154_D_XOR;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_A;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_A1;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_A2;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_A3;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_A4;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_A5;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_A6;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_AO5;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_AO6;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_AQ;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_A_CY;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_A_XOR;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_B;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_B1;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_B2;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_B3;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_B4;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_B5;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_B6;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_BO5;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_BO6;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_BQ;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_B_CY;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_B_XOR;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_C;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_C1;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_C2;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_C3;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_C4;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_C5;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_C6;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_CLK;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_CMUX;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_CO5;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_CO6;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_C_CY;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_C_XOR;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_D;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_D1;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_D2;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_D3;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_D4;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_D5;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_D6;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_DMUX;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_DO5;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_DO6;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_D_CY;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X18Y155_D_XOR;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_A;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_A1;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_A2;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_A3;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_A4;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_A5;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_A6;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_AO5;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_AO6;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_A_CY;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_A_XOR;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_B;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_B1;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_B2;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_B3;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_B4;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_B5;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_B6;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_BO5;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_BO6;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_B_CY;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_B_XOR;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_C;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_C1;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_C2;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_C3;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_C4;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_C5;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_C6;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_CO5;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_CO6;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_C_CY;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_C_XOR;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_D;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_D1;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_D2;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_D3;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_D4;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_D5;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_D6;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_DO5;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_DO6;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_D_CY;
  wire [0:0] CLBLM_R_X13Y155_SLICE_X19Y155_D_XOR;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_A;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_A1;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_A2;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_A3;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_A4;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_A5;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_A6;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_AO5;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_AO6;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_AQ;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_A_CY;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_A_XOR;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_B;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_B1;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_B2;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_B3;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_B4;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_B5;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_B6;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_BO5;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_BO6;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_B_CY;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_B_XOR;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_C;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_C1;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_C2;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_C3;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_C4;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_C5;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_C6;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_CLK;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_CO5;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_CO6;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_C_CY;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_C_XOR;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_D;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_D1;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_D2;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_D3;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_D4;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_D5;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_D6;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_DO5;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_DO6;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_D_CY;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X18Y156_D_XOR;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_A;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_A1;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_A2;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_A3;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_A4;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_A5;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_A6;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_AO5;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_AO6;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_AQ;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_A_CY;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_A_XOR;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_B;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_B1;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_B2;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_B3;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_B4;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_B5;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_B6;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_BO5;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_BO6;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_B_CY;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_B_XOR;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_C;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_C1;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_C2;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_C3;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_C4;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_C5;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_C6;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_CLK;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_CO5;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_CO6;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_C_CY;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_C_XOR;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_D;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_D1;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_D2;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_D3;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_D4;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_D5;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_D6;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_DO5;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_DO6;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_D_CY;
  wire [0:0] CLBLM_R_X13Y156_SLICE_X19Y156_D_XOR;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_A;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_A1;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_A2;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_A3;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_A4;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_A5;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_A6;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_AMUX;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_AO5;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_AO6;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_AQ;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_AX;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_A_CY;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_A_XOR;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_B;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_B1;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_B2;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_B3;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_B4;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_B5;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_B6;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_BMUX;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_BO5;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_BO6;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_B_CY;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_B_XOR;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_C;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_C1;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_C2;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_C3;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_C4;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_C5;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_C6;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_CE;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_CLK;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_CMUX;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_CO5;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_CO6;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_C_CY;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_C_XOR;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_D;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_D1;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_D2;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_D3;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_D4;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_D5;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_D6;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_DO5;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_DO6;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_D_CY;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_D_XOR;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X18Y157_SR;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_A;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_A1;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_A2;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_A3;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_A4;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_A5;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_A6;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_AO5;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_AO6;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_AQ;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_A_CY;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_A_XOR;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_B;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_B1;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_B2;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_B3;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_B4;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_B5;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_B6;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_BMUX;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_BO5;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_BO6;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_B_CY;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_B_XOR;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_C;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_C1;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_C2;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_C3;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_C4;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_C5;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_C6;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_CLK;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_CO5;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_CO6;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_C_CY;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_C_XOR;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_D;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_D1;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_D2;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_D3;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_D4;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_D5;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_D6;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_DO5;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_DO6;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_D_CY;
  wire [0:0] CLBLM_R_X13Y157_SLICE_X19Y157_D_XOR;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_A;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_A1;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_A2;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_A3;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_A4;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_A5;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_A6;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_AO5;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_AO6;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_AQ;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_A_CY;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_A_XOR;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_B;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_B1;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_B2;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_B3;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_B4;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_B5;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_B6;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_BO5;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_BO6;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_BQ;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_B_CY;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_B_XOR;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_C;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_C1;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_C2;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_C3;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_C4;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_C5;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_C6;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_CLK;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_CO5;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_CO6;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_C_CY;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_C_XOR;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_D;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_D1;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_D2;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_D3;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_D4;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_D5;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_D6;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_DO5;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_DO6;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_D_CY;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X18Y158_D_XOR;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_A;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_A1;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_A2;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_A3;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_A4;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_A5;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_A6;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_AMUX;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_AO5;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_AO6;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_A_CY;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_A_XOR;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_B;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_B1;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_B2;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_B3;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_B4;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_B5;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_B6;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_BMUX;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_BO5;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_BO6;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_B_CY;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_B_XOR;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_C;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_C1;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_C2;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_C3;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_C4;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_C5;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_C6;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_CO5;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_CO6;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_C_CY;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_C_XOR;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_D;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_D1;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_D2;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_D3;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_D4;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_D5;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_D6;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_DO5;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_DO6;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_D_CY;
  wire [0:0] CLBLM_R_X13Y158_SLICE_X19Y158_D_XOR;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_A;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_A1;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_A2;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_A3;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_A4;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_A5;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_A6;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_AO5;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_AO6;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_A_CY;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_A_XOR;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_B;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_B1;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_B2;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_B3;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_B4;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_B5;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_B6;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_BO5;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_BO6;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_B_CY;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_B_XOR;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_C;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_C1;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_C2;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_C3;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_C4;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_C5;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_C6;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_CO5;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_CO6;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_C_CY;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_C_XOR;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_D;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_D1;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_D2;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_D3;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_D4;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_D5;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_D6;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_DO5;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_DO6;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_D_CY;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X18Y159_D_XOR;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_A;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_A1;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_A2;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_A3;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_A4;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_A5;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_A6;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_AO5;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_AO6;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_A_CY;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_A_XOR;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_B;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_B1;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_B2;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_B3;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_B4;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_B5;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_B6;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_BO5;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_BO6;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_B_CY;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_B_XOR;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_C;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_C1;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_C2;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_C3;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_C4;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_C5;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_C6;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_CO5;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_CO6;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_C_CY;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_C_XOR;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_D;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_D1;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_D2;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_D3;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_D4;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_D5;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_D6;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_DO5;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_DO6;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_D_CY;
  wire [0:0] CLBLM_R_X13Y159_SLICE_X19Y159_D_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_AO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_A_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_BO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_BO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_B_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_CO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_CO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_C_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_DO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_DO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X2Y142_D_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_AO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_AO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_A_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_BO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_BO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_B_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_CO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_CO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_C_XOR;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D1;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D2;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D3;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D4;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_DO5;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_DO6;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D_CY;
  wire [0:0] CLBLM_R_X3Y142_SLICE_X3Y142_D_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A5Q;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_AMUX;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_AO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_AO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_AQ;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_AX;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_A_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_BMUX;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_BO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_BO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_B_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_CLK;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_CO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_CO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_C_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_DO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_DO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X2Y150_D_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_AO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_AQ;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_A_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_BO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_B_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_CLK;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_CO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_CQ;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_C_XOR;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D1;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D2;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D3;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D4;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_DO5;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D_CY;
  wire [0:0] CLBLM_R_X3Y150_SLICE_X3Y150_D_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_AMUX;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_AO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_AO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_AQ;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_A_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_BO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_BO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_BQ;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_B_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_CLK;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_CMUX;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_CO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_CO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_C_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_DO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_DO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X2Y151_D_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_AMUX;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_AO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_AO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_AQ;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_A_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_BMUX;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_BO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_BO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_B_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_CLK;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_CO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_CO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_C_XOR;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D1;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D2;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D3;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D4;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_DO5;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_DO6;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D_CY;
  wire [0:0] CLBLM_R_X3Y151_SLICE_X3Y151_D_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_AMUX;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_AO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_AO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_A_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_BO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_BO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_B_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_CO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_C_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_DMUX;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_DO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X2Y152_D_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_AMUX;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_AO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_AO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_A_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_BMUX;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_BO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_BO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_B_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_CO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_CO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_C_XOR;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D1;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D2;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D3;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D4;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_DO5;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_DO6;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D_CY;
  wire [0:0] CLBLM_R_X3Y152_SLICE_X3Y152_D_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_AMUX;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_AO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_AO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_A_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_BMUX;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_BO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_BO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_B_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_CO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_CO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_C_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_DO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_DO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X2Y153_D_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_AMUX;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_AO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_AO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_A_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_BO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_BO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_B_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_CO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_CO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_C_XOR;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D1;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D2;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D3;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D4;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_DO5;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_DO6;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D_CY;
  wire [0:0] CLBLM_R_X3Y153_SLICE_X3Y153_D_XOR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A1;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A2;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A3;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A4;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_AO5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_AO6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A_CY;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_A_XOR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B1;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B2;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B3;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B4;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_BO5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_BO6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B_CY;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_B_XOR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C1;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C2;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C3;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C4;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_CO5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_CO6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C_CY;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_C_XOR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D1;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D2;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D3;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D4;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_DO5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_DO6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D_CY;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X2Y154_D_XOR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A1;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A2;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A3;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A4;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_AMUX;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_AO5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_AO6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A_CY;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_A_XOR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B1;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B2;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B3;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B4;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_BO5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_BO6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B_CY;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_B_XOR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C1;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C2;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C3;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C4;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_CO5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_CO6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C_CY;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_C_XOR;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D1;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D2;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D3;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D4;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_DO5;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_DO6;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D_CY;
  wire [0:0] CLBLM_R_X3Y154_SLICE_X3Y154_D_XOR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A1;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A2;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A3;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A4;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_AO5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_AO6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A_CY;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_A_XOR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B1;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B2;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B3;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B4;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_BO5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_BO6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B_CY;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_B_XOR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C1;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C2;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C3;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C4;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_CMUX;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_CO5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_CO6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C_CY;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_C_XOR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D1;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D2;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D3;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D4;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_DO5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_DO6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D_CY;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X2Y155_D_XOR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A1;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A2;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A3;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A4;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_AO5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_AO6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A_CY;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_A_XOR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B1;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B2;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B3;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B4;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_BO5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_BO6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B_CY;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_B_XOR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C1;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C2;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C3;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C4;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_CMUX;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_CO5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_CO6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C_CY;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_C_XOR;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D1;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D2;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D3;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D4;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_DMUX;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_DO5;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_DO6;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D_CY;
  wire [0:0] CLBLM_R_X3Y155_SLICE_X3Y155_D_XOR;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_A;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_A1;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_A2;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_A3;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_A4;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_A5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_A6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_AO5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_AO6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_A_CY;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_A_XOR;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_B;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_B1;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_B2;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_B3;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_B4;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_B5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_B6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_BMUX;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_BO5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_BO6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_B_CY;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_B_XOR;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_C;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_C1;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_C2;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_C3;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_C4;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_C5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_C6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_CO5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_CO6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_C_CY;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_C_XOR;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_D;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_D1;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_D2;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_D3;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_D4;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_D5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_D6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_DO5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_DO6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_D_CY;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X2Y156_D_XOR;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_A;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_A1;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_A2;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_A3;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_A4;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_A5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_A6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_AMUX;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_AO5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_AO6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_A_CY;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_A_XOR;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_B;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_B1;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_B2;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_B3;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_B4;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_B5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_B6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_BO5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_BO6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_B_CY;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_B_XOR;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_C;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_C1;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_C2;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_C3;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_C4;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_C5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_C6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_CMUX;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_CO5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_CO6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_C_CY;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_C_XOR;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_D;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_D1;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_D2;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_D3;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_D4;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_D5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_D6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_DO5;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_DO6;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_D_CY;
  wire [0:0] CLBLM_R_X3Y156_SLICE_X3Y156_D_XOR;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_A;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_A1;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_A2;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_A3;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_A4;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_A5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_A6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_AMUX;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_AO5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_AO6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_A_CY;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_A_XOR;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_B;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_B1;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_B2;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_B3;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_B4;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_B5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_B6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_BO5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_BO6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_B_CY;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_B_XOR;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_C;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_C1;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_C2;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_C3;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_C4;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_C5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_C6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_CO5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_CO6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_C_CY;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_C_XOR;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_D;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_D1;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_D2;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_D3;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_D4;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_D5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_D6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_DO5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_DO6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_D_CY;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X2Y157_D_XOR;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_A;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_A1;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_A2;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_A3;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_A4;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_A5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_A6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_AO5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_AO6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_A_CY;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_A_XOR;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_B;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_B1;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_B2;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_B3;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_B4;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_B5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_B6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_BO5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_BO6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_B_CY;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_B_XOR;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_C;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_C1;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_C2;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_C3;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_C4;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_C5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_C6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_CO5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_CO6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_C_CY;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_C_XOR;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_D;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_D1;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_D2;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_D3;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_D4;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_D5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_D6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_DMUX;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_DO5;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_DO6;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_D_CY;
  wire [0:0] CLBLM_R_X3Y157_SLICE_X3Y157_D_XOR;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_A;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_A1;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_A2;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_A3;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_A4;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_A5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_A6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_AMUX;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_AO5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_AO6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_A_CY;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_A_XOR;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_B;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_B1;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_B2;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_B3;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_B4;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_B5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_B6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_BO5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_BO6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_B_CY;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_B_XOR;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_C;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_C1;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_C2;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_C3;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_C4;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_C5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_C6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_CO5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_CO6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_C_CY;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_C_XOR;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_D;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_D1;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_D2;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_D3;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_D4;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_D5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_D6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_DO5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_DO6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_D_CY;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X2Y158_D_XOR;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_A;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_A1;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_A2;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_A3;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_A4;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_A5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_A6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_AO5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_AO6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_A_CY;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_A_XOR;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_B;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_B1;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_B2;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_B3;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_B4;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_B5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_B6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_BO5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_BO6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_B_CY;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_B_XOR;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_C;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_C1;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_C2;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_C3;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_C4;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_C5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_C6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_CO5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_CO6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_C_CY;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_C_XOR;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_D;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_D1;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_D2;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_D3;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_D4;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_D5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_D6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_DO5;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_DO6;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_D_CY;
  wire [0:0] CLBLM_R_X3Y158_SLICE_X3Y158_D_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_AO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_AO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_AQ;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_A_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_BO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_BO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_BQ;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_B_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_CLK;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_CMUX;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_CO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_CO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_C_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_DO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_DO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X6Y144_D_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_AO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_AO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_A_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_BO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_B_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_CO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_CO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_C_XOR;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D1;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D2;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D3;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D4;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_DO5;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_DO6;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D_CY;
  wire [0:0] CLBLM_R_X5Y144_SLICE_X7Y144_D_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A5Q;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_AMUX;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_AO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_AO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_AQ;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_AX;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_A_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_BO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_BO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_BQ;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_B_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_CLK;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_CMUX;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_CO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_C_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_DO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X6Y146_D_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_AO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_AO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_A_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_BO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_BO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_B_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_CO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_CO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_C_XOR;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D1;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D2;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D3;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D4;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_DO5;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_DO6;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D_CY;
  wire [0:0] CLBLM_R_X5Y146_SLICE_X7Y146_D_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_AO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_AO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_A_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_BO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_BO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_BQ;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_B_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_CLK;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_CO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_C_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_DO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_DO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X6Y147_D_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_AO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_AO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_A_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_BO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_BO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_BQ;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_B_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C5Q;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_CLK;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_CMUX;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_CO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_CO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_CQ;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_C_XOR;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D1;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D2;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D3;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D4;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_DO5;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_DO6;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D_CY;
  wire [0:0] CLBLM_R_X5Y147_SLICE_X7Y147_D_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A5Q;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_AMUX;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_AO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_AO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_AQ;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_AX;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_A_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_BO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_BQ;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_B_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_CLK;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_CMUX;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_CO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_CO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_C_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_DO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_DO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X6Y148_D_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A5Q;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_AMUX;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_AO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_AO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_AQ;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_AX;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_A_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B5Q;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_BMUX;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_BO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_BO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_BQ;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_B_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_CLK;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_CO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_CO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_C_XOR;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D1;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D2;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D3;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D4;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_DO5;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_DO6;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D_CY;
  wire [0:0] CLBLM_R_X5Y148_SLICE_X7Y148_D_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A5Q;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_AMUX;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_AO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_AO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_AQ;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_A_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B5Q;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_BMUX;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_BO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_BO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_BQ;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_B_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_CLK;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_CMUX;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_CO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_CO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_C_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_DO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_DO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X6Y149_D_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A5Q;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_AMUX;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_AO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_AO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_AQ;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_AX;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_A_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_BO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_BO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_BQ;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_B_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_CLK;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_CO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_CO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_CQ;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_C_XOR;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D1;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D2;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D3;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D4;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_DMUX;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_DO5;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_DO6;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D_CY;
  wire [0:0] CLBLM_R_X5Y149_SLICE_X7Y149_D_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_AO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_AO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_AQ;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_A_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_BO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_BO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_BQ;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_B_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_CLK;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_CO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_CO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_CQ;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_C_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_DO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_DO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_DQ;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X6Y150_D_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A5Q;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_AMUX;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_AO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_AO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_AQ;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_A_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_BO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_BO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_BQ;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_B_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_CLK;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_CO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_CO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_CQ;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_C_XOR;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D1;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D2;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D3;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D4;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_DO5;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_DO6;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D_CY;
  wire [0:0] CLBLM_R_X5Y150_SLICE_X7Y150_D_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_AO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_AO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_AQ;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_A_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_BO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_BO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_BQ;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_B_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C5Q;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_CLK;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_CMUX;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_CO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_CO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_CQ;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_C_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_DO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_DO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_DQ;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X6Y151_D_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_AO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_AO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_AQ;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_A_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_BO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_BO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_BQ;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_B_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_CLK;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_CO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_CO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_CQ;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_C_XOR;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D1;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D2;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D3;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D4;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_DO5;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_DO6;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_DQ;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D_CY;
  wire [0:0] CLBLM_R_X5Y151_SLICE_X7Y151_D_XOR;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A1;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A2;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A3;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A4;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_AO5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_AO6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_AQ;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A_CY;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_A_XOR;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B1;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B2;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B3;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B4;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_BO5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_BO6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_BQ;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B_CY;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_B_XOR;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C1;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C2;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C3;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C4;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_CLK;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_CMUX;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_CO5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_CO6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C_CY;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_C_XOR;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D1;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D2;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D3;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D4;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_DMUX;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_DO5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_DO6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D_CY;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X6Y152_D_XOR;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A1;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A2;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A3;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A4;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_AO5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_AO6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_AQ;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A_CY;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_A_XOR;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B1;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B2;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B3;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B4;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_BO5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_BO6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_BQ;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B_CY;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_B_XOR;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C1;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C2;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C3;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C4;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_CLK;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_CO5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_CO6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_CQ;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C_CY;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_C_XOR;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D1;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D2;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D3;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D4;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_DO5;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_DO6;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_DQ;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D_CY;
  wire [0:0] CLBLM_R_X5Y152_SLICE_X7Y152_D_XOR;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A1;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A2;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A3;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A4;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_AO5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_AO6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_AQ;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A_CY;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_A_XOR;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B1;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B2;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B3;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B4;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_BMUX;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_BO5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_BO6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B_CY;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_B_XOR;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C1;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C2;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C3;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C4;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_CLK;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_CO5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_CO6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C_CY;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_C_XOR;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D1;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D2;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D3;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D4;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_DMUX;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_DO5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_DO6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D_CY;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X6Y153_D_XOR;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A1;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A2;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A3;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A4;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_AO5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_AO6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_AQ;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A_CY;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_A_XOR;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B1;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B2;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B3;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B4;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_BO5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_BO6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B_CY;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_B_XOR;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C1;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C2;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C3;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C4;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_CLK;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_CMUX;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_CO5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_CO6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C_CY;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_C_XOR;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D1;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D2;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D3;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D4;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_DO5;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_DO6;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D_CY;
  wire [0:0] CLBLM_R_X5Y153_SLICE_X7Y153_D_XOR;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A1;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A2;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A3;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A4;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_AO5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_AO6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_AQ;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A_CY;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_A_XOR;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B1;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B2;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B3;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B4;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_BO5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_BO6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B_CY;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_B_XOR;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C1;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C2;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C3;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C4;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_CLK;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_CO5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_CO6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C_CY;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_C_XOR;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D1;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D2;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D3;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D4;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_DO5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_DO6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D_CY;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X6Y154_D_XOR;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A1;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A2;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A3;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A4;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_AO5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_AO6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_AQ;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A_CY;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_A_XOR;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B1;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B2;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B3;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B4;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_BO5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_BO6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B_CY;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_B_XOR;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C1;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C2;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C3;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C4;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_CLK;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_CO5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_CO6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C_CY;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_C_XOR;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D1;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D2;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D3;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D4;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_DO5;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_DO6;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D_CY;
  wire [0:0] CLBLM_R_X5Y154_SLICE_X7Y154_D_XOR;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_A;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_A1;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_A2;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_A3;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_A4;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_A5;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_A6;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_AO5;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_AO6;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_AQ;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_A_CY;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_A_XOR;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_B;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_B1;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_B2;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_B3;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_B4;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_B5;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_B6;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_BO5;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_BO6;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_B_CY;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_B_XOR;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_C;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_C1;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_C2;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_C3;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_C4;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_C5;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_C6;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_CLK;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_CO5;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_CO6;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_C_CY;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_C_XOR;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_D;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_D1;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_D2;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_D3;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_D4;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_D5;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_D6;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_DO5;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_DO6;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_D_CY;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X6Y155_D_XOR;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_A;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_A1;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_A2;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_A3;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_A4;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_A5;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_A6;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_AO5;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_AO6;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_AQ;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_A_CY;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_A_XOR;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_B;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_B1;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_B2;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_B3;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_B4;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_B5;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_B6;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_BO5;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_BO6;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_BQ;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_B_CY;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_B_XOR;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_C;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_C1;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_C2;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_C3;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_C4;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_C5;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_C6;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_CLK;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_CO5;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_CO6;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_C_CY;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_C_XOR;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_D;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_D1;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_D2;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_D3;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_D4;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_D5;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_D6;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_DMUX;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_DO5;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_DO6;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_D_CY;
  wire [0:0] CLBLM_R_X5Y155_SLICE_X7Y155_D_XOR;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_A;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_A1;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_A2;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_A3;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_A4;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_A5;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_A6;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_AO5;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_AO6;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_A_CY;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_A_XOR;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_B;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_B1;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_B2;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_B3;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_B4;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_B5;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_B6;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_BO5;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_BO6;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_B_CY;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_B_XOR;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_C;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_C1;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_C2;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_C3;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_C4;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_C5;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_C6;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_CO5;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_CO6;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_C_CY;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_C_XOR;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_D;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_D1;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_D2;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_D3;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_D4;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_D5;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_D6;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_DO5;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_DO6;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_D_CY;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X6Y156_D_XOR;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_A;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_A1;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_A2;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_A3;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_A4;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_A5;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_A6;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_AO5;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_AO6;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_AQ;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_A_CY;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_A_XOR;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_B;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_B1;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_B2;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_B3;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_B4;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_B5;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_B6;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_BO5;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_BO6;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_B_CY;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_B_XOR;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_C;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_C1;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_C2;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_C3;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_C4;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_C5;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_C6;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_CLK;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_CO5;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_CO6;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_C_CY;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_C_XOR;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_D;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_D1;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_D2;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_D3;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_D4;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_D5;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_D6;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_DO5;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_DO6;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_D_CY;
  wire [0:0] CLBLM_R_X5Y156_SLICE_X7Y156_D_XOR;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_A;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_A1;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_A2;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_A3;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_A4;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_A5;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_A6;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_AO5;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_AO6;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_AQ;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_A_CY;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_A_XOR;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_B;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_B1;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_B2;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_B3;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_B4;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_B5;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_B6;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_BMUX;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_BO5;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_BO6;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_B_CY;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_B_XOR;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_C;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_C1;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_C2;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_C3;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_C4;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_C5;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_C6;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_CLK;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_CO5;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_CO6;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_C_CY;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_C_XOR;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_D;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_D1;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_D2;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_D3;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_D4;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_D5;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_D6;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_DO5;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_DO6;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_D_CY;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X6Y157_D_XOR;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_A;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_A1;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_A2;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_A3;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_A4;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_A5;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_A6;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_AO5;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_AO6;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_AQ;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_A_CY;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_A_XOR;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_B;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_B1;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_B2;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_B3;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_B4;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_B5;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_B6;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_BO5;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_BO6;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_BQ;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_B_CY;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_B_XOR;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_C;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_C1;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_C2;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_C3;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_C4;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_C5;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_C6;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_CLK;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_CO5;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_CO6;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_CQ;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_C_CY;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_C_XOR;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_D;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_D1;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_D2;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_D3;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_D4;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_D5;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_D6;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_DO5;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_DO6;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_DQ;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_D_CY;
  wire [0:0] CLBLM_R_X5Y157_SLICE_X7Y157_D_XOR;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_A;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_A1;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_A2;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_A3;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_A4;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_A5;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_A6;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_AO5;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_AO6;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_AQ;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_A_CY;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_A_XOR;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_B;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_B1;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_B2;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_B3;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_B4;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_B5;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_B6;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_BO5;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_BO6;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_BQ;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_B_CY;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_B_XOR;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_C;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_C1;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_C2;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_C3;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_C4;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_C5;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_C6;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_CLK;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_CO5;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_CO6;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_C_CY;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_C_XOR;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_D;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_D1;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_D2;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_D3;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_D4;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_D5;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_D6;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_DO5;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_DO6;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_D_CY;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X6Y158_D_XOR;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_A;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_A1;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_A2;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_A3;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_A4;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_A5;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_A6;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_AO5;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_AO6;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_A_CY;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_A_XOR;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_B;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_B1;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_B2;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_B3;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_B4;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_B5;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_B6;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_BO5;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_BO6;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_B_CY;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_B_XOR;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_C;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_C1;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_C2;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_C3;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_C4;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_C5;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_C6;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_CO5;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_CO6;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_C_CY;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_C_XOR;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_D;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_D1;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_D2;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_D3;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_D4;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_D5;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_D6;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_DO5;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_DO6;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_D_CY;
  wire [0:0] CLBLM_R_X5Y158_SLICE_X7Y158_D_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_AO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_A_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_BO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_BO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_B_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_CLK;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_CO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_CO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_C_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_DO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_DO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X8Y144_D_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_AO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_AO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_A_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_BO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_BO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_B_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_CO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_C_XOR;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D1;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D2;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D3;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D4;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_DO5;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_DO6;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D_CY;
  wire [0:0] CLBLM_R_X7Y144_SLICE_X9Y144_D_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_AO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_AO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_A_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_BO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_BO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_B_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_CLK;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_CO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_CO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_C_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_DO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_DO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X8Y145_D_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_AO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_AO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_A_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_BO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_BO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_B_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_CO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_CO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_C_XOR;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D1;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D2;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D3;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D4;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_DO5;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_DO6;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D_CY;
  wire [0:0] CLBLM_R_X7Y145_SLICE_X9Y145_D_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_AO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_AO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_A_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_BMUX;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_BO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_BO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_B_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_CLK;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_CO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_C_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_DMUX;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_DO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_DO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X8Y146_D_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_AO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_AO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_AQ;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_A_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_BMUX;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_BO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_BO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_B_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_CLK;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_CO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_CO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_C_XOR;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D1;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D2;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D3;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D4;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_DO5;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_DO6;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D_CY;
  wire [0:0] CLBLM_R_X7Y146_SLICE_X9Y146_D_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_AO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_AO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_AQ;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_A_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_BMUX;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_BO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_B_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_CLK;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_CO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_CO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_C_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_DMUX;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_DO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_DO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X8Y147_D_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A5Q;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_AMUX;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_AO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_AO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_A_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_BO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_BO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_BQ;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_B_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_CLK;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_CO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_CO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_CQ;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_C_XOR;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D1;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D2;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D3;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D4;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_DMUX;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_DO5;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_DO6;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D_CY;
  wire [0:0] CLBLM_R_X7Y147_SLICE_X9Y147_D_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A5Q;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_AMUX;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_AO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_AO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_AQ;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_AX;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_A_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_BO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_BO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_BQ;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_B_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_CLK;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_CO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_CO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_CQ;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_C_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_DMUX;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_DO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_DO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X8Y148_D_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_AO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_AO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_AQ;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_A_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_BO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_BO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_BQ;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_B_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_CLK;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_CMUX;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_CO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_CO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_C_XOR;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D1;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D2;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D3;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D4;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_DO5;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_DO6;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D_CY;
  wire [0:0] CLBLM_R_X7Y148_SLICE_X9Y148_D_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_AO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_AO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_A_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_BO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_BO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_BQ;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_B_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_CLK;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_CO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_CO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_CQ;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_C_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_DMUX;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_DO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_DO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X8Y149_D_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_AO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_AO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_A_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_BO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_BO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_BQ;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_B_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C5Q;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_CLK;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_CMUX;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_CO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_CO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_CQ;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_C_XOR;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D1;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D2;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D3;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D4;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_DMUX;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_DO5;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_DO6;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D_CY;
  wire [0:0] CLBLM_R_X7Y149_SLICE_X9Y149_D_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_AO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_AO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_A_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_BO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_BO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_BQ;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_B_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_CLK;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_CMUX;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_CO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_CO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_C_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_DO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_DO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X8Y150_D_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_AMUX;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_AO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_AO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_A_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_BO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_BO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_B_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_CO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_CO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_C_XOR;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D1;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D2;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D3;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D4;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_DO5;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_DO6;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D_CY;
  wire [0:0] CLBLM_R_X7Y150_SLICE_X9Y150_D_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_AO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_AO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_A_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_BO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_BO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_BQ;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_B_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_CLK;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_CO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_CO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_CQ;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_C_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_DO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_DO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_DQ;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X8Y151_D_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_AO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_AO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_AQ;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_A_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_BO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_BO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_BQ;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_B_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C5Q;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_CLK;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_CMUX;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_CO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_CO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_CQ;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_C_XOR;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D1;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D2;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D3;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D4;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_DMUX;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_DO5;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_DO6;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D_CY;
  wire [0:0] CLBLM_R_X7Y151_SLICE_X9Y151_D_XOR;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A1;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A2;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A3;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A4;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A5Q;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_AMUX;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_AO5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_AO6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_AQ;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_AX;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A_CY;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_A_XOR;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B1;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B2;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B3;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B4;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_BMUX;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_BO5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_BO6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B_CY;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_B_XOR;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C1;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C2;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C3;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C4;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_CLK;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_CO5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_CO6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C_CY;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_C_XOR;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D1;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D2;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D3;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D4;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_DO5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_DO6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D_CY;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X8Y152_D_XOR;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A1;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A2;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A3;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A4;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_AO5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_AO6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_AQ;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A_CY;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_A_XOR;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B1;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B2;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B3;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B4;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_BO5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_BO6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_BQ;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B_CY;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_B_XOR;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C1;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C2;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C3;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C4;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_CLK;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_CMUX;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_CO5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_CO6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C_CY;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_C_XOR;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D1;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D2;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D3;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D4;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_DO5;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_DO6;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D_CY;
  wire [0:0] CLBLM_R_X7Y152_SLICE_X9Y152_D_XOR;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A1;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A2;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A3;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A4;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_AMUX;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_AO5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_AO6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_AQ;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A_CY;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_A_XOR;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B1;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B2;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B3;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B4;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_BO5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_BO6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_BQ;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B_CY;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_B_XOR;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C1;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C2;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C3;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C4;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_CLK;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_CO5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_CO6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_CQ;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C_CY;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_C_XOR;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D1;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D2;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D3;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D4;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_DO5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_DO6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D_CY;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X8Y153_D_XOR;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A1;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A2;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A3;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A4;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_AO5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_AO6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_AQ;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A_CY;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_A_XOR;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B1;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B2;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B3;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B4;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_BO5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_BO6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_BQ;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B_CY;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_B_XOR;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C1;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C2;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C3;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C4;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_CLK;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_CMUX;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_CO5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_CO6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C_CY;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_C_XOR;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D1;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D2;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D3;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D4;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_DO5;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_DO6;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D_CY;
  wire [0:0] CLBLM_R_X7Y153_SLICE_X9Y153_D_XOR;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A1;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A2;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A3;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A4;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_AMUX;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_AO5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_AO6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_AQ;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A_CY;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_A_XOR;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B1;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B2;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B3;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B4;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_BO5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_BO6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B_CY;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_B_XOR;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C1;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C2;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C3;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C4;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_CLK;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_CO5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_CO6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_CQ;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C_CY;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_C_XOR;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D1;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D2;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D3;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D4;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_DO5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_DO6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D_CY;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X8Y154_D_XOR;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A1;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A2;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A3;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A4;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_AO5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_AO6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_AQ;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A_CY;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_A_XOR;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B1;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B2;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B3;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B4;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_BO5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_BO6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_BQ;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B_CY;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_B_XOR;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C1;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C2;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C3;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C4;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_CLK;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_CO5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_CO6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_CQ;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C_CY;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_C_XOR;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D1;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D2;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D3;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D4;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_DO5;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_DO6;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D_CY;
  wire [0:0] CLBLM_R_X7Y154_SLICE_X9Y154_D_XOR;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A1;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A2;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A3;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A4;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A5Q;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_AMUX;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_AO5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_AO6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_AQ;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A_CY;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_A_XOR;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B1;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B2;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B3;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B4;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_BMUX;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_BO5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_BO6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B_CY;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_B_XOR;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C1;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C2;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C3;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C4;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_CLK;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_CO5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_CO6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C_CY;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_C_XOR;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D1;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D2;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D3;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D4;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_DO5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_DO6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D_CY;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X8Y155_D_XOR;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A1;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A2;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A3;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A4;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A5Q;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_AMUX;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_AO5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_AO6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_AQ;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_AX;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A_CY;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_A_XOR;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B1;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B2;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B3;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B4;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_BO5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_BO6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_BQ;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B_CY;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_B_XOR;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C1;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C2;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C3;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C4;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_CLK;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_CMUX;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_CO5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_CO6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C_CY;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_C_XOR;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D1;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D2;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D3;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D4;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_DMUX;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_DO5;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_DO6;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D_CY;
  wire [0:0] CLBLM_R_X7Y155_SLICE_X9Y155_D_XOR;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_A;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_A1;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_A2;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_A3;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_A4;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_A5;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_A6;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_AO5;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_AO6;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_AQ;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_A_CY;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_A_XOR;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_B;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_B1;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_B2;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_B3;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_B4;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_B5;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_B6;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_BO5;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_BO6;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_BQ;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_B_CY;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_B_XOR;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_C;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_C1;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_C2;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_C3;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_C4;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_C5;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_C6;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_CLK;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_CO5;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_CO6;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_CQ;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_C_CY;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_C_XOR;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_D;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_D1;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_D2;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_D3;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_D4;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_D5;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_D6;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_DO5;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_DO6;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_DQ;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_D_CY;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X8Y156_D_XOR;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_A;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_A1;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_A2;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_A3;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_A4;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_A5;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_A6;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_AO5;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_AO6;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_AQ;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_A_CY;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_A_XOR;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_B;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_B1;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_B2;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_B3;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_B4;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_B5;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_B6;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_BO5;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_BO6;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_BQ;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_B_CY;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_B_XOR;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_C;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_C1;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_C2;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_C3;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_C4;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_C5;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_C6;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_CLK;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_CO5;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_CO6;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_CQ;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_C_CY;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_C_XOR;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_D;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_D1;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_D2;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_D3;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_D4;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_D5;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_D6;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_DO5;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_DO6;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_D_CY;
  wire [0:0] CLBLM_R_X7Y156_SLICE_X9Y156_D_XOR;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_A;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_A1;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_A2;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_A3;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_A4;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_A5;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_A6;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_AO5;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_AO6;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_AQ;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_A_CY;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_A_XOR;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_B;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_B1;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_B2;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_B3;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_B4;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_B5;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_B6;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_BO5;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_BO6;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_BQ;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_B_CY;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_B_XOR;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_C;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_C1;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_C2;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_C3;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_C4;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_C5;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_C6;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_CLK;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_CO5;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_CO6;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_CQ;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_C_CY;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_C_XOR;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_D;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_D1;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_D2;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_D3;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_D4;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_D5;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_D6;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_DO5;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_DO6;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_DQ;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_D_CY;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X8Y157_D_XOR;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_A;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_A1;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_A2;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_A3;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_A4;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_A5;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_A6;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_AO5;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_AO6;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_AQ;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_A_CY;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_A_XOR;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_B;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_B1;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_B2;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_B3;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_B4;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_B5;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_B6;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_BO5;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_BO6;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_BQ;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_B_CY;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_B_XOR;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_C;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_C1;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_C2;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_C3;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_C4;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_C5;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_C6;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_CLK;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_CO5;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_CO6;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_CQ;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_C_CY;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_C_XOR;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_D;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_D1;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_D2;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_D3;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_D4;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_D5;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_D6;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_DO5;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_DO6;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_DQ;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_D_CY;
  wire [0:0] CLBLM_R_X7Y157_SLICE_X9Y157_D_XOR;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_A;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_A1;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_A2;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_A3;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_A4;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_A5;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_A6;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_AO5;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_AO6;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_AQ;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_A_CY;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_A_XOR;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_B;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_B1;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_B2;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_B3;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_B4;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_B5;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_B6;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_BO5;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_BO6;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_BQ;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_B_CY;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_B_XOR;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_C;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_C1;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_C2;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_C3;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_C4;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_C5;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_C6;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_CLK;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_CMUX;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_CO5;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_CO6;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_C_CY;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_C_XOR;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_D;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_D1;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_D2;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_D3;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_D4;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_D5;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_D6;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_DO5;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_DO6;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_D_CY;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X8Y158_D_XOR;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_A;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_A1;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_A2;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_A3;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_A4;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_A5;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_A6;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_AO5;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_AO6;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_AQ;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_A_CY;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_A_XOR;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_B;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_B1;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_B2;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_B3;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_B4;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_B5;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_B6;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_BO5;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_BO6;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_B_CY;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_B_XOR;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_C;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_C1;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_C2;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_C3;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_C4;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_C5;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_C6;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_CLK;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_CO5;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_CO6;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_C_CY;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_C_XOR;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_D;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_D1;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_D2;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_D3;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_D4;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_D5;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_D6;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_DO5;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_DO6;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_D_CY;
  wire [0:0] CLBLM_R_X7Y158_SLICE_X9Y158_D_XOR;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_A;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_A1;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_A2;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_A3;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_A4;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_A5;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_A6;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_AO5;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_AO6;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_AQ;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_A_CY;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_A_XOR;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_B;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_B1;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_B2;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_B3;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_B4;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_B5;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_B6;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_BMUX;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_BO5;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_BO6;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_B_CY;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_B_XOR;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_C;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_C1;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_C2;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_C3;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_C4;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_C5;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_C6;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_CLK;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_CO5;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_CO6;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_C_CY;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_C_XOR;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_D;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_D1;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_D2;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_D3;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_D4;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_D5;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_D6;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_DO5;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_DO6;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_D_CY;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X8Y159_D_XOR;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_A;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_A1;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_A2;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_A3;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_A4;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_A5;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_A6;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_AO5;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_AO6;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_A_CY;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_A_XOR;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_B;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_B1;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_B2;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_B3;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_B4;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_B5;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_B6;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_BMUX;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_BO5;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_BO6;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_B_CY;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_B_XOR;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_C;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_C1;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_C2;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_C3;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_C4;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_C5;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_C6;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_CO5;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_CO6;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_C_CY;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_C_XOR;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_D;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_D1;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_D2;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_D3;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_D4;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_D5;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_D6;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_DO5;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_DO6;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_D_CY;
  wire [0:0] CLBLM_R_X7Y159_SLICE_X9Y159_D_XOR;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  wire [0:0] CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_CE;
  wire [0:0] CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_I;
  wire [0:0] CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_O;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_O;
  wire [0:0] LIOB33_SING_X0Y150_IOB_X0Y150_O;
  wire [0:0] LIOB33_SING_X0Y199_IOB_X0Y199_O;
  wire [0:0] LIOB33_SING_X0Y50_IOB_X0Y50_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_O;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_O;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_O;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_O;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_O;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_O;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_O;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_O;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y151_O;
  wire [0:0] LIOB33_X0Y151_IOB_X0Y152_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y153_O;
  wire [0:0] LIOB33_X0Y153_IOB_X0Y154_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y155_O;
  wire [0:0] LIOB33_X0Y155_IOB_X0Y156_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y157_O;
  wire [0:0] LIOB33_X0Y157_IOB_X0Y158_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y159_O;
  wire [0:0] LIOB33_X0Y159_IOB_X0Y160_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y161_O;
  wire [0:0] LIOB33_X0Y161_IOB_X0Y162_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y163_O;
  wire [0:0] LIOB33_X0Y163_IOB_X0Y164_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y165_O;
  wire [0:0] LIOB33_X0Y165_IOB_X0Y166_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y167_O;
  wire [0:0] LIOB33_X0Y167_IOB_X0Y168_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y169_O;
  wire [0:0] LIOB33_X0Y169_IOB_X0Y170_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y171_O;
  wire [0:0] LIOB33_X0Y171_IOB_X0Y172_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y173_O;
  wire [0:0] LIOB33_X0Y173_IOB_X0Y174_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y175_O;
  wire [0:0] LIOB33_X0Y175_IOB_X0Y176_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y177_O;
  wire [0:0] LIOB33_X0Y177_IOB_X0Y178_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y179_O;
  wire [0:0] LIOB33_X0Y179_IOB_X0Y180_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y181_O;
  wire [0:0] LIOB33_X0Y181_IOB_X0Y182_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y183_O;
  wire [0:0] LIOB33_X0Y183_IOB_X0Y184_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y185_O;
  wire [0:0] LIOB33_X0Y185_IOB_X0Y186_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y187_O;
  wire [0:0] LIOB33_X0Y187_IOB_X0Y188_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y189_O;
  wire [0:0] LIOB33_X0Y189_IOB_X0Y190_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y191_O;
  wire [0:0] LIOB33_X0Y191_IOB_X0Y192_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y193_O;
  wire [0:0] LIOB33_X0Y193_IOB_X0Y194_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y195_O;
  wire [0:0] LIOB33_X0Y195_IOB_X0Y196_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y197_O;
  wire [0:0] LIOB33_X0Y197_IOB_X0Y198_O;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y51_I;
  wire [0:0] LIOB33_X0Y51_IOB_X0Y52_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y53_I;
  wire [0:0] LIOB33_X0Y53_IOB_X0Y54_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y55_I;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y56_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y57_I;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y58_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y59_I;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y60_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y61_I;
  wire [0:0] LIOB33_X0Y61_IOB_X0Y62_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y63_I;
  wire [0:0] LIOB33_X0Y63_IOB_X0Y64_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y65_I;
  wire [0:0] LIOB33_X0Y65_IOB_X0Y66_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y67_I;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y68_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y69_I;
  wire [0:0] LIOB33_X0Y69_IOB_X0Y70_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y71_I;
  wire [0:0] LIOB33_X0Y71_IOB_X0Y72_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y73_I;
  wire [0:0] LIOB33_X0Y73_IOB_X0Y74_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y75_I;
  wire [0:0] LIOB33_X0Y75_IOB_X0Y76_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y77_I;
  wire [0:0] LIOB33_X0Y77_IOB_X0Y78_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y79_I;
  wire [0:0] LIOB33_X0Y79_IOB_X0Y80_O;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1;
  wire [0:0] LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1;
  wire [0:0] LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1;
  wire [0:0] LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_D;
  wire [0:0] LIOI3_SING_X0Y50_ILOGIC_X0Y50_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_O;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y101_TQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_D1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_OQ;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_T1;
  wire [0:0] LIOI3_X0Y101_OLOGIC_X0Y102_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y103_TQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_D1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_OQ;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_T1;
  wire [0:0] LIOI3_X0Y103_OLOGIC_X0Y104_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y105_TQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_D1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_OQ;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_T1;
  wire [0:0] LIOI3_X0Y105_OLOGIC_X0Y106_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y109_TQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_D1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_OQ;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_T1;
  wire [0:0] LIOI3_X0Y109_OLOGIC_X0Y110_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_TQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y112_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y115_TQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_D1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_OQ;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_T1;
  wire [0:0] LIOI3_X0Y115_OLOGIC_X0Y116_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y117_TQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y151_TQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_D1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_OQ;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_T1;
  wire [0:0] LIOI3_X0Y151_OLOGIC_X0Y152_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y153_TQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_D1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_OQ;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_T1;
  wire [0:0] LIOI3_X0Y153_OLOGIC_X0Y154_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y155_TQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_D1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_OQ;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_T1;
  wire [0:0] LIOI3_X0Y155_OLOGIC_X0Y156_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y159_TQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_D1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_OQ;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_T1;
  wire [0:0] LIOI3_X0Y159_OLOGIC_X0Y160_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y161_TQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_D1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_OQ;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_T1;
  wire [0:0] LIOI3_X0Y161_OLOGIC_X0Y162_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y165_TQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_D1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_OQ;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_T1;
  wire [0:0] LIOI3_X0Y165_OLOGIC_X0Y166_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y167_TQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_D1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_OQ;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_T1;
  wire [0:0] LIOI3_X0Y167_OLOGIC_X0Y168_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y171_TQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_D1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_OQ;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_T1;
  wire [0:0] LIOI3_X0Y171_OLOGIC_X0Y172_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y173_TQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_D1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_OQ;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_T1;
  wire [0:0] LIOI3_X0Y173_OLOGIC_X0Y174_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y175_TQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_D1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_OQ;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_T1;
  wire [0:0] LIOI3_X0Y175_OLOGIC_X0Y176_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y177_TQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_D1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_OQ;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_T1;
  wire [0:0] LIOI3_X0Y177_OLOGIC_X0Y178_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y179_TQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_D1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_OQ;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_T1;
  wire [0:0] LIOI3_X0Y179_OLOGIC_X0Y180_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y183_TQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_D1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_OQ;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_T1;
  wire [0:0] LIOI3_X0Y183_OLOGIC_X0Y184_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y185_TQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_D1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_OQ;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_T1;
  wire [0:0] LIOI3_X0Y185_OLOGIC_X0Y186_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y189_TQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_D1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_OQ;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_T1;
  wire [0:0] LIOI3_X0Y189_OLOGIC_X0Y190_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y191_TQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_D1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_OQ;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_T1;
  wire [0:0] LIOI3_X0Y191_OLOGIC_X0Y192_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y195_TQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_D1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_OQ;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_T1;
  wire [0:0] LIOI3_X0Y195_OLOGIC_X0Y196_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y197_TQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_D1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_OQ;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_T1;
  wire [0:0] LIOI3_X0Y197_OLOGIC_X0Y198_TQ;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y51_O;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_D;
  wire [0:0] LIOI3_X0Y51_ILOGIC_X0Y52_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y53_O;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_D;
  wire [0:0] LIOI3_X0Y53_ILOGIC_X0Y54_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y55_O;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_D;
  wire [0:0] LIOI3_X0Y55_ILOGIC_X0Y56_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y59_O;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_D;
  wire [0:0] LIOI3_X0Y59_ILOGIC_X0Y60_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y61_O;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_D;
  wire [0:0] LIOI3_X0Y61_ILOGIC_X0Y62_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y65_O;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_D;
  wire [0:0] LIOI3_X0Y65_ILOGIC_X0Y66_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y67_O;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_D;
  wire [0:0] LIOI3_X0Y67_ILOGIC_X0Y68_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y71_O;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_D;
  wire [0:0] LIOI3_X0Y71_ILOGIC_X0Y72_O;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y73_D;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y73_O;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_D;
  wire [0:0] LIOI3_X0Y73_ILOGIC_X0Y74_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y75_O;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_D;
  wire [0:0] LIOI3_X0Y75_ILOGIC_X0Y76_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y77_O;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_D;
  wire [0:0] LIOI3_X0Y77_ILOGIC_X0Y78_O;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_D;
  wire [0:0] LIOI3_X0Y79_ILOGIC_X0Y79_O;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_D1;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_OQ;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_T1;
  wire [0:0] LIOI3_X0Y79_OLOGIC_X0Y80_TQ;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_I;
  wire [0:0] RIOB33_SING_X105Y149_IOB_X1Y149_I;
  wire [0:0] RIOB33_SING_X105Y150_IOB_X1Y150_O;
  wire [0:0] RIOB33_SING_X105Y199_IOB_X1Y199_O;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y114_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y115_I;
  wire [0:0] RIOB33_X105Y115_IOB_X1Y116_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y117_I;
  wire [0:0] RIOB33_X105Y117_IOB_X1Y118_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y119_I;
  wire [0:0] RIOB33_X105Y119_IOB_X1Y120_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y121_I;
  wire [0:0] RIOB33_X105Y121_IOB_X1Y122_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y123_I;
  wire [0:0] RIOB33_X105Y123_IOB_X1Y124_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y125_I;
  wire [0:0] RIOB33_X105Y125_IOB_X1Y126_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y127_I;
  wire [0:0] RIOB33_X105Y127_IOB_X1Y128_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y129_I;
  wire [0:0] RIOB33_X105Y129_IOB_X1Y130_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y131_I;
  wire [0:0] RIOB33_X105Y131_IOB_X1Y132_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y133_I;
  wire [0:0] RIOB33_X105Y133_IOB_X1Y134_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y135_I;
  wire [0:0] RIOB33_X105Y135_IOB_X1Y136_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y137_I;
  wire [0:0] RIOB33_X105Y137_IOB_X1Y138_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y139_I;
  wire [0:0] RIOB33_X105Y139_IOB_X1Y140_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y141_I;
  wire [0:0] RIOB33_X105Y141_IOB_X1Y142_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y143_I;
  wire [0:0] RIOB33_X105Y143_IOB_X1Y144_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y145_I;
  wire [0:0] RIOB33_X105Y145_IOB_X1Y146_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y147_I;
  wire [0:0] RIOB33_X105Y147_IOB_X1Y148_I;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y151_O;
  wire [0:0] RIOB33_X105Y151_IOB_X1Y152_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y153_O;
  wire [0:0] RIOB33_X105Y153_IOB_X1Y154_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y155_O;
  wire [0:0] RIOB33_X105Y155_IOB_X1Y156_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y157_O;
  wire [0:0] RIOB33_X105Y157_IOB_X1Y158_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y159_O;
  wire [0:0] RIOB33_X105Y159_IOB_X1Y160_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y161_O;
  wire [0:0] RIOB33_X105Y161_IOB_X1Y162_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y163_O;
  wire [0:0] RIOB33_X105Y163_IOB_X1Y164_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y165_O;
  wire [0:0] RIOB33_X105Y165_IOB_X1Y166_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y167_O;
  wire [0:0] RIOB33_X105Y167_IOB_X1Y168_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y169_O;
  wire [0:0] RIOB33_X105Y169_IOB_X1Y170_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y171_O;
  wire [0:0] RIOB33_X105Y171_IOB_X1Y172_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y173_O;
  wire [0:0] RIOB33_X105Y173_IOB_X1Y174_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y175_O;
  wire [0:0] RIOB33_X105Y175_IOB_X1Y176_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y177_O;
  wire [0:0] RIOB33_X105Y177_IOB_X1Y178_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y179_O;
  wire [0:0] RIOB33_X105Y179_IOB_X1Y180_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y181_O;
  wire [0:0] RIOB33_X105Y181_IOB_X1Y182_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y183_O;
  wire [0:0] RIOB33_X105Y183_IOB_X1Y184_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y185_O;
  wire [0:0] RIOB33_X105Y185_IOB_X1Y186_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y187_O;
  wire [0:0] RIOB33_X105Y187_IOB_X1Y188_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y189_O;
  wire [0:0] RIOB33_X105Y189_IOB_X1Y190_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y191_O;
  wire [0:0] RIOB33_X105Y191_IOB_X1Y192_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y193_O;
  wire [0:0] RIOB33_X105Y193_IOB_X1Y194_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y195_O;
  wire [0:0] RIOB33_X105Y195_IOB_X1Y196_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y197_O;
  wire [0:0] RIOB33_X105Y197_IOB_X1Y198_O;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_D;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_O;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_D;
  wire [0:0] RIOI3_SING_X105Y149_ILOGIC_X1Y149_O;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1;
  wire [0:0] RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1;
  wire [0:0] RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1;
  wire [0:0] RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1;
  wire [0:0] RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y115_O;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_D;
  wire [0:0] RIOI3_X105Y115_ILOGIC_X1Y116_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y117_O;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_D;
  wire [0:0] RIOI3_X105Y117_ILOGIC_X1Y118_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y121_O;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_D;
  wire [0:0] RIOI3_X105Y121_ILOGIC_X1Y122_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y123_O;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_D;
  wire [0:0] RIOI3_X105Y123_ILOGIC_X1Y124_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y125_O;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_D;
  wire [0:0] RIOI3_X105Y125_ILOGIC_X1Y126_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y127_O;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_D;
  wire [0:0] RIOI3_X105Y127_ILOGIC_X1Y128_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y129_O;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_D;
  wire [0:0] RIOI3_X105Y129_ILOGIC_X1Y130_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y133_O;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_D;
  wire [0:0] RIOI3_X105Y133_ILOGIC_X1Y134_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y135_O;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_D;
  wire [0:0] RIOI3_X105Y135_ILOGIC_X1Y136_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y139_O;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_D;
  wire [0:0] RIOI3_X105Y139_ILOGIC_X1Y140_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y141_O;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_D;
  wire [0:0] RIOI3_X105Y141_ILOGIC_X1Y142_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y145_O;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_D;
  wire [0:0] RIOI3_X105Y145_ILOGIC_X1Y146_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y147_O;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_D;
  wire [0:0] RIOI3_X105Y147_ILOGIC_X1Y148_O;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y151_TQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_D1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_OQ;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_T1;
  wire [0:0] RIOI3_X105Y151_OLOGIC_X1Y152_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y153_TQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_D1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_OQ;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_T1;
  wire [0:0] RIOI3_X105Y153_OLOGIC_X1Y154_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y155_TQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_D1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_OQ;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_T1;
  wire [0:0] RIOI3_X105Y155_OLOGIC_X1Y156_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y159_TQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_D1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_OQ;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_T1;
  wire [0:0] RIOI3_X105Y159_OLOGIC_X1Y160_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y161_TQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_D1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_OQ;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_T1;
  wire [0:0] RIOI3_X105Y161_OLOGIC_X1Y162_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y165_TQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_D1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_OQ;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_T1;
  wire [0:0] RIOI3_X105Y165_OLOGIC_X1Y166_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y167_TQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_D1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_OQ;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_T1;
  wire [0:0] RIOI3_X105Y167_OLOGIC_X1Y168_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y171_TQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_D1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_OQ;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_T1;
  wire [0:0] RIOI3_X105Y171_OLOGIC_X1Y172_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y173_TQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_D1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_OQ;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_T1;
  wire [0:0] RIOI3_X105Y173_OLOGIC_X1Y174_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y175_TQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_D1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_OQ;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_T1;
  wire [0:0] RIOI3_X105Y175_OLOGIC_X1Y176_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y177_TQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_D1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_OQ;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_T1;
  wire [0:0] RIOI3_X105Y177_OLOGIC_X1Y178_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y179_TQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_D1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_OQ;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_T1;
  wire [0:0] RIOI3_X105Y179_OLOGIC_X1Y180_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y183_TQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_D1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_OQ;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_T1;
  wire [0:0] RIOI3_X105Y183_OLOGIC_X1Y184_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y185_TQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_D1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_OQ;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_T1;
  wire [0:0] RIOI3_X105Y185_OLOGIC_X1Y186_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y189_TQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_D1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_OQ;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_T1;
  wire [0:0] RIOI3_X105Y189_OLOGIC_X1Y190_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y191_TQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_D1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_OQ;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_T1;
  wire [0:0] RIOI3_X105Y191_OLOGIC_X1Y192_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y195_TQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_D1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_OQ;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_T1;
  wire [0:0] RIOI3_X105Y195_OLOGIC_X1Y196_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y197_TQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_D1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_OQ;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_T1;
  wire [0:0] RIOI3_X105Y197_OLOGIC_X1Y198_TQ;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y139_SLICE_X0Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y139_SLICE_X0Y139_DO5),
.O6(CLBLL_L_X2Y139_SLICE_X0Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y139_SLICE_X0Y139_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y139_SLICE_X0Y139_CO5),
.O6(CLBLL_L_X2Y139_SLICE_X0Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff5fffffffdfffd)
  ) CLBLL_L_X2Y139_SLICE_X0Y139_BLUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(CLBLL_L_X4Y154_SLICE_X5Y154_BO6),
.I2(RIOB33_X105Y129_IOB_X1Y129_I),
.I3(RIOB33_X105Y127_IOB_X1Y128_I),
.I4(CLBLL_L_X4Y153_SLICE_X4Y153_AO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y139_SLICE_X0Y139_BO5),
.O6(CLBLL_L_X2Y139_SLICE_X0Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffdfffdffffffdd)
  ) CLBLL_L_X2Y139_SLICE_X0Y139_ALUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(CLBLM_R_X3Y156_SLICE_X2Y156_DO6),
.I3(RIOB33_X105Y127_IOB_X1Y128_I),
.I4(CLBLL_L_X4Y154_SLICE_X4Y154_BO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y139_SLICE_X0Y139_AO5),
.O6(CLBLL_L_X2Y139_SLICE_X0Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y139_SLICE_X1Y139_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y139_SLICE_X1Y139_DO5),
.O6(CLBLL_L_X2Y139_SLICE_X1Y139_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y139_SLICE_X1Y139_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y139_SLICE_X1Y139_CO5),
.O6(CLBLL_L_X2Y139_SLICE_X1Y139_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y139_SLICE_X1Y139_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y139_SLICE_X1Y139_BO5),
.O6(CLBLL_L_X2Y139_SLICE_X1Y139_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y139_SLICE_X1Y139_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y139_SLICE_X1Y139_AO5),
.O6(CLBLL_L_X2Y139_SLICE_X1Y139_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y140_SLICE_X0Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y140_SLICE_X0Y140_DO5),
.O6(CLBLL_L_X2Y140_SLICE_X0Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y140_SLICE_X0Y140_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y140_SLICE_X0Y140_CO5),
.O6(CLBLL_L_X2Y140_SLICE_X0Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffafffffffcff)
  ) CLBLL_L_X2Y140_SLICE_X0Y140_BLUT (
.I0(CLBLL_L_X4Y154_SLICE_X5Y154_CO6),
.I1(CLBLL_L_X4Y153_SLICE_X4Y153_BO6),
.I2(RIOB33_X105Y127_IOB_X1Y128_I),
.I3(RIOB33_X105Y137_IOB_X1Y137_I),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y140_SLICE_X0Y140_BO5),
.O6(CLBLL_L_X2Y140_SLICE_X0Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffefefffffffcf)
  ) CLBLL_L_X2Y140_SLICE_X0Y140_ALUT (
.I0(CLBLM_R_X5Y155_SLICE_X6Y155_DO6),
.I1(RIOB33_X105Y127_IOB_X1Y128_I),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(CLBLM_R_X3Y155_SLICE_X2Y155_BO6),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y140_SLICE_X0Y140_AO5),
.O6(CLBLL_L_X2Y140_SLICE_X0Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y140_SLICE_X1Y140_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y140_SLICE_X1Y140_DO5),
.O6(CLBLL_L_X2Y140_SLICE_X1Y140_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y140_SLICE_X1Y140_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y140_SLICE_X1Y140_CO5),
.O6(CLBLL_L_X2Y140_SLICE_X1Y140_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y140_SLICE_X1Y140_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y140_SLICE_X1Y140_BO5),
.O6(CLBLL_L_X2Y140_SLICE_X1Y140_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y140_SLICE_X1Y140_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y140_SLICE_X1Y140_AO5),
.O6(CLBLL_L_X2Y140_SLICE_X1Y140_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y153_SLICE_X0Y153_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y153_SLICE_X0Y153_DO5),
.O6(CLBLL_L_X2Y153_SLICE_X0Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y153_SLICE_X0Y153_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y153_SLICE_X0Y153_CO5),
.O6(CLBLL_L_X2Y153_SLICE_X0Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y153_SLICE_X0Y153_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y153_SLICE_X0Y153_BO5),
.O6(CLBLL_L_X2Y153_SLICE_X0Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000200000)
  ) CLBLL_L_X2Y153_SLICE_X0Y153_ALUT (
.I0(LIOB33_X0Y71_IOB_X0Y71_I),
.I1(CLBLL_L_X4Y157_SLICE_X4Y157_CO6),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(RIOB33_X105Y133_IOB_X1Y134_I),
.O5(CLBLL_L_X2Y153_SLICE_X0Y153_AO5),
.O6(CLBLL_L_X2Y153_SLICE_X0Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fdf0fcf55dd00cc)
  ) CLBLL_L_X2Y153_SLICE_X1Y153_DLUT (
.I0(CLBLM_R_X3Y153_SLICE_X2Y153_AO6),
.I1(LIOB33_X0Y53_IOB_X0Y54_I),
.I2(CLBLM_R_X3Y151_SLICE_X2Y151_CO5),
.I3(CLBLL_L_X2Y154_SLICE_X1Y154_AO5),
.I4(CLBLL_L_X4Y155_SLICE_X4Y155_AQ),
.I5(CLBLM_R_X5Y156_SLICE_X7Y156_AQ),
.O5(CLBLL_L_X2Y153_SLICE_X1Y153_DO5),
.O6(CLBLL_L_X2Y153_SLICE_X1Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0200010102000000)
  ) CLBLL_L_X2Y153_SLICE_X1Y153_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLM_R_X3Y152_SLICE_X2Y152_AO5),
.I2(CLBLL_L_X4Y157_SLICE_X4Y157_CO6),
.I3(LIOB33_X0Y53_IOB_X0Y54_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_R_X5Y156_SLICE_X7Y156_AQ),
.O5(CLBLL_L_X2Y153_SLICE_X1Y153_CO5),
.O6(CLBLL_L_X2Y153_SLICE_X1Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f0ccfcaafaeefe)
  ) CLBLL_L_X2Y153_SLICE_X1Y153_BLUT (
.I0(LIOB33_X0Y55_IOB_X0Y55_I),
.I1(LIOB33_X0Y71_IOB_X0Y71_I),
.I2(RIOB33_X105Y115_IOB_X1Y115_I),
.I3(CLBLM_R_X3Y153_SLICE_X2Y153_CO6),
.I4(CLBLL_L_X2Y153_SLICE_X1Y153_AO6),
.I5(CLBLL_L_X2Y154_SLICE_X1Y154_AO5),
.O5(CLBLL_L_X2Y153_SLICE_X1Y153_BO5),
.O6(CLBLL_L_X2Y153_SLICE_X1Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffdfffffff7f)
  ) CLBLL_L_X2Y153_SLICE_X1Y153_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLL_L_X4Y157_SLICE_X4Y157_CO6),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y153_SLICE_X1Y153_AO5),
.O6(CLBLL_L_X2Y153_SLICE_X1Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y154_SLICE_X0Y154_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y154_SLICE_X0Y154_DO5),
.O6(CLBLL_L_X2Y154_SLICE_X0Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y154_SLICE_X0Y154_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y154_SLICE_X0Y154_CO5),
.O6(CLBLL_L_X2Y154_SLICE_X0Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y154_SLICE_X0Y154_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y154_SLICE_X0Y154_BO5),
.O6(CLBLL_L_X2Y154_SLICE_X0Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y154_SLICE_X0Y154_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y154_SLICE_X0Y154_AO5),
.O6(CLBLL_L_X2Y154_SLICE_X0Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y154_SLICE_X1Y154_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y154_SLICE_X1Y154_DO5),
.O6(CLBLL_L_X2Y154_SLICE_X1Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y154_SLICE_X1Y154_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y154_SLICE_X1Y154_CO5),
.O6(CLBLL_L_X2Y154_SLICE_X1Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y154_SLICE_X1Y154_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y154_SLICE_X1Y154_BO5),
.O6(CLBLL_L_X2Y154_SLICE_X1Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h15000100efffffff)
  ) CLBLL_L_X2Y154_SLICE_X1Y154_ALUT (
.I0(CLBLL_L_X4Y157_SLICE_X4Y157_CO6),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y154_SLICE_X1Y154_AO5),
.O6(CLBLL_L_X2Y154_SLICE_X1Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y155_SLICE_X0Y155_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y155_SLICE_X0Y155_DO5),
.O6(CLBLL_L_X2Y155_SLICE_X0Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y155_SLICE_X0Y155_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y155_SLICE_X0Y155_CO5),
.O6(CLBLL_L_X2Y155_SLICE_X0Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y155_SLICE_X0Y155_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y155_SLICE_X0Y155_BO5),
.O6(CLBLL_L_X2Y155_SLICE_X0Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y155_SLICE_X0Y155_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y155_SLICE_X0Y155_AO5),
.O6(CLBLL_L_X2Y155_SLICE_X0Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hedcceccccccccccc)
  ) CLBLL_L_X2Y155_SLICE_X1Y155_DLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(CLBLM_R_X3Y155_SLICE_X2Y155_DO6),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLM_R_X3Y158_SLICE_X2Y158_AO6),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLL_L_X2Y155_SLICE_X1Y155_DO5),
.O6(CLBLL_L_X2Y155_SLICE_X1Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff7f7ffbfbffff)
  ) CLBLL_L_X2Y155_SLICE_X1Y155_CLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(1'b1),
.I4(RIOB33_X105Y133_IOB_X1Y134_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y155_SLICE_X1Y155_CO5),
.O6(CLBLL_L_X2Y155_SLICE_X1Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha8000020dfffffff)
  ) CLBLL_L_X2Y155_SLICE_X1Y155_BLUT (
.I0(CLBLM_R_X3Y158_SLICE_X2Y158_AO6),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y155_SLICE_X1Y155_BO5),
.O6(CLBLL_L_X2Y155_SLICE_X1Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88000000fcffffff)
  ) CLBLL_L_X2Y155_SLICE_X1Y155_ALUT (
.I0(CLBLM_R_X3Y158_SLICE_X2Y158_AO6),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y155_SLICE_X1Y155_AO5),
.O6(CLBLL_L_X2Y155_SLICE_X1Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y146_SLICE_X4Y146_DO5),
.O6(CLBLL_L_X4Y146_SLICE_X4Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y146_SLICE_X4Y146_CO5),
.O6(CLBLL_L_X4Y146_SLICE_X4Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y146_SLICE_X4Y146_BO5),
.O6(CLBLL_L_X4Y146_SLICE_X4Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y146_SLICE_X4Y146_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y146_SLICE_X4Y146_AO5),
.O6(CLBLL_L_X4Y146_SLICE_X4Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y146_SLICE_X5Y146_AO6),
.Q(CLBLL_L_X4Y146_SLICE_X5Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y146_SLICE_X5Y146_DO5),
.O6(CLBLL_L_X4Y146_SLICE_X5Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y146_SLICE_X5Y146_CO5),
.O6(CLBLL_L_X4Y146_SLICE_X5Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y146_SLICE_X5Y146_BO5),
.O6(CLBLL_L_X4Y146_SLICE_X5Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaac000c000)
  ) CLBLL_L_X4Y146_SLICE_X5Y146_ALUT (
.I0(CLBLM_R_X5Y149_SLICE_X7Y149_CQ),
.I1(CLBLM_R_X5Y144_SLICE_X6Y144_CO6),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_BQ),
.I3(CLBLM_R_X5Y144_SLICE_X6Y144_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y146_SLICE_X5Y146_AO5),
.O6(CLBLL_L_X4Y146_SLICE_X5Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y147_SLICE_X4Y147_DO5),
.O6(CLBLL_L_X4Y147_SLICE_X4Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y147_SLICE_X4Y147_CO5),
.O6(CLBLL_L_X4Y147_SLICE_X4Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h50505050d0d0f0f0)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLL_L_X4Y151_SLICE_X4Y151_C5Q),
.I2(CLBLM_L_X8Y147_SLICE_X11Y147_CO6),
.I3(1'b1),
.I4(CLBLM_R_X3Y151_SLICE_X2Y151_AQ),
.I5(CLBLM_R_X5Y149_SLICE_X6Y149_B5Q),
.O5(CLBLL_L_X4Y147_SLICE_X4Y147_BO5),
.O6(CLBLL_L_X4Y147_SLICE_X4Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf222f00022220000)
  ) CLBLL_L_X4Y147_SLICE_X4Y147_ALUT (
.I0(CLBLL_L_X4Y154_SLICE_X5Y154_CO6),
.I1(CLBLL_L_X4Y151_SLICE_X4Y151_C5Q),
.I2(CLBLL_L_X4Y154_SLICE_X5Y154_BO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X3Y151_SLICE_X2Y151_AQ),
.I5(CLBLM_R_X5Y149_SLICE_X6Y149_B5Q),
.O5(CLBLL_L_X4Y147_SLICE_X4Y147_AO5),
.O6(CLBLL_L_X4Y147_SLICE_X4Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X5Y147_AO6),
.Q(CLBLL_L_X4Y147_SLICE_X5Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y147_SLICE_X5Y147_BO6),
.Q(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y147_SLICE_X5Y147_DO5),
.O6(CLBLL_L_X4Y147_SLICE_X5Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y147_SLICE_X5Y147_CO5),
.O6(CLBLL_L_X4Y147_SLICE_X5Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0002020808)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I2(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I3(CLBLM_R_X5Y149_SLICE_X6Y149_B5Q),
.I4(CLBLL_L_X4Y146_SLICE_X5Y146_AO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y147_SLICE_X5Y147_BO5),
.O6(CLBLL_L_X4Y147_SLICE_X5Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbefafafa14505050)
  ) CLBLL_L_X4Y147_SLICE_X5Y147_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I2(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I3(CLBLM_R_X5Y147_SLICE_X6Y147_AQ),
.I4(CLBLL_L_X4Y146_SLICE_X5Y146_AO5),
.I5(CLBLM_L_X10Y148_SLICE_X13Y148_BQ),
.O5(CLBLL_L_X4Y147_SLICE_X5Y147_AO5),
.O6(CLBLL_L_X4Y147_SLICE_X5Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y148_SLICE_X4Y148_AO6),
.Q(CLBLL_L_X4Y148_SLICE_X4Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y148_SLICE_X4Y148_DO5),
.O6(CLBLL_L_X4Y148_SLICE_X4Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f03035fff53f3)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_CLUT (
.I0(CLBLL_L_X4Y150_SLICE_X5Y150_C5Q),
.I1(CLBLM_R_X5Y155_SLICE_X6Y155_DO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLL_L_X4Y154_SLICE_X5Y154_BO6),
.I4(CLBLL_L_X4Y148_SLICE_X4Y148_BO5),
.I5(CLBLL_L_X4Y149_SLICE_X5Y149_DO6),
.O5(CLBLL_L_X4Y148_SLICE_X4Y148_CO5),
.O6(CLBLL_L_X4Y148_SLICE_X4Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdc10cc000f0fffff)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y151_SLICE_X4Y151_BQ),
.I3(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I4(CLBLM_L_X10Y151_SLICE_X12Y151_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y148_SLICE_X4Y148_BO5),
.O6(CLBLL_L_X4Y148_SLICE_X4Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ff33ce02df13)
  ) CLBLL_L_X4Y148_SLICE_X4Y148_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y152_SLICE_X4Y152_AQ),
.I3(CLBLM_R_X11Y148_SLICE_X15Y148_AQ),
.I4(LIOB33_X0Y53_IOB_X0Y53_I),
.I5(CLBLL_L_X4Y151_SLICE_X4Y151_CQ),
.O5(CLBLL_L_X4Y148_SLICE_X4Y148_AO5),
.O6(CLBLL_L_X4Y148_SLICE_X4Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y148_SLICE_X5Y148_AO6),
.Q(CLBLL_L_X4Y148_SLICE_X5Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y148_SLICE_X5Y148_BO6),
.Q(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y148_SLICE_X5Y148_CO6),
.Q(CLBLL_L_X4Y148_SLICE_X5Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y148_SLICE_X5Y148_DO6),
.Q(CLBLL_L_X4Y148_SLICE_X5Y148_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff480048ffc000c0)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_DLUT (
.I0(CLBLM_L_X10Y149_SLICE_X12Y149_BQ),
.I1(CLBLM_L_X10Y149_SLICE_X12Y149_DO5),
.I2(CLBLL_L_X4Y148_SLICE_X5Y148_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y148_SLICE_X5Y148_AQ),
.I5(CLBLM_R_X7Y148_SLICE_X8Y148_A5Q),
.O5(CLBLL_L_X4Y148_SLICE_X5Y148_DO5),
.O6(CLBLL_L_X4Y148_SLICE_X5Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaa00eeccaa00)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_CLUT (
.I0(CLBLM_R_X5Y148_SLICE_X7Y148_BQ),
.I1(CLBLL_L_X4Y148_SLICE_X5Y148_CQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y152_SLICE_X6Y152_CO6),
.I5(CLBLM_L_X10Y150_SLICE_X13Y150_CQ),
.O5(CLBLL_L_X4Y148_SLICE_X5Y148_CO5),
.O6(CLBLL_L_X4Y148_SLICE_X5Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeeef000feeef000)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_BLUT (
.I0(CLBLL_L_X4Y150_SLICE_X5Y150_DQ),
.I1(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I2(CLBLM_L_X8Y147_SLICE_X10Y147_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y152_SLICE_X6Y152_CO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y148_SLICE_X5Y148_BO5),
.O6(CLBLL_L_X4Y148_SLICE_X5Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbfff8000bf0080)
  ) CLBLL_L_X4Y148_SLICE_X5Y148_ALUT (
.I0(CLBLL_L_X4Y148_SLICE_X5Y148_AQ),
.I1(CLBLL_L_X4Y151_SLICE_X4Y151_BQ),
.I2(CLBLM_L_X10Y151_SLICE_X12Y151_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y152_SLICE_X15Y152_DQ),
.I5(CLBLL_L_X4Y150_SLICE_X5Y150_BQ),
.O5(CLBLL_L_X4Y148_SLICE_X5Y148_AO5),
.O6(CLBLL_L_X4Y148_SLICE_X5Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y148_SLICE_X4Y148_BO6),
.Q(CLBLL_L_X4Y149_SLICE_X4Y149_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X4Y149_AO6),
.Q(CLBLL_L_X4Y149_SLICE_X4Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X4Y149_BO6),
.Q(CLBLL_L_X4Y149_SLICE_X4Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf040f040f0f0f0f0)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_DLUT (
.I0(CLBLL_L_X4Y151_SLICE_X4Y151_C5Q),
.I1(CLBLM_R_X3Y151_SLICE_X2Y151_AQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X5Y149_SLICE_X6Y149_B5Q),
.I4(1'b1),
.I5(CLBLM_L_X10Y154_SLICE_X13Y154_CQ),
.O5(CLBLL_L_X4Y149_SLICE_X4Y149_DO5),
.O6(CLBLL_L_X4Y149_SLICE_X4Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccffffcfcdffff)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_CLUT (
.I0(CLBLL_L_X4Y152_SLICE_X4Y152_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(LIOB33_X0Y53_IOB_X0Y53_I),
.I3(CLBLL_L_X4Y151_SLICE_X4Y151_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X5Y149_SLICE_X6Y149_A5Q),
.O5(CLBLL_L_X4Y149_SLICE_X4Y149_CO5),
.O6(CLBLL_L_X4Y149_SLICE_X4Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000aa0088)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_BLUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I1(CLBLL_L_X4Y149_SLICE_X4Y149_BQ),
.I2(CLBLL_L_X4Y151_SLICE_X4Y151_C5Q),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X11Y148_SLICE_X15Y148_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y149_SLICE_X4Y149_BO5),
.O6(CLBLL_L_X4Y149_SLICE_X4Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000fcfcf0f0)
  ) CLBLL_L_X4Y149_SLICE_X4Y149_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y149_SLICE_X4Y149_AQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y146_SLICE_X12Y146_CQ),
.I5(CLBLL_L_X4Y149_SLICE_X4Y149_CO6),
.O5(CLBLL_L_X4Y149_SLICE_X4Y149_AO5),
.O6(CLBLL_L_X4Y149_SLICE_X4Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X5Y149_BO6),
.Q(CLBLL_L_X4Y149_SLICE_X5Y149_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y149_SLICE_X5Y149_AO6),
.Q(CLBLL_L_X4Y149_SLICE_X5Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdc50dc50ffffdc50)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_DLUT (
.I0(CLBLL_L_X4Y149_SLICE_X5Y149_CO5),
.I1(CLBLM_R_X3Y155_SLICE_X2Y155_BO6),
.I2(CLBLL_L_X4Y154_SLICE_X5Y154_CO6),
.I3(CLBLL_L_X4Y147_SLICE_X5Y147_AQ),
.I4(CLBLL_L_X4Y153_SLICE_X4Y153_BO6),
.I5(CLBLM_L_X10Y149_SLICE_X13Y149_A5Q),
.O5(CLBLL_L_X4Y149_SLICE_X5Y149_DO5),
.O6(CLBLL_L_X4Y149_SLICE_X5Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7f50000ccffffff)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_CLUT (
.I0(CLBLM_R_X7Y153_SLICE_X8Y153_AQ),
.I1(CLBLM_L_X8Y148_SLICE_X11Y148_BQ),
.I2(CLBLL_L_X4Y150_SLICE_X5Y150_C5Q),
.I3(CLBLL_L_X4Y151_SLICE_X5Y151_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y149_SLICE_X5Y149_CO5),
.O6(CLBLL_L_X4Y149_SLICE_X5Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d8cc000000)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y150_SLICE_X5Y150_AQ),
.I2(RIOB33_X105Y127_IOB_X1Y127_I),
.I3(CLBLM_R_X5Y149_SLICE_X6Y149_DO6),
.I4(CLBLL_L_X4Y150_SLICE_X5Y150_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y149_SLICE_X5Y149_BO5),
.O6(CLBLL_L_X4Y149_SLICE_X5Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcfffc00fc00fc)
  ) CLBLL_L_X4Y149_SLICE_X5Y149_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y153_SLICE_X8Y153_AQ),
.I2(CLBLL_L_X4Y149_SLICE_X5Y149_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(LIOB33_X0Y79_IOB_X0Y79_I),
.O5(CLBLL_L_X4Y149_SLICE_X5Y149_AO5),
.O6(CLBLL_L_X4Y149_SLICE_X5Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y150_SLICE_X4Y150_AO6),
.Q(CLBLL_L_X4Y150_SLICE_X4Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y150_SLICE_X4Y150_BO6),
.Q(CLBLL_L_X4Y150_SLICE_X4Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y150_SLICE_X4Y150_CO6),
.Q(CLBLL_L_X4Y150_SLICE_X4Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff23ff00ff)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_DLUT (
.I0(CLBLM_L_X8Y148_SLICE_X11Y148_BQ),
.I1(CLBLL_L_X4Y150_SLICE_X5Y150_C5Q),
.I2(CLBLL_L_X4Y151_SLICE_X5Y151_CQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X7Y153_SLICE_X8Y153_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y150_SLICE_X4Y150_DO5),
.O6(CLBLL_L_X4Y150_SLICE_X4Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0003300cc)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y151_SLICE_X9Y151_BQ),
.I2(CLBLM_R_X5Y148_SLICE_X7Y148_B5Q),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X8Y150_SLICE_X10Y150_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y150_SLICE_X4Y150_CO5),
.O6(CLBLL_L_X4Y150_SLICE_X4Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00eeeee0e0)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_BLUT (
.I0(CLBLM_L_X8Y150_SLICE_X10Y150_DO6),
.I1(CLBLL_L_X4Y150_SLICE_X4Y150_BQ),
.I2(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y150_SLICE_X4Y150_BO5),
.O6(CLBLL_L_X4Y150_SLICE_X4Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccf0aaaaaa)
  ) CLBLL_L_X4Y150_SLICE_X4Y150_ALUT (
.I0(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.I1(CLBLL_L_X4Y150_SLICE_X4Y150_BQ),
.I2(CLBLL_L_X4Y150_SLICE_X4Y150_AQ),
.I3(CLBLL_L_X4Y151_SLICE_X4Y151_BQ),
.I4(CLBLM_L_X10Y151_SLICE_X12Y151_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y150_SLICE_X4Y150_AO5),
.O6(CLBLL_L_X4Y150_SLICE_X4Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y150_SLICE_X5Y150_CO5),
.Q(CLBLL_L_X4Y150_SLICE_X5Y150_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_D5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y150_SLICE_X5Y150_DO5),
.Q(CLBLL_L_X4Y150_SLICE_X5Y150_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y150_SLICE_X5Y150_AO6),
.Q(CLBLL_L_X4Y150_SLICE_X5Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y150_SLICE_X5Y150_BO6),
.Q(CLBLL_L_X4Y150_SLICE_X5Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y150_SLICE_X5Y150_CO6),
.Q(CLBLL_L_X4Y150_SLICE_X5Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y150_SLICE_X5Y150_DO6),
.Q(CLBLL_L_X4Y150_SLICE_X5Y150_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha3a3a0a0fff00f00)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_DLUT (
.I0(CLBLL_L_X4Y155_SLICE_X5Y155_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y149_SLICE_X4Y149_A5Q),
.I4(CLBLM_R_X5Y148_SLICE_X6Y148_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y150_SLICE_X5Y150_DO5),
.O6(CLBLL_L_X4Y150_SLICE_X5Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff000f0cc55cc55)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_CLUT (
.I0(CLBLM_L_X12Y155_SLICE_X16Y155_CO6),
.I1(CLBLM_R_X13Y151_SLICE_X18Y151_AQ),
.I2(CLBLM_R_X5Y155_SLICE_X6Y155_DO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y149_SLICE_X4Y149_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y150_SLICE_X5Y150_CO5),
.O6(CLBLL_L_X4Y150_SLICE_X5Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00003c003c00)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y150_SLICE_X5Y150_BQ),
.I2(CLBLM_R_X5Y149_SLICE_X6Y149_DO6),
.I3(CLBLM_L_X10Y149_SLICE_X12Y149_DO5),
.I4(CLBLM_R_X5Y157_SLICE_X6Y157_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y150_SLICE_X5Y150_BO5),
.O6(CLBLL_L_X4Y150_SLICE_X5Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa3c00f000)
  ) CLBLL_L_X4Y150_SLICE_X5Y150_ALUT (
.I0(CLBLM_R_X5Y152_SLICE_X7Y152_CQ),
.I1(CLBLL_L_X4Y150_SLICE_X5Y150_BQ),
.I2(CLBLL_L_X4Y150_SLICE_X5Y150_AQ),
.I3(CLBLM_L_X10Y149_SLICE_X12Y149_DO5),
.I4(CLBLM_R_X5Y149_SLICE_X6Y149_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y150_SLICE_X5Y150_AO5),
.O6(CLBLL_L_X4Y150_SLICE_X5Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y151_SLICE_X4Y151_CO5),
.Q(CLBLL_L_X4Y151_SLICE_X4Y151_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_D5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y151_SLICE_X4Y151_DO5),
.Q(CLBLL_L_X4Y151_SLICE_X4Y151_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y151_SLICE_X4Y151_AO6),
.Q(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y151_SLICE_X4Y151_BO6),
.Q(CLBLL_L_X4Y151_SLICE_X4Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y151_SLICE_X4Y151_CO6),
.Q(CLBLL_L_X4Y151_SLICE_X4Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y151_SLICE_X4Y151_DO6),
.Q(CLBLL_L_X4Y151_SLICE_X4Y151_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000aaccaacc)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_DLUT (
.I0(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I1(CLBLM_R_X3Y155_SLICE_X2Y155_BO6),
.I2(CLBLM_L_X10Y149_SLICE_X12Y149_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y154_SLICE_X5Y154_BO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y151_SLICE_X4Y151_DO5),
.O6(CLBLL_L_X4Y151_SLICE_X4Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaaaff00f0f0)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_CLUT (
.I0(CLBLL_L_X4Y152_SLICE_X4Y152_AQ),
.I1(CLBLM_R_X5Y151_SLICE_X7Y151_BQ),
.I2(CLBLM_R_X3Y151_SLICE_X2Y151_AQ),
.I3(CLBLL_L_X4Y158_SLICE_X5Y158_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y151_SLICE_X4Y151_CO5),
.O6(CLBLL_L_X4Y151_SLICE_X4Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cf03cc00cf03)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y151_SLICE_X12Y151_CQ),
.I3(CLBLL_L_X4Y151_SLICE_X4Y151_D5Q),
.I4(CLBLL_L_X4Y150_SLICE_X5Y150_D5Q),
.I5(1'b1),
.O5(CLBLL_L_X4Y151_SLICE_X4Y151_BO5),
.O6(CLBLL_L_X4Y151_SLICE_X4Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000eeec2220)
  ) CLBLL_L_X4Y151_SLICE_X4Y151_ALUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.I3(CLBLM_R_X13Y150_SLICE_X18Y150_CQ),
.I4(CLBLL_L_X4Y152_SLICE_X4Y152_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLL_L_X4Y151_SLICE_X4Y151_AO5),
.O6(CLBLL_L_X4Y151_SLICE_X4Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y151_SLICE_X5Y151_AO6),
.Q(CLBLL_L_X4Y151_SLICE_X5Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y151_SLICE_X5Y151_BO6),
.Q(CLBLL_L_X4Y151_SLICE_X5Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y151_SLICE_X5Y151_CO6),
.Q(CLBLL_L_X4Y151_SLICE_X5Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f330f00bfbbafaa)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_DLUT (
.I0(CLBLM_R_X5Y147_SLICE_X6Y147_BQ),
.I1(CLBLL_L_X2Y153_SLICE_X1Y153_AO5),
.I2(CLBLL_L_X4Y157_SLICE_X4Y157_BO6),
.I3(CLBLL_L_X4Y152_SLICE_X5Y152_BQ),
.I4(LIOB33_X0Y65_IOB_X0Y65_I),
.I5(CLBLM_R_X3Y151_SLICE_X2Y151_CO5),
.O5(CLBLL_L_X4Y151_SLICE_X5Y151_DO5),
.O6(CLBLL_L_X4Y151_SLICE_X5Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb888888888888888)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_CLUT (
.I0(CLBLM_R_X7Y151_SLICE_X9Y151_C5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y156_SLICE_X4Y156_AQ),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_AQ),
.I4(CLBLM_R_X3Y151_SLICE_X3Y151_AQ),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.O5(CLBLL_L_X4Y151_SLICE_X5Y151_CO5),
.O6(CLBLL_L_X4Y151_SLICE_X5Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaff00cccc)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_BLUT (
.I0(CLBLM_L_X12Y149_SLICE_X16Y149_DQ),
.I1(CLBLL_L_X4Y151_SLICE_X5Y151_BQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y150_SLICE_X11Y150_AQ),
.I4(CLBLM_R_X5Y152_SLICE_X6Y152_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLL_L_X4Y151_SLICE_X5Y151_BO5),
.O6(CLBLL_L_X4Y151_SLICE_X5Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcfcfcff000000)
  ) CLBLL_L_X4Y151_SLICE_X5Y151_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y151_SLICE_X9Y151_BQ),
.I2(CLBLL_L_X4Y151_SLICE_X5Y151_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X12Y151_SLICE_X16Y151_C5Q),
.I5(CLBLM_R_X5Y152_SLICE_X6Y152_CO6),
.O5(CLBLL_L_X4Y151_SLICE_X5Y151_AO5),
.O6(CLBLL_L_X4Y151_SLICE_X5Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y152_SLICE_X4Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y152_SLICE_X4Y152_AO6),
.Q(CLBLL_L_X4Y152_SLICE_X4Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff005033730050)
  ) CLBLL_L_X4Y152_SLICE_X4Y152_DLUT (
.I0(CLBLL_L_X4Y157_SLICE_X4Y157_CO6),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(LIOB33_X0Y65_IOB_X0Y66_I),
.I3(CLBLL_L_X2Y155_SLICE_X1Y155_CO6),
.I4(CLBLM_R_X5Y149_SLICE_X6Y149_BQ),
.I5(RIOB33_X105Y129_IOB_X1Y129_I),
.O5(CLBLL_L_X4Y152_SLICE_X4Y152_DO5),
.O6(CLBLL_L_X4Y152_SLICE_X4Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0300000003000a0a)
  ) CLBLL_L_X4Y152_SLICE_X4Y152_CLUT (
.I0(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.I1(CLBLL_L_X2Y155_SLICE_X1Y155_CO6),
.I2(CLBLM_R_X3Y158_SLICE_X2Y158_AO5),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(CLBLL_L_X2Y155_SLICE_X1Y155_CO5),
.O5(CLBLL_L_X4Y152_SLICE_X4Y152_CO5),
.O6(CLBLL_L_X4Y152_SLICE_X4Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffefffee)
  ) CLBLL_L_X4Y152_SLICE_X4Y152_BLUT (
.I0(CLBLL_L_X4Y152_SLICE_X4Y152_DO6),
.I1(CLBLL_L_X4Y152_SLICE_X5Y152_DO6),
.I2(CLBLM_R_X3Y151_SLICE_X2Y151_CO5),
.I3(CLBLM_R_X5Y152_SLICE_X6Y152_DO6),
.I4(CLBLM_R_X7Y153_SLICE_X9Y153_BQ),
.I5(CLBLL_L_X4Y152_SLICE_X4Y152_CO6),
.O5(CLBLL_L_X4Y152_SLICE_X4Y152_BO5),
.O6(CLBLL_L_X4Y152_SLICE_X4Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccca000cccc0000)
  ) CLBLL_L_X4Y152_SLICE_X4Y152_ALUT (
.I0(CLBLM_R_X7Y155_SLICE_X9Y155_A5Q),
.I1(CLBLM_L_X12Y149_SLICE_X16Y149_AQ),
.I2(CLBLL_L_X4Y155_SLICE_X4Y155_AQ),
.I3(CLBLL_L_X4Y155_SLICE_X4Y155_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y149_SLICE_X4Y149_AQ),
.O5(CLBLL_L_X4Y152_SLICE_X4Y152_AO5),
.O6(CLBLL_L_X4Y152_SLICE_X4Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y152_SLICE_X5Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y152_SLICE_X5Y152_AO6),
.Q(CLBLL_L_X4Y152_SLICE_X5Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y152_SLICE_X5Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y152_SLICE_X5Y152_BO6),
.Q(CLBLL_L_X4Y152_SLICE_X5Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y152_SLICE_X5Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y152_SLICE_X5Y152_CO6),
.Q(CLBLL_L_X4Y152_SLICE_X5Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000022f200002222)
  ) CLBLL_L_X4Y152_SLICE_X5Y152_DLUT (
.I0(CLBLM_R_X5Y149_SLICE_X7Y149_BQ),
.I1(CLBLM_R_X3Y156_SLICE_X3Y156_AO5),
.I2(CLBLL_L_X4Y148_SLICE_X5Y148_CQ),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLL_L_X4Y157_SLICE_X4Y157_CO5),
.I5(CLBLL_L_X4Y157_SLICE_X5Y157_AO6),
.O5(CLBLL_L_X4Y152_SLICE_X5Y152_DO5),
.O6(CLBLL_L_X4Y152_SLICE_X5Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55aa00ee44aa00)
  ) CLBLL_L_X4Y152_SLICE_X5Y152_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y152_SLICE_X5Y152_CQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y151_SLICE_X5Y151_BQ),
.I4(CLBLL_L_X4Y147_SLICE_X4Y147_BO6),
.I5(CLBLM_L_X8Y153_SLICE_X11Y153_C5Q),
.O5(CLBLL_L_X4Y152_SLICE_X5Y152_CO5),
.O6(CLBLL_L_X4Y152_SLICE_X5Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa8a8a8ffa8a8a8)
  ) CLBLL_L_X4Y152_SLICE_X5Y152_BLUT (
.I0(CLBLM_R_X5Y152_SLICE_X6Y152_CO6),
.I1(CLBLL_L_X4Y152_SLICE_X5Y152_BQ),
.I2(CLBLM_R_X5Y150_SLICE_X6Y150_AQ),
.I3(CLBLM_R_X7Y152_SLICE_X9Y152_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y152_SLICE_X5Y152_BO5),
.O6(CLBLL_L_X4Y152_SLICE_X5Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf5ccffcca0cc00)
  ) CLBLL_L_X4Y152_SLICE_X5Y152_ALUT (
.I0(CLBLL_L_X4Y151_SLICE_X4Y151_BQ),
.I1(CLBLL_L_X4Y148_SLICE_X5Y148_CQ),
.I2(CLBLL_L_X4Y152_SLICE_X5Y152_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y151_SLICE_X12Y151_CQ),
.I5(CLBLM_L_X10Y148_SLICE_X13Y148_BQ),
.O5(CLBLL_L_X4Y152_SLICE_X5Y152_AO5),
.O6(CLBLL_L_X4Y152_SLICE_X5Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafaaaaffafffaa)
  ) CLBLL_L_X4Y153_SLICE_X4Y153_DLUT (
.I0(CLBLL_L_X4Y153_SLICE_X5Y153_BO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y153_SLICE_X2Y153_CO6),
.I3(CLBLM_R_X7Y155_SLICE_X9Y155_A5Q),
.I4(RIOB33_X105Y115_IOB_X1Y116_I),
.I5(CLBLM_R_X3Y153_SLICE_X2Y153_AO6),
.O5(CLBLL_L_X4Y153_SLICE_X4Y153_DO5),
.O6(CLBLL_L_X4Y153_SLICE_X4Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8fff88ff8f8f8888)
  ) CLBLL_L_X4Y153_SLICE_X4Y153_CLUT (
.I0(CLBLM_R_X5Y149_SLICE_X6Y149_BQ),
.I1(CLBLM_R_X3Y152_SLICE_X3Y152_AO6),
.I2(CLBLL_L_X2Y153_SLICE_X1Y153_AO5),
.I3(CLBLM_R_X3Y151_SLICE_X2Y151_CO5),
.I4(LIOB33_X0Y65_IOB_X0Y66_I),
.I5(CLBLM_R_X7Y153_SLICE_X9Y153_BQ),
.O5(CLBLL_L_X4Y153_SLICE_X4Y153_CO5),
.O6(CLBLL_L_X4Y153_SLICE_X4Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffff1)
  ) CLBLL_L_X4Y153_SLICE_X4Y153_BLUT (
.I0(CLBLM_R_X3Y154_SLICE_X3Y154_DO6),
.I1(CLBLM_R_X3Y155_SLICE_X2Y155_DO6),
.I2(CLBLM_R_X5Y153_SLICE_X6Y153_DO6),
.I3(CLBLM_R_X5Y154_SLICE_X7Y154_CO6),
.I4(CLBLL_L_X4Y152_SLICE_X5Y152_DO6),
.I5(CLBLL_L_X4Y153_SLICE_X4Y153_CO6),
.O5(CLBLL_L_X4Y153_SLICE_X4Y153_BO5),
.O6(CLBLL_L_X4Y153_SLICE_X4Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLL_L_X4Y153_SLICE_X4Y153_ALUT (
.I0(CLBLL_L_X4Y153_SLICE_X4Y153_DO6),
.I1(CLBLL_L_X4Y154_SLICE_X4Y154_DO6),
.I2(CLBLM_R_X5Y156_SLICE_X7Y156_DO6),
.I3(CLBLM_R_X3Y151_SLICE_X2Y151_DO6),
.I4(CLBLM_R_X3Y155_SLICE_X3Y155_DO6),
.I5(CLBLM_R_X5Y153_SLICE_X6Y153_CO6),
.O5(CLBLL_L_X4Y153_SLICE_X4Y153_AO5),
.O6(CLBLL_L_X4Y153_SLICE_X4Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y153_SLICE_X5Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y153_SLICE_X5Y153_AO6),
.Q(CLBLL_L_X4Y153_SLICE_X5Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3b3b3b3b0a0a0a0a)
  ) CLBLL_L_X4Y153_SLICE_X5Y153_DLUT (
.I0(CLBLL_L_X4Y150_SLICE_X4Y150_AQ),
.I1(CLBLM_R_X5Y153_SLICE_X6Y153_BO5),
.I2(CLBLL_L_X2Y155_SLICE_X1Y155_BO5),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X13Y153_SLICE_X18Y153_C5Q),
.O5(CLBLL_L_X4Y153_SLICE_X5Y153_DO5),
.O6(CLBLL_L_X4Y153_SLICE_X5Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4fff4f4f44ff4444)
  ) CLBLL_L_X4Y153_SLICE_X5Y153_CLUT (
.I0(CLBLM_R_X3Y154_SLICE_X3Y154_AO6),
.I1(CLBLL_L_X4Y148_SLICE_X5Y148_BQ),
.I2(CLBLM_R_X3Y157_SLICE_X2Y157_AO6),
.I3(CLBLL_L_X4Y156_SLICE_X4Y156_CO6),
.I4(CLBLM_R_X5Y150_SLICE_X6Y150_DQ),
.I5(RIOB33_X105Y109_IOB_X1Y110_I),
.O5(CLBLL_L_X4Y153_SLICE_X5Y153_CO5),
.O6(CLBLL_L_X4Y153_SLICE_X5Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcd05cdcdcc00cccc)
  ) CLBLL_L_X4Y153_SLICE_X5Y153_BLUT (
.I0(CLBLM_R_X3Y156_SLICE_X3Y156_AO5),
.I1(CLBLM_R_X7Y155_SLICE_X8Y155_A5Q),
.I2(CLBLL_L_X4Y157_SLICE_X4Y157_CO6),
.I3(RIOB33_X105Y129_IOB_X1Y129_I),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(CLBLM_R_X7Y147_SLICE_X8Y147_AQ),
.O5(CLBLL_L_X4Y153_SLICE_X5Y153_BO5),
.O6(CLBLL_L_X4Y153_SLICE_X5Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf055f000f055f000)
  ) CLBLL_L_X4Y153_SLICE_X5Y153_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(CLBLL_L_X4Y150_SLICE_X4Y150_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y152_SLICE_X7Y152_DQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y153_SLICE_X5Y153_AO5),
.O6(CLBLL_L_X4Y153_SLICE_X5Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f0f5f0f55005500)
  ) CLBLL_L_X4Y154_SLICE_X4Y154_DLUT (
.I0(CLBLM_R_X3Y153_SLICE_X3Y153_AO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y154_SLICE_X3Y154_AO5),
.I3(CLBLM_L_X8Y154_SLICE_X11Y154_BQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y154_SLICE_X15Y154_AQ),
.O5(CLBLL_L_X4Y154_SLICE_X4Y154_DO5),
.O6(CLBLL_L_X4Y154_SLICE_X4Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3fff0fff3f3f0f0)
  ) CLBLL_L_X4Y154_SLICE_X4Y154_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y156_SLICE_X4Y156_CO6),
.I2(CLBLL_L_X4Y155_SLICE_X4Y155_DO6),
.I3(CLBLL_L_X4Y157_SLICE_X4Y157_BO5),
.I4(CLBLM_R_X11Y151_SLICE_X15Y151_BQ),
.I5(CLBLM_R_X7Y154_SLICE_X9Y154_BQ),
.O5(CLBLL_L_X4Y154_SLICE_X4Y154_CO5),
.O6(CLBLL_L_X4Y154_SLICE_X4Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLL_L_X4Y154_SLICE_X4Y154_BLUT (
.I0(CLBLM_R_X3Y153_SLICE_X3Y153_DO6),
.I1(CLBLM_R_X3Y155_SLICE_X3Y155_DO6),
.I2(CLBLL_L_X4Y156_SLICE_X5Y156_CO6),
.I3(CLBLM_R_X3Y153_SLICE_X3Y153_CO6),
.I4(CLBLM_R_X5Y154_SLICE_X6Y154_BO6),
.I5(CLBLL_L_X4Y154_SLICE_X4Y154_CO6),
.O5(CLBLL_L_X4Y154_SLICE_X4Y154_BO5),
.O6(CLBLL_L_X4Y154_SLICE_X4Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLL_L_X4Y154_SLICE_X4Y154_ALUT (
.I0(CLBLM_R_X3Y155_SLICE_X3Y155_AO6),
.I1(CLBLM_R_X7Y155_SLICE_X9Y155_DO6),
.I2(CLBLM_R_X5Y156_SLICE_X6Y156_AO6),
.I3(CLBLL_L_X4Y152_SLICE_X4Y152_BO6),
.I4(CLBLM_R_X3Y154_SLICE_X3Y154_BO6),
.I5(CLBLM_R_X5Y154_SLICE_X7Y154_CO6),
.O5(CLBLL_L_X4Y154_SLICE_X4Y154_AO5),
.O6(CLBLL_L_X4Y154_SLICE_X4Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y154_SLICE_X5Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y154_SLICE_X5Y154_AO6),
.Q(CLBLL_L_X4Y154_SLICE_X5Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd5d5d5c0c0d5c0c0)
  ) CLBLL_L_X4Y154_SLICE_X5Y154_DLUT (
.I0(CLBLM_R_X3Y153_SLICE_X3Y153_AO5),
.I1(CLBLL_L_X4Y155_SLICE_X5Y155_A5Q),
.I2(CLBLM_R_X3Y152_SLICE_X3Y152_AO6),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLM_R_X7Y154_SLICE_X8Y154_CQ),
.I5(CLBLM_R_X11Y154_SLICE_X14Y154_D5Q),
.O5(CLBLL_L_X4Y154_SLICE_X5Y154_DO5),
.O6(CLBLL_L_X4Y154_SLICE_X5Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLL_L_X4Y154_SLICE_X5Y154_CLUT (
.I0(CLBLM_R_X3Y154_SLICE_X3Y154_CO6),
.I1(CLBLL_L_X4Y153_SLICE_X5Y153_CO6),
.I2(CLBLM_R_X5Y154_SLICE_X7Y154_DO6),
.I3(CLBLM_R_X5Y154_SLICE_X6Y154_DO6),
.I4(CLBLL_L_X4Y154_SLICE_X5Y154_DO6),
.I5(CLBLL_L_X4Y151_SLICE_X5Y151_DO6),
.O5(CLBLL_L_X4Y154_SLICE_X5Y154_CO5),
.O6(CLBLL_L_X4Y154_SLICE_X5Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLL_L_X4Y154_SLICE_X5Y154_BLUT (
.I0(CLBLM_R_X5Y154_SLICE_X6Y154_CO6),
.I1(CLBLM_R_X3Y155_SLICE_X3Y155_DO6),
.I2(CLBLL_L_X4Y153_SLICE_X5Y153_DO6),
.I3(CLBLM_R_X5Y155_SLICE_X7Y155_DO6),
.I4(CLBLM_R_X5Y157_SLICE_X6Y157_DO6),
.I5(CLBLM_R_X3Y151_SLICE_X3Y151_CO6),
.O5(CLBLL_L_X4Y154_SLICE_X5Y154_BO5),
.O6(CLBLL_L_X4Y154_SLICE_X5Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb11ba10bb11ba10)
  ) CLBLL_L_X4Y154_SLICE_X5Y154_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y152_SLICE_X6Y152_CO5),
.I2(CLBLL_L_X4Y154_SLICE_X5Y154_AQ),
.I3(CLBLM_R_X7Y154_SLICE_X8Y154_AQ),
.I4(CLBLM_R_X5Y152_SLICE_X7Y152_DQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y154_SLICE_X5Y154_AO5),
.O6(CLBLL_L_X4Y154_SLICE_X5Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y155_SLICE_X4Y155_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y155_SLICE_X4Y155_AO6),
.Q(CLBLL_L_X4Y155_SLICE_X4Y155_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y155_SLICE_X4Y155_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y155_SLICE_X4Y155_BO6),
.Q(CLBLL_L_X4Y155_SLICE_X4Y155_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0032003200020002)
  ) CLBLL_L_X4Y155_SLICE_X4Y155_DLUT (
.I0(CLBLL_L_X4Y154_SLICE_X5Y154_AQ),
.I1(CLBLM_R_X3Y158_SLICE_X2Y158_AO5),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(CLBLL_L_X2Y155_SLICE_X1Y155_CO6),
.I4(1'b1),
.I5(RIOB33_X105Y107_IOB_X1Y107_I),
.O5(CLBLL_L_X4Y155_SLICE_X4Y155_DO5),
.O6(CLBLL_L_X4Y155_SLICE_X4Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff007f807f80)
  ) CLBLL_L_X4Y155_SLICE_X4Y155_CLUT (
.I0(CLBLM_R_X3Y151_SLICE_X3Y151_AQ),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_AQ),
.I3(CLBLL_L_X4Y156_SLICE_X4Y156_AQ),
.I4(1'b1),
.I5(CLBLM_L_X12Y155_SLICE_X16Y155_CO6),
.O5(CLBLL_L_X4Y155_SLICE_X4Y155_CO5),
.O6(CLBLL_L_X4Y155_SLICE_X4Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000fcfccccc)
  ) CLBLL_L_X4Y155_SLICE_X4Y155_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y155_SLICE_X4Y155_BQ),
.I2(CLBLM_R_X5Y153_SLICE_X6Y153_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y149_SLICE_X4Y149_CO6),
.O5(CLBLL_L_X4Y155_SLICE_X4Y155_BO5),
.O6(CLBLL_L_X4Y155_SLICE_X4Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00fcf0fcf0)
  ) CLBLL_L_X4Y155_SLICE_X4Y155_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y155_SLICE_X4Y155_AQ),
.I3(CLBLM_R_X7Y155_SLICE_X8Y155_A5Q),
.I4(1'b1),
.I5(CLBLL_L_X4Y149_SLICE_X4Y149_CO6),
.O5(CLBLL_L_X4Y155_SLICE_X4Y155_AO5),
.O6(CLBLL_L_X4Y155_SLICE_X4Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y155_SLICE_X5Y155_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y155_SLICE_X5Y155_AO5),
.Q(CLBLL_L_X4Y155_SLICE_X5Y155_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y155_SLICE_X5Y155_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y155_SLICE_X5Y155_AO6),
.Q(CLBLL_L_X4Y155_SLICE_X5Y155_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y155_SLICE_X5Y155_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y155_SLICE_X5Y155_BO6),
.Q(CLBLL_L_X4Y155_SLICE_X5Y155_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1010005510100000)
  ) CLBLL_L_X4Y155_SLICE_X5Y155_DLUT (
.I0(CLBLM_R_X3Y158_SLICE_X2Y158_AO5),
.I1(CLBLL_L_X2Y155_SLICE_X1Y155_CO6),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(CLBLL_L_X2Y155_SLICE_X1Y155_AO5),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(CLBLL_L_X4Y151_SLICE_X5Y151_BQ),
.O5(CLBLL_L_X4Y155_SLICE_X5Y155_DO5),
.O6(CLBLL_L_X4Y155_SLICE_X5Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f222ff00ff22)
  ) CLBLL_L_X4Y155_SLICE_X5Y155_CLUT (
.I0(CLBLL_L_X4Y155_SLICE_X5Y155_BQ),
.I1(CLBLM_R_X3Y156_SLICE_X3Y156_AO5),
.I2(RIOB33_X105Y129_IOB_X1Y129_I),
.I3(CLBLL_L_X4Y150_SLICE_X5Y150_CQ),
.I4(CLBLL_L_X4Y157_SLICE_X4Y157_CO6),
.I5(RIOB33_X105Y137_IOB_X1Y137_I),
.O5(CLBLL_L_X4Y155_SLICE_X5Y155_CO5),
.O6(CLBLL_L_X4Y155_SLICE_X5Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fffc00000f0c)
  ) CLBLL_L_X4Y155_SLICE_X5Y155_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y155_SLICE_X5Y155_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y146_SLICE_X5Y146_AQ),
.I4(CLBLL_L_X4Y147_SLICE_X4Y147_BO6),
.I5(CLBLL_L_X4Y155_SLICE_X5Y155_A5Q),
.O5(CLBLL_L_X4Y155_SLICE_X5Y155_BO5),
.O6(CLBLL_L_X4Y155_SLICE_X5Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2e2e2ff33cc00)
  ) CLBLL_L_X4Y155_SLICE_X5Y155_ALUT (
.I0(CLBLM_R_X3Y156_SLICE_X2Y156_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y155_SLICE_X14Y155_BQ),
.I3(CLBLM_R_X7Y155_SLICE_X9Y155_BQ),
.I4(CLBLL_L_X4Y154_SLICE_X5Y154_CO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y155_SLICE_X5Y155_AO5),
.O6(CLBLL_L_X4Y155_SLICE_X5Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y156_SLICE_X4Y156_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLL_L_X4Y156_SLICE_X4Y156_AO6),
.Q(CLBLL_L_X4Y156_SLICE_X4Y156_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000080)
  ) CLBLL_L_X4Y156_SLICE_X4Y156_DLUT (
.I0(CLBLM_L_X8Y154_SLICE_X11Y154_AQ),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(CLBLL_L_X4Y157_SLICE_X4Y157_CO5),
.O5(CLBLL_L_X4Y156_SLICE_X4Y156_DO5),
.O6(CLBLL_L_X4Y156_SLICE_X4Y156_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffbfffbffffff)
  ) CLBLL_L_X4Y156_SLICE_X4Y156_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLM_R_X3Y158_SLICE_X2Y158_AO6),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y156_SLICE_X4Y156_CO5),
.O6(CLBLL_L_X4Y156_SLICE_X4Y156_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffeffffffe55)
  ) CLBLL_L_X4Y156_SLICE_X4Y156_BLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(CLBLL_L_X4Y157_SLICE_X4Y157_CO5),
.I5(1'b1),
.O5(CLBLL_L_X4Y156_SLICE_X4Y156_BO5),
.O6(CLBLL_L_X4Y156_SLICE_X4Y156_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00fcf022222222)
  ) CLBLL_L_X4Y156_SLICE_X4Y156_ALUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLL_L_X4Y155_SLICE_X4Y155_CO6),
.I3(CLBLL_L_X4Y154_SLICE_X5Y154_AQ),
.I4(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y156_SLICE_X4Y156_AO5),
.O6(CLBLL_L_X4Y156_SLICE_X4Y156_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00003f0f00003300)
  ) CLBLL_L_X4Y156_SLICE_X5Y156_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y155_SLICE_X1Y155_CO6),
.I2(CLBLL_L_X2Y155_SLICE_X1Y155_CO5),
.I3(LIOB33_X0Y67_IOB_X0Y67_I),
.I4(CLBLL_L_X4Y157_SLICE_X4Y157_CO6),
.I5(CLBLM_R_X7Y156_SLICE_X8Y156_DQ),
.O5(CLBLL_L_X4Y156_SLICE_X5Y156_DO5),
.O6(CLBLL_L_X4Y156_SLICE_X5Y156_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff3f0fbfa)
  ) CLBLL_L_X4Y156_SLICE_X5Y156_CLUT (
.I0(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.I1(CLBLM_R_X3Y154_SLICE_X3Y154_AO6),
.I2(CLBLL_L_X4Y157_SLICE_X5Y157_CO6),
.I3(CLBLM_R_X7Y157_SLICE_X8Y157_DQ),
.I4(CLBLL_L_X4Y156_SLICE_X4Y156_CO5),
.I5(CLBLL_L_X4Y156_SLICE_X5Y156_BO6),
.O5(CLBLL_L_X4Y156_SLICE_X5Y156_CO5),
.O6(CLBLL_L_X4Y156_SLICE_X5Y156_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010000000000)
  ) CLBLL_L_X4Y156_SLICE_X5Y156_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLL_L_X4Y157_SLICE_X4Y157_CO5),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLM_R_X7Y152_SLICE_X9Y152_AQ),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(RIOB33_X105Y133_IOB_X1Y134_I),
.O5(CLBLL_L_X4Y156_SLICE_X5Y156_BO5),
.O6(CLBLL_L_X4Y156_SLICE_X5Y156_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffdc)
  ) CLBLL_L_X4Y156_SLICE_X5Y156_ALUT (
.I0(CLBLL_L_X4Y156_SLICE_X4Y156_CO5),
.I1(CLBLL_L_X4Y155_SLICE_X5Y155_DO6),
.I2(CLBLM_R_X3Y151_SLICE_X3Y151_AQ),
.I3(CLBLM_R_X3Y156_SLICE_X2Y156_CO6),
.I4(CLBLM_R_X5Y158_SLICE_X6Y158_CO6),
.I5(CLBLM_R_X5Y157_SLICE_X6Y157_CO6),
.O5(CLBLL_L_X4Y156_SLICE_X5Y156_AO5),
.O6(CLBLL_L_X4Y156_SLICE_X5Y156_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000400000000000)
  ) CLBLL_L_X4Y157_SLICE_X4Y157_DLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(CLBLM_R_X3Y158_SLICE_X2Y158_AO6),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(CLBLM_L_X8Y152_SLICE_X10Y152_CQ),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLL_L_X4Y157_SLICE_X4Y157_DO5),
.O6(CLBLL_L_X4Y157_SLICE_X4Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffbfffffffffb)
  ) CLBLL_L_X4Y157_SLICE_X4Y157_CLUT (
.I0(RIOB33_X105Y129_IOB_X1Y130_I),
.I1(RIOB33_X105Y137_IOB_X1Y137_I),
.I2(RIOB33_X105Y129_IOB_X1Y129_I),
.I3(RIOB33_X105Y135_IOB_X1Y135_I),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y157_SLICE_X4Y157_CO5),
.O6(CLBLL_L_X4Y157_SLICE_X4Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbfffffffffbf)
  ) CLBLL_L_X4Y157_SLICE_X4Y157_BLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLL_L_X4Y157_SLICE_X4Y157_CO5),
.I5(1'b1),
.O5(CLBLL_L_X4Y157_SLICE_X4Y157_BO5),
.O6(CLBLL_L_X4Y157_SLICE_X4Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaaaaaaaaffff)
  ) CLBLL_L_X4Y157_SLICE_X4Y157_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y157_SLICE_X4Y157_AO5),
.O6(CLBLL_L_X4Y157_SLICE_X4Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y157_SLICE_X5Y157_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y157_SLICE_X5Y157_DO5),
.O6(CLBLL_L_X4Y157_SLICE_X5Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f4ffff00440044)
  ) CLBLL_L_X4Y157_SLICE_X5Y157_CLUT (
.I0(CLBLL_L_X4Y157_SLICE_X4Y157_CO6),
.I1(CLBLM_R_X7Y156_SLICE_X9Y156_CQ),
.I2(RIOB33_X105Y129_IOB_X1Y129_I),
.I3(CLBLM_R_X3Y156_SLICE_X3Y156_AO5),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(CLBLM_L_X8Y156_SLICE_X11Y156_B5Q),
.O5(CLBLL_L_X4Y157_SLICE_X5Y157_CO5),
.O6(CLBLL_L_X4Y157_SLICE_X5Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000005010400)
  ) CLBLL_L_X4Y157_SLICE_X5Y157_BLUT (
.I0(CLBLL_L_X4Y157_SLICE_X4Y157_AO5),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLL_L_X4Y157_SLICE_X4Y157_CO5),
.I3(CLBLM_R_X5Y157_SLICE_X6Y157_AQ),
.I4(CLBLM_R_X5Y157_SLICE_X7Y157_AQ),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLL_L_X4Y157_SLICE_X5Y157_BO5),
.O6(CLBLL_L_X4Y157_SLICE_X5Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h50005000fff5fff5)
  ) CLBLL_L_X4Y157_SLICE_X5Y157_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(1'b1),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y157_SLICE_X5Y157_AO5),
.O6(CLBLL_L_X4Y157_SLICE_X5Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y158_SLICE_X4Y158_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y158_SLICE_X4Y158_DO5),
.O6(CLBLL_L_X4Y158_SLICE_X4Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y158_SLICE_X4Y158_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y158_SLICE_X4Y158_CO5),
.O6(CLBLL_L_X4Y158_SLICE_X4Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y158_SLICE_X4Y158_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y158_SLICE_X4Y158_BO5),
.O6(CLBLL_L_X4Y158_SLICE_X4Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffefffe)
  ) CLBLL_L_X4Y158_SLICE_X4Y158_ALUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(RIOB33_X105Y127_IOB_X1Y128_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLL_L_X4Y157_SLICE_X4Y157_AO6),
.I4(1'b1),
.I5(RIOB33_X105Y129_IOB_X1Y130_I),
.O5(CLBLL_L_X4Y158_SLICE_X4Y158_AO5),
.O6(CLBLL_L_X4Y158_SLICE_X4Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y158_SLICE_X5Y158_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y159_SLICE_X16Y159_CO5),
.Q(CLBLL_L_X4Y158_SLICE_X5Y158_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y158_SLICE_X5Y158_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y158_SLICE_X5Y158_DO5),
.O6(CLBLL_L_X4Y158_SLICE_X5Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y158_SLICE_X5Y158_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y158_SLICE_X5Y158_CO5),
.O6(CLBLL_L_X4Y158_SLICE_X5Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y158_SLICE_X5Y158_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y158_SLICE_X5Y158_BO5),
.O6(CLBLL_L_X4Y158_SLICE_X5Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y158_SLICE_X5Y158_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y158_SLICE_X5Y158_AO5),
.O6(CLBLL_L_X4Y158_SLICE_X5Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y150_SLICE_X54Y150_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y150_SLICE_X54Y150_DO5),
.O6(CLBLL_L_X36Y150_SLICE_X54Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y150_SLICE_X54Y150_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y150_SLICE_X54Y150_CO5),
.O6(CLBLL_L_X36Y150_SLICE_X54Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y150_SLICE_X54Y150_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y150_SLICE_X54Y150_BO5),
.O6(CLBLL_L_X36Y150_SLICE_X54Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000033003300)
  ) CLBLL_L_X36Y150_SLICE_X54Y150_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(1'b1),
.I3(RIOB33_X105Y119_IOB_X1Y119_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y149_SLICE_X9Y149_CQ),
.O5(CLBLL_L_X36Y150_SLICE_X54Y150_AO5),
.O6(CLBLL_L_X36Y150_SLICE_X54Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y150_SLICE_X55Y150_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y150_SLICE_X55Y150_DO5),
.O6(CLBLL_L_X36Y150_SLICE_X55Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y150_SLICE_X55Y150_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y150_SLICE_X55Y150_CO5),
.O6(CLBLL_L_X36Y150_SLICE_X55Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y150_SLICE_X55Y150_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y150_SLICE_X55Y150_BO5),
.O6(CLBLL_L_X36Y150_SLICE_X55Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X36Y150_SLICE_X55Y150_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X36Y150_SLICE_X55Y150_AO5),
.O6(CLBLL_L_X36Y150_SLICE_X55Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_DO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_CO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_BO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00ff)
  ) CLBLL_L_X52Y126_SLICE_X78Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y123_IOB_X1Y124_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X78Y126_AO5),
.O6(CLBLL_L_X52Y126_SLICE_X78Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_DO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_CO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_BO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X52Y126_SLICE_X79Y126_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X52Y126_SLICE_X79Y126_AO5),
.O6(CLBLL_L_X52Y126_SLICE_X79Y126_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X10Y146_BO5),
.Q(CLBLM_L_X8Y146_SLICE_X10Y146_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X10Y146_AO6),
.Q(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X10Y146_BO6),
.Q(CLBLM_L_X8Y146_SLICE_X10Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y146_SLICE_X10Y146_DO5),
.O6(CLBLM_L_X8Y146_SLICE_X10Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y146_SLICE_X10Y146_CO5),
.O6(CLBLM_L_X8Y146_SLICE_X10Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000ccffcc00)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y154_SLICE_X9Y154_BQ),
.I2(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y146_SLICE_X10Y146_BO5),
.O6(CLBLM_L_X8Y146_SLICE_X10Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff220022ff200020)
  ) CLBLM_L_X8Y146_SLICE_X10Y146_ALUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y150_SLICE_X11Y150_BQ),
.I5(CLBLM_R_X11Y146_SLICE_X14Y146_CQ),
.O5(CLBLM_L_X8Y146_SLICE_X10Y146_AO5),
.O6(CLBLM_L_X8Y146_SLICE_X10Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X11Y146_AO6),
.Q(CLBLM_L_X8Y146_SLICE_X11Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X11Y146_BO6),
.Q(CLBLM_L_X8Y146_SLICE_X11Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y146_SLICE_X11Y146_CO6),
.Q(CLBLM_L_X8Y146_SLICE_X11Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y146_SLICE_X11Y146_DO5),
.O6(CLBLM_L_X8Y146_SLICE_X11Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00fc000000fc)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y146_SLICE_X11Y146_CQ),
.I2(CLBLM_L_X8Y146_SLICE_X11Y146_BQ),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y146_SLICE_X10Y146_BQ),
.O5(CLBLM_L_X8Y146_SLICE_X11Y146_CO5),
.O6(CLBLM_L_X8Y146_SLICE_X11Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0f5e4f5e4)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y146_SLICE_X11Y146_BQ),
.I2(CLBLM_L_X8Y148_SLICE_X11Y148_AQ),
.I3(CLBLM_R_X7Y146_SLICE_X9Y146_AQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y146_SLICE_X8Y146_DO6),
.O5(CLBLM_L_X8Y146_SLICE_X11Y146_BO5),
.O6(CLBLM_L_X8Y146_SLICE_X11Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888ddddd8d8)
  ) CLBLM_L_X8Y146_SLICE_X11Y146_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y154_SLICE_X11Y154_BQ),
.I2(CLBLM_L_X8Y146_SLICE_X11Y146_AQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y146_SLICE_X12Y146_AQ),
.I5(CLBLM_R_X7Y146_SLICE_X9Y146_DO6),
.O5(CLBLM_L_X8Y146_SLICE_X11Y146_AO5),
.O6(CLBLM_L_X8Y146_SLICE_X11Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y147_SLICE_X10Y147_AO6),
.Q(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y147_SLICE_X10Y147_BO6),
.Q(CLBLM_L_X8Y147_SLICE_X10Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y147_SLICE_X10Y147_CO6),
.Q(CLBLM_L_X8Y147_SLICE_X10Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3319339980800000)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_DLUT (
.I0(CLBLM_L_X8Y147_SLICE_X10Y147_BQ),
.I1(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.I2(CLBLM_R_X7Y147_SLICE_X9Y147_BQ),
.I3(CLBLM_R_X7Y146_SLICE_X9Y146_DO6),
.I4(CLBLM_R_X7Y147_SLICE_X9Y147_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y147_SLICE_X10Y147_DO5),
.O6(CLBLM_L_X8Y147_SLICE_X10Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00ccaaaa0000)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_CLUT (
.I0(CLBLM_R_X5Y144_SLICE_X6Y144_BQ),
.I1(CLBLM_L_X8Y147_SLICE_X10Y147_CQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y151_SLICE_X9Y151_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y147_SLICE_X10Y147_CO5),
.O6(CLBLM_L_X8Y147_SLICE_X10Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0ffecb3b3)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_BLUT (
.I0(CLBLM_R_X7Y156_SLICE_X8Y156_BQ),
.I1(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y147_SLICE_X10Y147_DO5),
.I4(CLBLM_L_X8Y147_SLICE_X10Y147_BQ),
.I5(CLBLM_L_X8Y147_SLICE_X10Y147_AO5),
.O5(CLBLM_L_X8Y147_SLICE_X10Y147_BO5),
.O6(CLBLM_L_X8Y147_SLICE_X10Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcd01cc00fcfcffff)
  ) CLBLM_L_X8Y147_SLICE_X10Y147_ALUT (
.I0(CLBLM_L_X8Y147_SLICE_X10Y147_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y154_SLICE_X13Y154_CQ),
.I3(CLBLM_L_X10Y148_SLICE_X13Y148_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y147_SLICE_X10Y147_AO5),
.O6(CLBLM_L_X8Y147_SLICE_X10Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y147_SLICE_X11Y147_AO6),
.Q(CLBLM_L_X8Y147_SLICE_X11Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y147_SLICE_X11Y147_BO6),
.Q(CLBLM_L_X8Y147_SLICE_X11Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffdfffdf)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_DLUT (
.I0(CLBLL_L_X4Y154_SLICE_X5Y154_BO6),
.I1(CLBLM_R_X3Y156_SLICE_X2Y156_DO6),
.I2(CLBLM_R_X3Y152_SLICE_X3Y152_BO5),
.I3(CLBLM_R_X7Y148_SLICE_X9Y148_CO5),
.I4(1'b1),
.I5(CLBLM_R_X13Y155_SLICE_X19Y155_AO6),
.O5(CLBLM_L_X8Y147_SLICE_X11Y147_DO5),
.O6(CLBLM_L_X8Y147_SLICE_X11Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000000000000000)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_CLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.I1(CLBLM_R_X11Y147_SLICE_X14Y147_CO6),
.I2(CLBLM_R_X7Y147_SLICE_X9Y147_CQ),
.I3(CLBLM_R_X7Y147_SLICE_X9Y147_BQ),
.I4(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.I5(CLBLM_L_X8Y147_SLICE_X10Y147_BQ),
.O5(CLBLM_L_X8Y147_SLICE_X11Y147_CO5),
.O6(CLBLM_L_X8Y147_SLICE_X11Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f0f0e4e4)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_BLUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I1(CLBLM_L_X8Y147_SLICE_X11Y147_BQ),
.I2(CLBLM_L_X8Y148_SLICE_X11Y148_AQ),
.I3(CLBLM_L_X10Y146_SLICE_X12Y146_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y147_SLICE_X11Y147_BO5),
.O6(CLBLM_L_X8Y147_SLICE_X11Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ccffccf0)
  ) CLBLM_L_X8Y147_SLICE_X11Y147_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y148_SLICE_X6Y148_BQ),
.I2(CLBLM_L_X8Y147_SLICE_X11Y147_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y146_SLICE_X15Y146_AQ),
.I5(CLBLM_R_X7Y146_SLICE_X9Y146_DO6),
.O5(CLBLM_L_X8Y147_SLICE_X11Y147_AO5),
.O6(CLBLM_L_X8Y147_SLICE_X11Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y148_SLICE_X10Y148_AO6),
.Q(CLBLM_L_X8Y148_SLICE_X10Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y148_SLICE_X10Y148_BO6),
.Q(CLBLM_L_X8Y148_SLICE_X10Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y148_SLICE_X10Y148_CO6),
.Q(CLBLM_L_X8Y148_SLICE_X10Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffbf)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_DLUT (
.I0(CLBLM_L_X8Y148_SLICE_X11Y148_AQ),
.I1(CLBLM_L_X8Y147_SLICE_X10Y147_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y151_SLICE_X9Y151_CQ),
.I4(CLBLM_R_X7Y145_SLICE_X8Y145_AQ),
.I5(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.O5(CLBLM_L_X8Y148_SLICE_X10Y148_DO5),
.O6(CLBLM_L_X8Y148_SLICE_X10Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0ffccfff0ff88)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_CLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X8Y148_SLICE_X10Y148_CQ),
.I2(CLBLM_L_X8Y146_SLICE_X10Y146_B5Q),
.I3(CLBLM_L_X8Y152_SLICE_X11Y152_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.O5(CLBLM_L_X8Y148_SLICE_X10Y148_CO5),
.O6(CLBLM_L_X8Y148_SLICE_X10Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff05ff0400050004)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_BLUT (
.I0(CLBLM_L_X8Y149_SLICE_X10Y149_BO5),
.I1(CLBLM_L_X8Y148_SLICE_X10Y148_BQ),
.I2(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y148_SLICE_X11Y148_CO6),
.I5(CLBLM_L_X10Y151_SLICE_X12Y151_CQ),
.O5(CLBLM_L_X8Y148_SLICE_X10Y148_BO5),
.O6(CLBLM_L_X8Y148_SLICE_X10Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00e2e2ff00aaaa)
  ) CLBLM_L_X8Y148_SLICE_X10Y148_ALUT (
.I0(CLBLM_R_X11Y149_SLICE_X14Y149_DQ),
.I1(CLBLL_L_X4Y151_SLICE_X4Y151_BQ),
.I2(CLBLM_L_X8Y148_SLICE_X10Y148_AQ),
.I3(CLBLM_L_X12Y152_SLICE_X16Y152_B5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y151_SLICE_X12Y151_CQ),
.O5(CLBLM_L_X8Y148_SLICE_X10Y148_AO5),
.O6(CLBLM_L_X8Y148_SLICE_X10Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y148_SLICE_X12Y148_BO6),
.Q(CLBLM_L_X8Y148_SLICE_X11Y148_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y148_SLICE_X11Y148_BO5),
.Q(CLBLM_L_X8Y148_SLICE_X11Y148_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y148_SLICE_X11Y148_AO6),
.Q(CLBLM_L_X8Y148_SLICE_X11Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y148_SLICE_X11Y148_BO6),
.Q(CLBLM_L_X8Y148_SLICE_X11Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00220022dcdc1010)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y151_SLICE_X8Y151_BQ),
.I3(CLBLM_R_X11Y154_SLICE_X14Y154_DQ),
.I4(CLBLM_L_X8Y149_SLICE_X11Y149_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y148_SLICE_X11Y148_DO5),
.O6(CLBLM_L_X8Y148_SLICE_X11Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000000000ffffff)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_L_X10Y148_SLICE_X13Y148_DO6),
.I3(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.I4(CLBLM_R_X11Y149_SLICE_X14Y149_DQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y148_SLICE_X11Y148_CO5),
.O6(CLBLM_L_X8Y148_SLICE_X11Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888e4e4e4e4)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y148_SLICE_X11Y148_A5Q),
.I2(CLBLM_R_X7Y148_SLICE_X9Y148_AQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y151_SLICE_X5Y151_CQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y148_SLICE_X11Y148_BO5),
.O6(CLBLM_L_X8Y148_SLICE_X11Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaeeea00004440)
  ) CLBLM_L_X8Y148_SLICE_X11Y148_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I2(CLBLM_L_X8Y148_SLICE_X11Y148_AQ),
.I3(CLBLM_L_X10Y147_SLICE_X12Y147_BQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLL_L_X4Y150_SLICE_X5Y150_DQ),
.O5(CLBLM_L_X8Y148_SLICE_X11Y148_AO5),
.O6(CLBLM_L_X8Y148_SLICE_X11Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y149_SLICE_X10Y149_AO6),
.Q(CLBLM_L_X8Y149_SLICE_X10Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h80007fff0000ffff)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_DLUT (
.I0(CLBLM_L_X10Y148_SLICE_X13Y148_DO6),
.I1(CLBLM_R_X11Y149_SLICE_X14Y149_DQ),
.I2(CLBLM_L_X8Y149_SLICE_X10Y149_AQ),
.I3(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.I4(CLBLM_L_X8Y155_SLICE_X10Y155_B5Q),
.I5(CLBLM_L_X8Y148_SLICE_X10Y148_BQ),
.O5(CLBLM_L_X8Y149_SLICE_X10Y149_DO5),
.O6(CLBLM_L_X8Y149_SLICE_X10Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffffffffffff)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_CLUT (
.I0(CLBLM_L_X10Y150_SLICE_X13Y150_BQ),
.I1(CLBLM_L_X10Y148_SLICE_X13Y148_BQ),
.I2(CLBLM_L_X8Y155_SLICE_X10Y155_B5Q),
.I3(CLBLM_R_X7Y149_SLICE_X9Y149_C5Q),
.I4(CLBLM_L_X10Y148_SLICE_X13Y148_AQ),
.I5(CLBLM_L_X10Y155_SLICE_X12Y155_BQ),
.O5(CLBLM_L_X8Y149_SLICE_X10Y149_CO5),
.O6(CLBLM_L_X8Y149_SLICE_X10Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffff88000000)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_BLUT (
.I0(CLBLM_R_X11Y149_SLICE_X14Y149_DQ),
.I1(CLBLM_L_X8Y148_SLICE_X10Y148_BQ),
.I2(CLBLM_L_X8Y149_SLICE_X10Y149_AQ),
.I3(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.I4(CLBLM_L_X10Y148_SLICE_X13Y148_DO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y149_SLICE_X10Y149_BO5),
.O6(CLBLM_L_X8Y149_SLICE_X10Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfecc00003200)
  ) CLBLM_L_X8Y149_SLICE_X10Y149_ALUT (
.I0(CLBLM_L_X8Y149_SLICE_X10Y149_BO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y149_SLICE_X10Y149_AQ),
.I3(CLBLM_L_X8Y149_SLICE_X10Y149_BO6),
.I4(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I5(CLBLM_L_X10Y155_SLICE_X12Y155_BQ),
.O5(CLBLM_L_X8Y149_SLICE_X10Y149_AO5),
.O6(CLBLM_L_X8Y149_SLICE_X10Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y149_SLICE_X11Y149_AO6),
.Q(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y149_SLICE_X11Y149_BO6),
.Q(CLBLM_L_X8Y149_SLICE_X11Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y149_SLICE_X11Y149_CO6),
.Q(CLBLM_L_X8Y149_SLICE_X11Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555ffffffff)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_DLUT (
.I0(CLBLM_L_X10Y148_SLICE_X13Y148_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y155_SLICE_X12Y155_BQ),
.O5(CLBLM_L_X8Y149_SLICE_X11Y149_DO5),
.O6(CLBLM_L_X8Y149_SLICE_X11Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haf05aa00ae04aa00)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y149_SLICE_X11Y149_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_R_X7Y147_SLICE_X9Y147_A5Q),
.I4(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I5(CLBLM_L_X10Y147_SLICE_X13Y147_AQ),
.O5(CLBLM_L_X8Y149_SLICE_X11Y149_CO5),
.O6(CLBLM_L_X8Y149_SLICE_X11Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf808fc0cf808fc0c)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_BLUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I1(CLBLM_L_X8Y149_SLICE_X11Y149_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y150_SLICE_X5Y150_CQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y149_SLICE_X11Y149_BO5),
.O6(CLBLM_L_X8Y149_SLICE_X11Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffccccf0a0)
  ) CLBLM_L_X8Y149_SLICE_X11Y149_ALUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I1(CLBLM_R_X5Y151_SLICE_X6Y151_CQ),
.I2(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y150_SLICE_X9Y150_CO6),
.O5(CLBLM_L_X8Y149_SLICE_X11Y149_AO5),
.O6(CLBLM_L_X8Y149_SLICE_X11Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y150_SLICE_X10Y150_CO6),
.Q(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y150_SLICE_X10Y150_AO6),
.Q(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y150_SLICE_X10Y150_BO6),
.Q(CLBLM_L_X8Y150_SLICE_X10Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaaaccccaa55)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_DLUT (
.I0(CLBLM_L_X10Y148_SLICE_X12Y148_AQ),
.I1(CLBLM_R_X5Y151_SLICE_X6Y151_CQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y147_SLICE_X10Y147_CQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_L_X10Y150_SLICE_X12Y150_BO5),
.O5(CLBLM_L_X8Y150_SLICE_X10Y150_DO5),
.O6(CLBLM_L_X8Y150_SLICE_X10Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heaea4040ff000000)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y151_SLICE_X13Y151_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X8Y148_SLICE_X10Y148_BQ),
.I4(CLBLM_L_X8Y149_SLICE_X10Y149_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y150_SLICE_X10Y150_CO5),
.O6(CLBLM_L_X8Y150_SLICE_X10Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f808f808)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y150_SLICE_X10Y150_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y151_SLICE_X10Y151_BQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y151_SLICE_X9Y151_CQ),
.O5(CLBLM_L_X8Y150_SLICE_X10Y150_BO5),
.O6(CLBLM_L_X8Y150_SLICE_X10Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f1f0f000010000)
  ) CLBLM_L_X8Y150_SLICE_X10Y150_ALUT (
.I0(CLBLM_L_X8Y148_SLICE_X11Y148_CO5),
.I1(CLBLM_R_X11Y152_SLICE_X15Y152_DQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y149_SLICE_X10Y149_CO6),
.I4(CLBLM_L_X8Y150_SLICE_X10Y150_CO5),
.I5(CLBLM_R_X7Y156_SLICE_X9Y156_CQ),
.O5(CLBLM_L_X8Y150_SLICE_X10Y150_AO5),
.O6(CLBLM_L_X8Y150_SLICE_X10Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y150_SLICE_X11Y150_AO6),
.Q(CLBLM_L_X8Y150_SLICE_X11Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y150_SLICE_X11Y150_BO6),
.Q(CLBLM_L_X8Y150_SLICE_X11Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y150_SLICE_X11Y150_CO6),
.Q(CLBLM_L_X8Y150_SLICE_X11Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2020002033330033)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_DLUT (
.I0(CLBLM_L_X10Y148_SLICE_X13Y148_AQ),
.I1(CLBLM_L_X10Y150_SLICE_X13Y150_BQ),
.I2(CLBLM_R_X11Y152_SLICE_X15Y152_DQ),
.I3(CLBLM_L_X8Y148_SLICE_X11Y148_CO5),
.I4(CLBLM_L_X8Y150_SLICE_X10Y150_CO5),
.I5(CLBLM_L_X8Y149_SLICE_X11Y149_DO6),
.O5(CLBLM_L_X8Y150_SLICE_X11Y150_DO5),
.O6(CLBLM_L_X8Y150_SLICE_X11Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff0fff000f044)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_CLUT (
.I0(CLBLM_R_X7Y148_SLICE_X9Y148_CO6),
.I1(CLBLM_R_X7Y158_SLICE_X8Y158_CO5),
.I2(CLBLM_L_X8Y146_SLICE_X11Y146_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y150_SLICE_X11Y150_DO6),
.I5(CLBLM_L_X8Y156_SLICE_X11Y156_CO6),
.O5(CLBLM_L_X8Y150_SLICE_X11Y150_CO5),
.O6(CLBLM_L_X8Y150_SLICE_X11Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaffccf0c0)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_BLUT (
.I0(CLBLM_L_X8Y157_SLICE_X10Y157_BQ),
.I1(CLBLM_L_X8Y150_SLICE_X11Y150_BQ),
.I2(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I3(CLBLM_L_X8Y151_SLICE_X11Y151_BO6),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y150_SLICE_X11Y150_BO5),
.O6(CLBLM_L_X8Y150_SLICE_X11Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c5c0c5c5c0c5c0)
  ) CLBLM_L_X8Y150_SLICE_X11Y150_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y146_SLICE_X11Y146_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y152_SLICE_X7Y152_CQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y152_SLICE_X14Y152_DO6),
.O5(CLBLM_L_X8Y150_SLICE_X11Y150_AO5),
.O6(CLBLM_L_X8Y150_SLICE_X11Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y151_SLICE_X10Y151_AO6),
.Q(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y151_SLICE_X10Y151_BO6),
.Q(CLBLM_L_X8Y151_SLICE_X10Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y151_SLICE_X10Y151_CO6),
.Q(CLBLM_L_X8Y151_SLICE_X10Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699669999669966)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_DLUT (
.I0(CLBLM_L_X10Y157_SLICE_X12Y157_AQ),
.I1(CLBLM_L_X8Y151_SLICE_X10Y151_CQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y152_SLICE_X8Y152_A5Q),
.I4(1'b1),
.I5(CLBLM_L_X10Y150_SLICE_X12Y150_CQ),
.O5(CLBLM_L_X8Y151_SLICE_X10Y151_DO5),
.O6(CLBLM_L_X8Y151_SLICE_X10Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00f0f000)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_CLUT (
.I0(CLBLM_R_X7Y153_SLICE_X8Y153_BQ),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y149_SLICE_X13Y149_CO6),
.I4(CLBLM_L_X8Y151_SLICE_X10Y151_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y151_SLICE_X10Y151_CO5),
.O6(CLBLM_L_X8Y151_SLICE_X10Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff440044ff440044)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y151_SLICE_X10Y151_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y151_SLICE_X11Y151_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y151_SLICE_X10Y151_BO5),
.O6(CLBLM_L_X8Y151_SLICE_X10Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfaccfaccfacc00)
  ) CLBLM_L_X8Y151_SLICE_X10Y151_ALUT (
.I0(CLBLM_L_X8Y151_SLICE_X11Y151_CO6),
.I1(CLBLM_L_X12Y154_SLICE_X17Y154_BQ),
.I2(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X8Y151_SLICE_X10Y151_AO5),
.O6(CLBLM_L_X8Y151_SLICE_X10Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y151_SLICE_X11Y151_AO6),
.Q(CLBLM_L_X8Y151_SLICE_X11Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ff00ff00)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X8Y152_SLICE_X10Y152_BQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y150_SLICE_X10Y150_BQ),
.O5(CLBLM_L_X8Y151_SLICE_X11Y151_DO5),
.O6(CLBLM_L_X8Y151_SLICE_X11Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc5cfcfc0cac0c0)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_CLUT (
.I0(CLBLM_R_X7Y151_SLICE_X8Y151_CQ),
.I1(CLBLM_L_X10Y151_SLICE_X13Y151_BQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X8Y147_SLICE_X10Y147_CQ),
.I4(CLBLM_L_X8Y151_SLICE_X11Y151_DO6),
.I5(CLBLM_L_X8Y151_SLICE_X10Y151_BQ),
.O5(CLBLM_L_X8Y151_SLICE_X11Y151_CO5),
.O6(CLBLM_L_X8Y151_SLICE_X11Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff78fff0007800f0)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_BLUT (
.I0(CLBLM_L_X8Y152_SLICE_X11Y152_BO6),
.I1(CLBLM_L_X8Y150_SLICE_X10Y150_BQ),
.I2(CLBLM_R_X5Y150_SLICE_X7Y150_AQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X8Y152_SLICE_X10Y152_BQ),
.I5(CLBLM_R_X7Y151_SLICE_X8Y151_DQ),
.O5(CLBLM_L_X8Y151_SLICE_X11Y151_BO5),
.O6(CLBLM_L_X8Y151_SLICE_X11Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f40104f1f40104)
  ) CLBLM_L_X8Y151_SLICE_X11Y151_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y152_SLICE_X9Y152_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y151_SLICE_X11Y151_BO6),
.I4(CLBLM_R_X13Y150_SLICE_X19Y150_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y151_SLICE_X11Y151_AO5),
.O6(CLBLM_L_X8Y151_SLICE_X11Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y152_SLICE_X10Y152_AO6),
.Q(CLBLM_L_X8Y152_SLICE_X10Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y152_SLICE_X10Y152_BO6),
.Q(CLBLM_L_X8Y152_SLICE_X10Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y152_SLICE_X10Y152_CO6),
.Q(CLBLM_L_X8Y152_SLICE_X10Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccd8881cccc8888)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_DLUT (
.I0(CLBLM_R_X5Y151_SLICE_X7Y151_CQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X8Y152_SLICE_X11Y152_BO5),
.I3(CLBLM_L_X8Y152_SLICE_X10Y152_BQ),
.I4(CLBLM_R_X11Y151_SLICE_X15Y151_AQ),
.I5(CLBLM_L_X8Y150_SLICE_X10Y150_BQ),
.O5(CLBLM_L_X8Y152_SLICE_X10Y152_DO5),
.O6(CLBLM_L_X8Y152_SLICE_X10Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0aaaaccaa)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_CLUT (
.I0(CLBLM_L_X10Y148_SLICE_X13Y148_BQ),
.I1(CLBLM_L_X8Y152_SLICE_X10Y152_CQ),
.I2(CLBLM_R_X13Y153_SLICE_X19Y153_AQ),
.I3(CLBLM_L_X10Y150_SLICE_X12Y150_A5Q),
.I4(CLBLM_L_X12Y155_SLICE_X16Y155_CO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y152_SLICE_X10Y152_CO5),
.O6(CLBLM_L_X8Y152_SLICE_X10Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f088f088)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X8Y152_SLICE_X10Y152_BQ),
.I2(CLBLM_L_X8Y153_SLICE_X10Y153_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y151_SLICE_X9Y151_CQ),
.O5(CLBLM_L_X8Y152_SLICE_X10Y152_BO5),
.O6(CLBLM_L_X8Y152_SLICE_X10Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfaccfaccfacc00)
  ) CLBLM_L_X8Y152_SLICE_X10Y152_ALUT (
.I0(CLBLM_L_X8Y152_SLICE_X10Y152_DO6),
.I1(CLBLL_L_X4Y146_SLICE_X5Y146_AQ),
.I2(CLBLM_L_X8Y152_SLICE_X10Y152_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.O5(CLBLM_L_X8Y152_SLICE_X10Y152_AO5),
.O6(CLBLM_L_X8Y152_SLICE_X10Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc33cc33cc639c)
  ) CLBLM_L_X8Y152_SLICE_X11Y152_DLUT (
.I0(CLBLM_L_X8Y147_SLICE_X10Y147_CQ),
.I1(CLBLM_L_X10Y151_SLICE_X12Y151_CQ),
.I2(CLBLM_L_X8Y152_SLICE_X10Y152_BQ),
.I3(CLBLM_L_X8Y155_SLICE_X11Y155_DO6),
.I4(CLBLM_R_X7Y151_SLICE_X8Y151_CQ),
.I5(CLBLM_L_X8Y150_SLICE_X10Y150_BQ),
.O5(CLBLM_L_X8Y152_SLICE_X11Y152_DO5),
.O6(CLBLM_L_X8Y152_SLICE_X11Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff8aaa00000000)
  ) CLBLM_L_X8Y152_SLICE_X11Y152_CLUT (
.I0(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.I1(CLBLL_L_X4Y153_SLICE_X4Y153_BO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X8Y152_SLICE_X11Y152_AO5),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I5(CLBLM_L_X10Y149_SLICE_X13Y149_BO5),
.O5(CLBLM_L_X8Y152_SLICE_X11Y152_CO5),
.O6(CLBLM_L_X8Y152_SLICE_X11Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f000ff0fff0ff)
  ) CLBLM_L_X8Y152_SLICE_X11Y152_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X7Y151_SLICE_X8Y151_CQ),
.I3(CLBLM_L_X8Y147_SLICE_X10Y147_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y152_SLICE_X11Y152_BO5),
.O6(CLBLM_L_X8Y152_SLICE_X11Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a5a50f555555ff)
  ) CLBLM_L_X8Y152_SLICE_X11Y152_ALUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(1'b1),
.I2(CLBLM_L_X8Y150_SLICE_X11Y150_AQ),
.I3(CLBLM_R_X5Y151_SLICE_X6Y151_CQ),
.I4(CLBLM_L_X8Y152_SLICE_X10Y152_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y152_SLICE_X11Y152_AO5),
.O6(CLBLM_L_X8Y152_SLICE_X11Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y153_SLICE_X10Y153_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y153_SLICE_X10Y153_AO5),
.Q(CLBLM_L_X8Y153_SLICE_X10Y153_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y153_SLICE_X10Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y153_SLICE_X10Y153_AO6),
.Q(CLBLM_L_X8Y153_SLICE_X10Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbf3fffffffffffff)
  ) CLBLM_L_X8Y153_SLICE_X10Y153_DLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X10Y153_SLICE_X12Y153_CO6),
.I2(CLBLM_R_X7Y153_SLICE_X9Y153_CO6),
.I3(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I4(CLBLM_L_X8Y155_SLICE_X11Y155_DO6),
.I5(CLBLM_R_X5Y151_SLICE_X7Y151_BQ),
.O5(CLBLM_L_X8Y153_SLICE_X10Y153_DO5),
.O6(CLBLM_L_X8Y153_SLICE_X10Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0f7f000000088)
  ) CLBLM_L_X8Y153_SLICE_X10Y153_CLUT (
.I0(CLBLM_L_X8Y152_SLICE_X10Y152_BQ),
.I1(CLBLM_L_X8Y150_SLICE_X10Y150_BQ),
.I2(CLBLM_R_X5Y152_SLICE_X6Y152_BQ),
.I3(CLBLM_R_X7Y157_SLICE_X9Y157_DQ),
.I4(CLBLM_L_X8Y152_SLICE_X11Y152_BO5),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_L_X8Y153_SLICE_X10Y153_CO5),
.O6(CLBLM_L_X8Y153_SLICE_X10Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccefcc00000050)
  ) CLBLM_L_X8Y153_SLICE_X10Y153_BLUT (
.I0(CLBLM_L_X8Y152_SLICE_X11Y152_BO5),
.I1(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I2(CLBLM_L_X8Y152_SLICE_X10Y152_BQ),
.I3(CLBLM_L_X8Y158_SLICE_X10Y158_BQ),
.I4(CLBLM_L_X8Y150_SLICE_X10Y150_BQ),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_L_X8Y153_SLICE_X10Y153_BO5),
.O6(CLBLM_L_X8Y153_SLICE_X10Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00ccf0f0aaaa)
  ) CLBLM_L_X8Y153_SLICE_X10Y153_ALUT (
.I0(CLBLM_L_X8Y154_SLICE_X10Y154_CQ),
.I1(CLBLM_L_X8Y157_SLICE_X10Y157_DQ),
.I2(CLBLM_L_X10Y151_SLICE_X13Y151_BQ),
.I3(CLBLM_R_X11Y159_SLICE_X15Y159_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y153_SLICE_X10Y153_AO5),
.O6(CLBLM_L_X8Y153_SLICE_X10Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y153_SLICE_X11Y153_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y153_SLICE_X11Y153_CO5),
.Q(CLBLM_L_X8Y153_SLICE_X11Y153_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y153_SLICE_X11Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y153_SLICE_X11Y153_AO6),
.Q(CLBLM_L_X8Y153_SLICE_X11Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y153_SLICE_X11Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y153_SLICE_X11Y153_BO6),
.Q(CLBLM_L_X8Y153_SLICE_X11Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y153_SLICE_X11Y153_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y153_SLICE_X11Y153_CO6),
.Q(CLBLM_L_X8Y153_SLICE_X11Y153_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y153_SLICE_X11Y153_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y153_SLICE_X11Y153_DO6),
.Q(CLBLM_L_X8Y153_SLICE_X11Y153_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc005a005a)
  ) CLBLM_L_X8Y153_SLICE_X11Y153_DLUT (
.I0(CLBLM_L_X10Y152_SLICE_X13Y152_BO5),
.I1(CLBLM_L_X8Y153_SLICE_X10Y153_A5Q),
.I2(CLBLM_R_X5Y152_SLICE_X6Y152_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y153_SLICE_X11Y153_DO5),
.O6(CLBLM_L_X8Y153_SLICE_X11Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0e4a0e4dddd8888)
  ) CLBLM_L_X8Y153_SLICE_X11Y153_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y154_SLICE_X12Y154_DQ),
.I2(CLBLM_L_X8Y153_SLICE_X11Y153_DQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X7Y148_SLICE_X8Y148_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y153_SLICE_X11Y153_CO5),
.O6(CLBLM_L_X8Y153_SLICE_X11Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcccc00330000)
  ) CLBLM_L_X8Y153_SLICE_X11Y153_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_R_X11Y159_SLICE_X15Y159_CO6),
.I4(CLBLM_L_X8Y153_SLICE_X10Y153_AQ),
.I5(CLBLM_L_X10Y153_SLICE_X13Y153_DQ),
.O5(CLBLM_L_X8Y153_SLICE_X11Y153_BO5),
.O6(CLBLM_L_X8Y153_SLICE_X11Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33ee22cf03fc30)
  ) CLBLM_L_X8Y153_SLICE_X11Y153_ALUT (
.I0(CLBLM_L_X10Y153_SLICE_X13Y153_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y153_SLICE_X11Y153_AQ),
.I3(CLBLL_L_X4Y148_SLICE_X5Y148_DQ),
.I4(CLBLM_R_X13Y150_SLICE_X18Y150_BQ),
.I5(CLBLM_R_X7Y153_SLICE_X9Y153_CO6),
.O5(CLBLM_L_X8Y153_SLICE_X11Y153_AO5),
.O6(CLBLM_L_X8Y153_SLICE_X11Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y154_SLICE_X10Y154_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y154_SLICE_X10Y154_AO5),
.Q(CLBLM_L_X8Y154_SLICE_X10Y154_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y154_SLICE_X10Y154_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y154_SLICE_X10Y154_BO5),
.Q(CLBLM_L_X8Y154_SLICE_X10Y154_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y154_SLICE_X10Y154_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y154_SLICE_X10Y154_CO5),
.Q(CLBLM_L_X8Y154_SLICE_X10Y154_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y154_SLICE_X10Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y154_SLICE_X10Y154_AO6),
.Q(CLBLM_L_X8Y154_SLICE_X10Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y154_SLICE_X10Y154_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y154_SLICE_X10Y154_BO6),
.Q(CLBLM_L_X8Y154_SLICE_X10Y154_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y154_SLICE_X10Y154_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y154_SLICE_X10Y154_CO6),
.Q(CLBLM_L_X8Y154_SLICE_X10Y154_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y154_SLICE_X10Y154_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y154_SLICE_X10Y154_DO6),
.Q(CLBLM_L_X8Y154_SLICE_X10Y154_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefeaafe54540054)
  ) CLBLM_L_X8Y154_SLICE_X10Y154_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y149_SLICE_X14Y149_DQ),
.I2(CLBLM_L_X8Y154_SLICE_X10Y154_DQ),
.I3(CLBLM_L_X10Y150_SLICE_X12Y150_A5Q),
.I4(CLBLM_L_X12Y155_SLICE_X16Y155_CO6),
.I5(CLBLM_L_X8Y158_SLICE_X10Y158_BQ),
.O5(CLBLM_L_X8Y154_SLICE_X10Y154_DO5),
.O6(CLBLM_L_X8Y154_SLICE_X10Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0a0fc0cfc0c)
  ) CLBLM_L_X8Y154_SLICE_X10Y154_CLUT (
.I0(CLBLM_L_X8Y157_SLICE_X11Y157_AQ),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I4(CLBLM_L_X8Y154_SLICE_X10Y154_B5Q),
.I5(1'b1),
.O5(CLBLM_L_X8Y154_SLICE_X10Y154_CO5),
.O6(CLBLM_L_X8Y154_SLICE_X10Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaf0fff000f0)
  ) CLBLM_L_X8Y154_SLICE_X10Y154_BLUT (
.I0(CLBLM_R_X3Y150_SLICE_X2Y150_A5Q),
.I1(1'b1),
.I2(RIOB33_X105Y143_IOB_X1Y144_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y158_SLICE_X12Y158_BQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y154_SLICE_X10Y154_BO5),
.O6(CLBLM_L_X8Y154_SLICE_X10Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff000f0eeaaeeaa)
  ) CLBLM_L_X8Y154_SLICE_X10Y154_ALUT (
.I0(CLBLM_R_X7Y156_SLICE_X9Y156_DO6),
.I1(CLBLL_L_X4Y152_SLICE_X5Y152_CQ),
.I2(CLBLM_L_X12Y156_SLICE_X16Y156_CO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y147_SLICE_X11Y147_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y154_SLICE_X10Y154_AO5),
.O6(CLBLM_L_X8Y154_SLICE_X10Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y154_SLICE_X11Y154_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y154_SLICE_X14Y154_BO6),
.Q(CLBLM_L_X8Y154_SLICE_X11Y154_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y154_SLICE_X11Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y154_SLICE_X11Y154_AO6),
.Q(CLBLM_L_X8Y154_SLICE_X11Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y154_SLICE_X11Y154_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y154_SLICE_X11Y154_BO6),
.Q(CLBLM_L_X8Y154_SLICE_X11Y154_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y154_SLICE_X11Y154_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y154_SLICE_X11Y154_CO6),
.Q(CLBLM_L_X8Y154_SLICE_X11Y154_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeeeeffffeeee)
  ) CLBLM_L_X8Y154_SLICE_X11Y154_DLUT (
.I0(CLBLM_R_X5Y151_SLICE_X7Y151_CQ),
.I1(CLBLM_R_X7Y157_SLICE_X9Y157_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X5Y150_SLICE_X7Y150_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y154_SLICE_X11Y154_DO5),
.O6(CLBLM_L_X8Y154_SLICE_X11Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaffccf0c0)
  ) CLBLM_L_X8Y154_SLICE_X11Y154_CLUT (
.I0(CLBLM_L_X10Y157_SLICE_X12Y157_AQ),
.I1(CLBLM_L_X8Y154_SLICE_X11Y154_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X8Y153_SLICE_X10Y153_CO6),
.I4(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y154_SLICE_X11Y154_CO5),
.O6(CLBLM_L_X8Y154_SLICE_X11Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaf0aac0aac0)
  ) CLBLM_L_X8Y154_SLICE_X11Y154_BLUT (
.I0(CLBLM_L_X8Y155_SLICE_X10Y155_BQ),
.I1(CLBLM_L_X8Y154_SLICE_X11Y154_BQ),
.I2(CLBLM_R_X7Y153_SLICE_X9Y153_CO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X10Y154_SLICE_X12Y154_DQ),
.O5(CLBLM_L_X8Y154_SLICE_X11Y154_BO5),
.O6(CLBLM_L_X8Y154_SLICE_X11Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00e4e4e4e4)
  ) CLBLM_L_X8Y154_SLICE_X11Y154_ALUT (
.I0(CLBLM_R_X7Y153_SLICE_X9Y153_CO6),
.I1(CLBLM_L_X10Y156_SLICE_X13Y156_BQ),
.I2(CLBLM_L_X8Y154_SLICE_X11Y154_AQ),
.I3(CLBLM_R_X7Y154_SLICE_X8Y154_CQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y154_SLICE_X11Y154_AO5),
.O6(CLBLM_L_X8Y154_SLICE_X11Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y155_SLICE_X10Y155_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y155_SLICE_X10Y155_BO5),
.Q(CLBLM_L_X8Y155_SLICE_X10Y155_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y155_SLICE_X10Y155_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y155_SLICE_X10Y155_AO6),
.Q(CLBLM_L_X8Y155_SLICE_X10Y155_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y155_SLICE_X10Y155_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y155_SLICE_X10Y155_BO6),
.Q(CLBLM_L_X8Y155_SLICE_X10Y155_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y155_SLICE_X10Y155_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y155_SLICE_X10Y155_CO6),
.Q(CLBLM_L_X8Y155_SLICE_X10Y155_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0020000000000000)
  ) CLBLM_L_X8Y155_SLICE_X10Y155_DLUT (
.I0(CLBLM_L_X8Y152_SLICE_X10Y152_CQ),
.I1(CLBLM_L_X8Y153_SLICE_X10Y153_DO6),
.I2(CLBLM_L_X8Y149_SLICE_X10Y149_DO6),
.I3(CLBLL_L_X4Y156_SLICE_X4Y156_CO5),
.I4(CLBLM_R_X7Y155_SLICE_X9Y155_CO6),
.I5(CLBLM_R_X13Y152_SLICE_X19Y152_CO6),
.O5(CLBLM_L_X8Y155_SLICE_X10Y155_DO5),
.O6(CLBLM_L_X8Y155_SLICE_X10Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff5c40000f5c4)
  ) CLBLM_L_X8Y155_SLICE_X10Y155_CLUT (
.I0(CLBLM_L_X10Y150_SLICE_X12Y150_A5Q),
.I1(CLBLM_L_X8Y155_SLICE_X10Y155_CQ),
.I2(CLBLM_L_X12Y155_SLICE_X16Y155_CO6),
.I3(CLBLM_L_X10Y155_SLICE_X12Y155_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y155_SLICE_X10Y155_AQ),
.O5(CLBLM_L_X8Y155_SLICE_X10Y155_CO5),
.O6(CLBLM_L_X8Y155_SLICE_X10Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f0f0cccc0055)
  ) CLBLM_L_X8Y155_SLICE_X10Y155_BLUT (
.I0(CLBLM_L_X8Y149_SLICE_X10Y149_DO6),
.I1(CLBLM_R_X5Y155_SLICE_X6Y155_AQ),
.I2(CLBLM_L_X8Y154_SLICE_X11Y154_A5Q),
.I3(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y155_SLICE_X10Y155_BO5),
.O6(CLBLM_L_X8Y155_SLICE_X10Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ff00f0f0cccc)
  ) CLBLM_L_X8Y155_SLICE_X10Y155_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y155_SLICE_X12Y155_CQ),
.I2(CLBLM_R_X5Y152_SLICE_X6Y152_BQ),
.I3(CLBLM_L_X8Y155_SLICE_X10Y155_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y153_SLICE_X9Y153_CO6),
.O5(CLBLM_L_X8Y155_SLICE_X10Y155_AO5),
.O6(CLBLM_L_X8Y155_SLICE_X10Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y155_SLICE_X11Y155_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y155_SLICE_X11Y155_AO6),
.Q(CLBLM_L_X8Y155_SLICE_X11Y155_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y155_SLICE_X11Y155_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y155_SLICE_X11Y155_BO6),
.Q(CLBLM_L_X8Y155_SLICE_X11Y155_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y155_SLICE_X11Y155_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y155_SLICE_X11Y155_CO6),
.Q(CLBLM_L_X8Y155_SLICE_X11Y155_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc33cc33cc33cf)
  ) CLBLM_L_X8Y155_SLICE_X11Y155_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y157_SLICE_X11Y157_CQ),
.I2(CLBLM_L_X10Y155_SLICE_X12Y155_DO6),
.I3(CLBLM_L_X8Y156_SLICE_X11Y156_BQ),
.I4(CLBLM_L_X8Y154_SLICE_X11Y154_DO6),
.I5(CLBLM_L_X10Y150_SLICE_X12Y150_DO6),
.O5(CLBLM_L_X8Y155_SLICE_X11Y155_DO5),
.O6(CLBLM_L_X8Y155_SLICE_X11Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000030303030)
  ) CLBLM_L_X8Y155_SLICE_X11Y155_CLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y156_SLICE_X10Y156_CQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y154_SLICE_X9Y154_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y155_SLICE_X11Y155_CO5),
.O6(CLBLM_L_X8Y155_SLICE_X11Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000ddee1122)
  ) CLBLM_L_X8Y155_SLICE_X11Y155_BLUT (
.I0(CLBLM_L_X10Y153_SLICE_X13Y153_DQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_L_X12Y153_SLICE_X17Y153_DO5),
.I4(CLBLM_R_X5Y155_SLICE_X7Y155_BQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y155_SLICE_X11Y155_BO5),
.O6(CLBLM_L_X8Y155_SLICE_X11Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haafcaafcaa00aa00)
  ) CLBLM_L_X8Y155_SLICE_X11Y155_ALUT (
.I0(CLBLM_R_X7Y151_SLICE_X8Y151_CQ),
.I1(CLBLM_R_X13Y155_SLICE_X18Y155_BQ),
.I2(CLBLM_L_X8Y155_SLICE_X11Y155_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y153_SLICE_X9Y153_CO6),
.O5(CLBLM_L_X8Y155_SLICE_X11Y155_AO5),
.O6(CLBLM_L_X8Y155_SLICE_X11Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y156_SLICE_X10Y156_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y156_SLICE_X10Y156_AO6),
.Q(CLBLM_L_X8Y156_SLICE_X10Y156_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y156_SLICE_X10Y156_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y156_SLICE_X10Y156_BO6),
.Q(CLBLM_L_X8Y156_SLICE_X10Y156_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y156_SLICE_X10Y156_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y156_SLICE_X10Y156_CO6),
.Q(CLBLM_L_X8Y156_SLICE_X10Y156_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aa55aa55aa)
  ) CLBLM_L_X8Y156_SLICE_X10Y156_DLUT (
.I0(CLBLM_L_X8Y155_SLICE_X11Y155_BQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X12Y158_SLICE_X16Y158_A5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y156_SLICE_X10Y156_DO5),
.O6(CLBLM_L_X8Y156_SLICE_X10Y156_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa03c0003c)
  ) CLBLM_L_X8Y156_SLICE_X10Y156_CLUT (
.I0(CLBLM_L_X8Y154_SLICE_X10Y154_BQ),
.I1(CLBLM_L_X8Y156_SLICE_X10Y156_CQ),
.I2(CLBLM_L_X10Y154_SLICE_X12Y154_DQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X8Y156_SLICE_X10Y156_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y156_SLICE_X10Y156_CO5),
.O6(CLBLM_L_X8Y156_SLICE_X10Y156_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0afacafacafac)
  ) CLBLM_L_X8Y156_SLICE_X10Y156_BLUT (
.I0(CLBLM_L_X12Y157_SLICE_X16Y157_BQ),
.I1(CLBLM_L_X8Y156_SLICE_X10Y156_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y155_SLICE_X10Y155_B5Q),
.I4(CLBLL_L_X4Y151_SLICE_X4Y151_BQ),
.I5(CLBLM_L_X10Y151_SLICE_X12Y151_CQ),
.O5(CLBLM_L_X8Y156_SLICE_X10Y156_BO5),
.O6(CLBLM_L_X8Y156_SLICE_X10Y156_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00fcaaaafcfc)
  ) CLBLM_L_X8Y156_SLICE_X10Y156_ALUT (
.I0(CLBLM_R_X11Y159_SLICE_X14Y159_DQ),
.I1(CLBLM_L_X10Y155_SLICE_X12Y155_BQ),
.I2(CLBLM_L_X8Y156_SLICE_X10Y156_AQ),
.I3(CLBLL_L_X4Y151_SLICE_X4Y151_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y151_SLICE_X12Y151_CQ),
.O5(CLBLM_L_X8Y156_SLICE_X10Y156_AO5),
.O6(CLBLM_L_X8Y156_SLICE_X10Y156_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y156_SLICE_X11Y156_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y156_SLICE_X11Y156_BO5),
.Q(CLBLM_L_X8Y156_SLICE_X11Y156_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y156_SLICE_X11Y156_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y156_SLICE_X11Y156_AO6),
.Q(CLBLM_L_X8Y156_SLICE_X11Y156_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y156_SLICE_X11Y156_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y156_SLICE_X11Y156_BO6),
.Q(CLBLM_L_X8Y156_SLICE_X11Y156_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0f7707ffffffff)
  ) CLBLM_L_X8Y156_SLICE_X11Y156_DLUT (
.I0(CLBLM_L_X8Y158_SLICE_X10Y158_AQ),
.I1(CLBLM_L_X8Y154_SLICE_X10Y154_A5Q),
.I2(CLBLM_L_X8Y150_SLICE_X11Y150_CQ),
.I3(CLBLM_L_X10Y156_SLICE_X13Y156_AO6),
.I4(CLBLM_R_X7Y155_SLICE_X8Y155_AQ),
.I5(CLBLM_R_X7Y155_SLICE_X8Y155_BO5),
.O5(CLBLM_L_X8Y156_SLICE_X11Y156_DO5),
.O6(CLBLM_L_X8Y156_SLICE_X11Y156_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555aaaa5554aa00)
  ) CLBLM_L_X8Y156_SLICE_X11Y156_CLUT (
.I0(CLBLM_R_X7Y155_SLICE_X8Y155_BO5),
.I1(CLBLM_L_X8Y154_SLICE_X10Y154_A5Q),
.I2(CLBLM_L_X8Y158_SLICE_X10Y158_AQ),
.I3(CLBLM_R_X7Y148_SLICE_X8Y148_AQ),
.I4(CLBLM_L_X8Y150_SLICE_X11Y150_CQ),
.I5(CLBLM_R_X7Y148_SLICE_X8Y148_BQ),
.O5(CLBLM_L_X8Y156_SLICE_X11Y156_CO5),
.O6(CLBLM_L_X8Y156_SLICE_X11Y156_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0acaccfc0cfc0)
  ) CLBLM_L_X8Y156_SLICE_X11Y156_BLUT (
.I0(CLBLM_R_X13Y155_SLICE_X18Y155_BQ),
.I1(CLBLM_L_X8Y156_SLICE_X11Y156_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y154_SLICE_X4Y154_BO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y156_SLICE_X11Y156_BO5),
.O6(CLBLM_L_X8Y156_SLICE_X11Y156_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88dd8888d8ddd888)
  ) CLBLM_L_X8Y156_SLICE_X11Y156_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y153_SLICE_X11Y153_C5Q),
.I2(CLBLM_L_X8Y156_SLICE_X11Y156_AQ),
.I3(CLBLM_R_X7Y155_SLICE_X8Y155_CO6),
.I4(CLBLM_L_X10Y153_SLICE_X12Y153_AQ),
.I5(CLBLM_R_X7Y158_SLICE_X8Y158_CO5),
.O5(CLBLM_L_X8Y156_SLICE_X11Y156_AO5),
.O6(CLBLM_L_X8Y156_SLICE_X11Y156_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y157_SLICE_X10Y157_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y157_SLICE_X10Y157_AO6),
.Q(CLBLM_L_X8Y157_SLICE_X10Y157_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y157_SLICE_X10Y157_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y157_SLICE_X10Y157_BO6),
.Q(CLBLM_L_X8Y157_SLICE_X10Y157_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y157_SLICE_X10Y157_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y157_SLICE_X10Y157_CO6),
.Q(CLBLM_L_X8Y157_SLICE_X10Y157_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y157_SLICE_X10Y157_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y157_SLICE_X10Y157_DO6),
.Q(CLBLM_L_X8Y157_SLICE_X10Y157_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00cc00cc)
  ) CLBLM_L_X8Y157_SLICE_X10Y157_DLUT (
.I0(CLBLM_R_X5Y149_SLICE_X6Y149_BQ),
.I1(CLBLM_R_X11Y158_SLICE_X14Y158_CQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y159_SLICE_X15Y159_CO6),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y157_SLICE_X10Y157_DO5),
.O6(CLBLM_L_X8Y157_SLICE_X10Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000d0c0d0c0)
  ) CLBLM_L_X8Y157_SLICE_X10Y157_CLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_L_X8Y157_SLICE_X10Y157_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X12Y149_SLICE_X16Y149_CQ),
.I4(CLBLM_L_X8Y150_SLICE_X11Y150_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y157_SLICE_X10Y157_CO5),
.O6(CLBLM_L_X8Y157_SLICE_X10Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00f0ccf0)
  ) CLBLM_L_X8Y157_SLICE_X10Y157_BLUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I1(CLBLM_L_X8Y157_SLICE_X10Y157_BQ),
.I2(CLBLM_L_X8Y156_SLICE_X11Y156_AQ),
.I3(CLBLM_R_X7Y155_SLICE_X8Y155_CO6),
.I4(CLBLM_R_X7Y158_SLICE_X8Y158_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y157_SLICE_X10Y157_BO5),
.O6(CLBLM_L_X8Y157_SLICE_X10Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaffaaf3aaff)
  ) CLBLM_L_X8Y157_SLICE_X10Y157_ALUT (
.I0(CLBLM_R_X11Y158_SLICE_X14Y158_CQ),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLL_L_X4Y158_SLICE_X4Y158_AO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(RIOB33_X105Y135_IOB_X1Y135_I),
.O5(CLBLM_L_X8Y157_SLICE_X10Y157_AO5),
.O6(CLBLM_L_X8Y157_SLICE_X10Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y157_SLICE_X11Y157_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y157_SLICE_X11Y157_AO6),
.Q(CLBLM_L_X8Y157_SLICE_X11Y157_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y157_SLICE_X11Y157_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y157_SLICE_X11Y157_BO6),
.Q(CLBLM_L_X8Y157_SLICE_X11Y157_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y157_SLICE_X11Y157_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y157_SLICE_X11Y157_CO6),
.Q(CLBLM_L_X8Y157_SLICE_X11Y157_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff0f0fffbf)
  ) CLBLM_L_X8Y157_SLICE_X11Y157_DLUT (
.I0(CLBLM_R_X7Y148_SLICE_X8Y148_AQ),
.I1(CLBLM_L_X8Y158_SLICE_X10Y158_AQ),
.I2(CLBLM_R_X7Y155_SLICE_X8Y155_BO5),
.I3(CLBLM_L_X8Y154_SLICE_X10Y154_A5Q),
.I4(CLBLM_R_X7Y155_SLICE_X8Y155_AQ),
.I5(CLBLM_R_X7Y148_SLICE_X8Y148_BQ),
.O5(CLBLM_L_X8Y157_SLICE_X11Y157_DO5),
.O6(CLBLM_L_X8Y157_SLICE_X11Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000cc00cc)
  ) CLBLM_L_X8Y157_SLICE_X11Y157_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y157_SLICE_X11Y157_CQ),
.I2(CLBLM_R_X13Y158_SLICE_X18Y158_BQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y157_SLICE_X11Y157_CO5),
.O6(CLBLM_L_X8Y157_SLICE_X11Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd11dd11cc00cc00)
  ) CLBLM_L_X8Y157_SLICE_X11Y157_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_L_X10Y156_SLICE_X13Y156_BQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y157_SLICE_X12Y157_AQ),
.O5(CLBLM_L_X8Y157_SLICE_X11Y157_BO5),
.O6(CLBLM_L_X8Y157_SLICE_X11Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8bbb8b8888bb8888)
  ) CLBLM_L_X8Y157_SLICE_X11Y157_ALUT (
.I0(CLBLM_R_X11Y149_SLICE_X15Y149_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y158_SLICE_X8Y158_CO5),
.I3(CLBLM_R_X7Y155_SLICE_X8Y155_CO6),
.I4(CLBLM_L_X8Y158_SLICE_X11Y158_AQ),
.I5(CLBLM_L_X8Y157_SLICE_X11Y157_AQ),
.O5(CLBLM_L_X8Y157_SLICE_X11Y157_AO5),
.O6(CLBLM_L_X8Y157_SLICE_X11Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y158_SLICE_X10Y158_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y158_SLICE_X10Y158_AO6),
.Q(CLBLM_L_X8Y158_SLICE_X10Y158_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y158_SLICE_X10Y158_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y158_SLICE_X10Y158_BO6),
.Q(CLBLM_L_X8Y158_SLICE_X10Y158_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y158_SLICE_X10Y158_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y158_SLICE_X10Y158_DO5),
.O6(CLBLM_L_X8Y158_SLICE_X10Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y158_SLICE_X10Y158_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y158_SLICE_X10Y158_CO5),
.O6(CLBLM_L_X8Y158_SLICE_X10Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00ee44ee44)
  ) CLBLM_L_X8Y158_SLICE_X10Y158_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y158_SLICE_X10Y158_BQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y158_SLICE_X9Y158_AQ),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X8Y158_SLICE_X10Y158_BO5),
.O6(CLBLM_L_X8Y158_SLICE_X10Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00b4000000b4)
  ) CLBLM_L_X8Y158_SLICE_X10Y158_ALUT (
.I0(CLBLM_L_X8Y159_SLICE_X10Y159_BO5),
.I1(CLBLM_L_X10Y159_SLICE_X12Y159_AO6),
.I2(CLBLM_L_X8Y158_SLICE_X10Y158_AQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y156_SLICE_X10Y156_CQ),
.O5(CLBLM_L_X8Y158_SLICE_X10Y158_AO5),
.O6(CLBLM_L_X8Y158_SLICE_X10Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y158_SLICE_X11Y158_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y158_SLICE_X11Y158_AO6),
.Q(CLBLM_L_X8Y158_SLICE_X11Y158_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y158_SLICE_X11Y158_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y158_SLICE_X11Y158_BO6),
.Q(CLBLM_L_X8Y158_SLICE_X11Y158_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y158_SLICE_X11Y158_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y158_SLICE_X11Y158_DO5),
.O6(CLBLM_L_X8Y158_SLICE_X11Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y158_SLICE_X11Y158_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y158_SLICE_X11Y158_CO5),
.O6(CLBLM_L_X8Y158_SLICE_X11Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f0f0cccc)
  ) CLBLM_L_X8Y158_SLICE_X11Y158_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X8Y158_SLICE_X11Y158_BQ),
.I2(CLBLM_L_X10Y153_SLICE_X12Y153_BQ),
.I3(CLBLM_R_X11Y152_SLICE_X14Y152_B5Q),
.I4(CLBLM_R_X5Y152_SLICE_X6Y152_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X8Y158_SLICE_X11Y158_BO5),
.O6(CLBLM_L_X8Y158_SLICE_X11Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcceefcee00223022)
  ) CLBLM_L_X8Y158_SLICE_X11Y158_ALUT (
.I0(CLBLM_L_X8Y157_SLICE_X10Y157_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y158_SLICE_X11Y158_AQ),
.I3(CLBLM_R_X7Y155_SLICE_X8Y155_CO6),
.I4(CLBLM_R_X7Y158_SLICE_X8Y158_CO5),
.I5(CLBLM_R_X7Y156_SLICE_X8Y156_DQ),
.O5(CLBLM_L_X8Y158_SLICE_X11Y158_AO5),
.O6(CLBLM_L_X8Y158_SLICE_X11Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X8Y159_SLICE_X10Y159_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X8Y159_SLICE_X10Y159_AO6),
.Q(CLBLM_L_X8Y159_SLICE_X10Y159_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y159_SLICE_X10Y159_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y159_SLICE_X10Y159_DO5),
.O6(CLBLM_L_X8Y159_SLICE_X10Y159_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y159_SLICE_X10Y159_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y159_SLICE_X10Y159_CO5),
.O6(CLBLM_L_X8Y159_SLICE_X10Y159_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h22f26767bb0b5555)
  ) CLBLM_L_X8Y159_SLICE_X10Y159_BLUT (
.I0(CLBLM_R_X7Y148_SLICE_X8Y148_AQ),
.I1(CLBLM_R_X7Y148_SLICE_X8Y148_BQ),
.I2(CLBLM_L_X8Y154_SLICE_X10Y154_A5Q),
.I3(CLBLM_R_X7Y155_SLICE_X8Y155_AQ),
.I4(CLBLM_L_X8Y158_SLICE_X10Y158_AQ),
.I5(1'b1),
.O5(CLBLM_L_X8Y159_SLICE_X10Y159_BO5),
.O6(CLBLM_L_X8Y159_SLICE_X10Y159_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffcfc00000cfc0)
  ) CLBLM_L_X8Y159_SLICE_X10Y159_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y149_SLICE_X9Y149_DO6),
.I2(CLBLM_R_X7Y158_SLICE_X8Y158_CO5),
.I3(CLBLM_R_X7Y159_SLICE_X9Y159_AO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y159_SLICE_X15Y159_AQ),
.O5(CLBLM_L_X8Y159_SLICE_X10Y159_AO5),
.O6(CLBLM_L_X8Y159_SLICE_X10Y159_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y159_SLICE_X11Y159_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y159_SLICE_X11Y159_DO5),
.O6(CLBLM_L_X8Y159_SLICE_X11Y159_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y159_SLICE_X11Y159_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y159_SLICE_X11Y159_CO5),
.O6(CLBLM_L_X8Y159_SLICE_X11Y159_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y159_SLICE_X11Y159_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y159_SLICE_X11Y159_BO5),
.O6(CLBLM_L_X8Y159_SLICE_X11Y159_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafaea55550515)
  ) CLBLM_L_X8Y159_SLICE_X11Y159_ALUT (
.I0(CLBLM_L_X8Y157_SLICE_X11Y157_DO6),
.I1(CLBLM_L_X10Y159_SLICE_X12Y159_BO6),
.I2(CLBLM_L_X8Y157_SLICE_X11Y157_AQ),
.I3(CLBLM_L_X10Y159_SLICE_X13Y159_BO5),
.I4(CLBLM_L_X8Y156_SLICE_X11Y156_DO6),
.I5(CLBLM_R_X11Y159_SLICE_X14Y159_DQ),
.O5(CLBLM_L_X8Y159_SLICE_X11Y159_AO5),
.O6(CLBLM_L_X8Y159_SLICE_X11Y159_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y144_SLICE_X12Y144_AO6),
.Q(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y144_SLICE_X12Y144_DO5),
.O6(CLBLM_L_X10Y144_SLICE_X12Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y144_SLICE_X12Y144_CO5),
.O6(CLBLM_L_X10Y144_SLICE_X12Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y144_SLICE_X12Y144_BO5),
.O6(CLBLM_L_X10Y144_SLICE_X12Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hec20ee220000aaaa)
  ) CLBLM_L_X10Y144_SLICE_X12Y144_ALUT (
.I0(CLBLM_L_X8Y153_SLICE_X10Y153_A5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.I3(CLBLM_L_X10Y147_SLICE_X12Y147_CQ),
.I4(RIOB33_X105Y141_IOB_X1Y142_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y144_SLICE_X12Y144_AO5),
.O6(CLBLM_L_X10Y144_SLICE_X12Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y144_SLICE_X13Y144_DO5),
.O6(CLBLM_L_X10Y144_SLICE_X13Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y144_SLICE_X13Y144_CO5),
.O6(CLBLM_L_X10Y144_SLICE_X13Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y144_SLICE_X13Y144_BO5),
.O6(CLBLM_L_X10Y144_SLICE_X13Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y144_SLICE_X13Y144_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y144_SLICE_X13Y144_AO5),
.O6(CLBLM_L_X10Y144_SLICE_X13Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y145_SLICE_X12Y145_AO6),
.Q(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y145_SLICE_X12Y145_BO6),
.Q(CLBLM_L_X10Y145_SLICE_X12Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y145_SLICE_X12Y145_CO6),
.Q(CLBLM_L_X10Y145_SLICE_X12Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbaaa00009aaa0000)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_DLUT (
.I0(CLBLM_L_X10Y146_SLICE_X12Y146_C5Q),
.I1(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.I2(CLBLM_L_X10Y146_SLICE_X12Y146_CQ),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_CQ),
.I4(CLBLM_L_X8Y148_SLICE_X11Y148_DO6),
.I5(CLBLM_L_X10Y145_SLICE_X13Y145_BQ),
.O5(CLBLM_L_X10Y145_SLICE_X12Y145_DO5),
.O6(CLBLM_L_X10Y145_SLICE_X12Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00fc00fc)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_CLUT (
.I0(CLBLL_L_X4Y151_SLICE_X5Y151_CQ),
.I1(CLBLM_L_X10Y145_SLICE_X12Y145_CQ),
.I2(CLBLM_L_X10Y145_SLICE_X12Y145_BQ),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y145_SLICE_X12Y145_CO5),
.O6(CLBLM_L_X10Y145_SLICE_X12Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000fffc00fc)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y145_SLICE_X12Y145_BQ),
.I2(CLBLM_L_X10Y147_SLICE_X12Y147_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y144_SLICE_X15Y144_AQ),
.I5(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.O5(CLBLM_L_X10Y145_SLICE_X12Y145_BO5),
.O6(CLBLM_L_X10Y145_SLICE_X12Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd11dd11dc10dc10)
  ) CLBLM_L_X10Y145_SLICE_X12Y145_ALUT (
.I0(CLBLM_R_X7Y146_SLICE_X9Y146_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I3(CLBLM_R_X5Y148_SLICE_X7Y148_A5Q),
.I4(1'b1),
.I5(CLBLM_L_X12Y146_SLICE_X16Y146_AQ),
.O5(CLBLM_L_X10Y145_SLICE_X12Y145_AO5),
.O6(CLBLM_L_X10Y145_SLICE_X12Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y145_SLICE_X13Y145_AO6),
.Q(CLBLM_L_X10Y145_SLICE_X13Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y145_SLICE_X13Y145_BO6),
.Q(CLBLM_L_X10Y145_SLICE_X13Y145_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y145_SLICE_X13Y145_CO6),
.Q(CLBLM_L_X10Y145_SLICE_X13Y145_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8080000000080000)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_DLUT (
.I0(CLBLM_L_X10Y146_SLICE_X12Y146_C5Q),
.I1(CLBLM_L_X10Y145_SLICE_X13Y145_CQ),
.I2(CLBLM_L_X10Y145_SLICE_X13Y145_BQ),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.I4(CLBLM_L_X10Y146_SLICE_X12Y146_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y145_SLICE_X13Y145_DO5),
.O6(CLBLM_L_X10Y145_SLICE_X13Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc0ff90c0c09090)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_CLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.I1(CLBLM_L_X10Y145_SLICE_X13Y145_CQ),
.I2(CLBLM_L_X8Y148_SLICE_X11Y148_DO6),
.I3(CLBLM_R_X11Y146_SLICE_X14Y146_CQ),
.I4(CLBLM_L_X10Y145_SLICE_X13Y145_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y145_SLICE_X13Y145_CO5),
.O6(CLBLM_L_X10Y145_SLICE_X13Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0000f0c0)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_BLUT (
.I0(CLBLM_L_X10Y145_SLICE_X12Y145_BQ),
.I1(CLBLM_L_X10Y145_SLICE_X13Y145_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_DO5),
.I4(CLBLM_R_X11Y154_SLICE_X14Y154_DQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y145_SLICE_X13Y145_BO5),
.O6(CLBLM_L_X10Y145_SLICE_X13Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaf0aa30aa30)
  ) CLBLM_L_X10Y145_SLICE_X13Y145_ALUT (
.I0(CLBLM_L_X10Y147_SLICE_X13Y147_CQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X10Y145_SLICE_X13Y145_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.O5(CLBLM_L_X10Y145_SLICE_X13Y145_AO5),
.O6(CLBLM_L_X10Y145_SLICE_X13Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y146_SLICE_X12Y146_CO5),
.Q(CLBLM_L_X10Y146_SLICE_X12Y146_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y146_SLICE_X12Y146_AO6),
.Q(CLBLM_L_X10Y146_SLICE_X12Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y146_SLICE_X12Y146_BO6),
.Q(CLBLM_L_X10Y146_SLICE_X12Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y146_SLICE_X12Y146_CO6),
.Q(CLBLM_L_X10Y146_SLICE_X12Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0b0c0c0c030c0)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_DLUT (
.I0(CLBLM_L_X10Y146_SLICE_X12Y146_C5Q),
.I1(CLBLM_L_X10Y146_SLICE_X12Y146_CQ),
.I2(CLBLM_L_X8Y148_SLICE_X11Y148_DO6),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_CQ),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.I5(CLBLM_L_X10Y145_SLICE_X13Y145_BQ),
.O5(CLBLM_L_X10Y146_SLICE_X12Y146_DO5),
.O6(CLBLM_L_X10Y146_SLICE_X12Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffc0c0ffa0ffa0)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_CLUT (
.I0(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.I1(CLBLM_R_X11Y158_SLICE_X14Y158_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y145_SLICE_X12Y145_DO6),
.I4(CLBLM_L_X10Y146_SLICE_X12Y146_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y146_SLICE_X12Y146_CO5),
.O6(CLBLM_L_X10Y146_SLICE_X12Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fffc000000fc)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y146_SLICE_X12Y146_BQ),
.I2(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_DO6),
.I5(CLBLM_R_X11Y152_SLICE_X14Y152_BQ),
.O5(CLBLM_L_X10Y146_SLICE_X12Y146_BO5),
.O6(CLBLM_L_X10Y146_SLICE_X12Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aaffaa00aaf0)
  ) CLBLM_L_X10Y146_SLICE_X12Y146_ALUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y146_SLICE_X12Y146_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y146_SLICE_X9Y146_DO6),
.I5(CLBLM_L_X8Y147_SLICE_X11Y147_AQ),
.O5(CLBLM_L_X10Y146_SLICE_X12Y146_AO5),
.O6(CLBLM_L_X10Y146_SLICE_X12Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h66ff66ffff66ff66)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_DLUT (
.I0(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I1(CLBLM_R_X11Y152_SLICE_X14Y152_BQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y149_SLICE_X12Y149_CQ),
.I4(1'b1),
.I5(CLBLM_L_X12Y146_SLICE_X16Y146_AQ),
.O5(CLBLM_L_X10Y146_SLICE_X13Y146_DO5),
.O6(CLBLM_L_X10Y146_SLICE_X13Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffeeffee)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_CLUT (
.I0(CLBLM_L_X10Y146_SLICE_X12Y146_AQ),
.I1(CLBLM_L_X10Y147_SLICE_X12Y147_AQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y147_SLICE_X11Y147_AQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y146_SLICE_X9Y146_AQ),
.O5(CLBLM_L_X10Y146_SLICE_X13Y146_CO5),
.O6(CLBLM_L_X10Y146_SLICE_X13Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_BLUT (
.I0(CLBLM_R_X11Y146_SLICE_X15Y146_CQ),
.I1(CLBLM_L_X10Y147_SLICE_X13Y147_BQ),
.I2(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.I3(CLBLM_L_X10Y146_SLICE_X12Y146_BQ),
.I4(CLBLM_L_X8Y146_SLICE_X11Y146_BQ),
.I5(CLBLM_L_X8Y146_SLICE_X11Y146_CQ),
.O5(CLBLM_L_X10Y146_SLICE_X13Y146_BO5),
.O6(CLBLM_L_X10Y146_SLICE_X13Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00ff00fd)
  ) CLBLM_L_X10Y146_SLICE_X13Y146_ALUT (
.I0(CLBLM_L_X10Y146_SLICE_X13Y146_BO6),
.I1(CLBLM_R_X11Y146_SLICE_X15Y146_AQ),
.I2(CLBLM_L_X8Y146_SLICE_X11Y146_AQ),
.I3(CLBLM_R_X11Y146_SLICE_X15Y146_BQ),
.I4(CLBLM_L_X12Y146_SLICE_X16Y146_AQ),
.I5(CLBLM_L_X10Y146_SLICE_X13Y146_CO6),
.O5(CLBLM_L_X10Y146_SLICE_X13Y146_AO5),
.O6(CLBLM_L_X10Y146_SLICE_X13Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y147_SLICE_X12Y147_AO6),
.Q(CLBLM_L_X10Y147_SLICE_X12Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y147_SLICE_X12Y147_BO6),
.Q(CLBLM_L_X10Y147_SLICE_X12Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y147_SLICE_X12Y147_CO6),
.Q(CLBLM_L_X10Y147_SLICE_X12Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y147_SLICE_X12Y147_DO6),
.Q(CLBLM_L_X10Y147_SLICE_X12Y147_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaaaafffff0c0)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_DLUT (
.I0(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.I1(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I2(CLBLM_L_X10Y147_SLICE_X12Y147_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X10Y148_SLICE_X12Y148_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y147_SLICE_X12Y147_DO5),
.O6(CLBLM_L_X10Y147_SLICE_X12Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000fc00fc)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y147_SLICE_X12Y147_CQ),
.I2(CLBLM_L_X12Y148_SLICE_X16Y148_DO6),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.I4(CLBLM_R_X7Y148_SLICE_X8Y148_A5Q),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y147_SLICE_X12Y147_CO5),
.O6(CLBLM_L_X10Y147_SLICE_X12Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff22ff3300220033)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_BLUT (
.I0(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.I1(CLBLM_R_X11Y147_SLICE_X14Y147_BO6),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y141_IOB_X1Y142_I),
.I5(CLBLM_R_X5Y155_SLICE_X7Y155_AQ),
.O5(CLBLM_L_X10Y147_SLICE_X12Y147_BO5),
.O6(CLBLM_L_X10Y147_SLICE_X12Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000fff300f3)
  ) CLBLM_L_X10Y147_SLICE_X12Y147_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y147_SLICE_X13Y147_DO6),
.I2(CLBLM_L_X10Y147_SLICE_X12Y147_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y154_SLICE_X11Y154_AQ),
.I5(CLBLM_R_X7Y146_SLICE_X9Y146_DO6),
.O5(CLBLM_L_X10Y147_SLICE_X12Y147_AO5),
.O6(CLBLM_L_X10Y147_SLICE_X12Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y147_SLICE_X13Y147_AO6),
.Q(CLBLM_L_X10Y147_SLICE_X13Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y147_SLICE_X13Y147_BO6),
.Q(CLBLM_L_X10Y147_SLICE_X13Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y147_SLICE_X13Y147_CO6),
.Q(CLBLM_L_X10Y147_SLICE_X13Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0a0a0cfcfafaf)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_DLUT (
.I0(CLBLM_L_X10Y146_SLICE_X13Y146_AO6),
.I1(CLBLM_R_X11Y146_SLICE_X15Y146_BQ),
.I2(CLBLM_L_X8Y147_SLICE_X10Y147_DO5),
.I3(1'b1),
.I4(CLBLM_R_X11Y146_SLICE_X14Y146_DQ),
.I5(CLBLM_R_X13Y153_SLICE_X18Y153_CQ),
.O5(CLBLM_L_X10Y147_SLICE_X13Y147_DO5),
.O6(CLBLM_L_X10Y147_SLICE_X13Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00cecec4c4)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_CLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X10Y147_SLICE_X13Y147_CQ),
.I2(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I3(CLBLM_R_X11Y146_SLICE_X15Y146_CQ),
.I4(CLBLM_L_X8Y147_SLICE_X11Y147_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y147_SLICE_X13Y147_CO5),
.O6(CLBLM_L_X10Y147_SLICE_X13Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0f000fff0c000c)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y147_SLICE_X13Y147_BQ),
.I2(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y156_SLICE_X12Y156_AQ),
.I5(CLBLM_R_X11Y146_SLICE_X15Y146_CQ),
.O5(CLBLM_L_X10Y147_SLICE_X13Y147_BO5),
.O6(CLBLM_L_X10Y147_SLICE_X13Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ccaaccff)
  ) CLBLM_L_X10Y147_SLICE_X13Y147_ALUT (
.I0(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.I1(CLBLM_L_X10Y150_SLICE_X13Y150_CQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y141_IOB_X1Y142_I),
.I5(CLBLM_R_X11Y147_SLICE_X15Y147_BO6),
.O5(CLBLM_L_X10Y147_SLICE_X13Y147_AO5),
.O6(CLBLM_L_X10Y147_SLICE_X13Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y148_SLICE_X12Y148_AO6),
.Q(CLBLM_L_X10Y148_SLICE_X12Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf100f100f1001100)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_DLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I1(CLBLM_R_X3Y152_SLICE_X3Y152_BO5),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X10Y148_SLICE_X12Y148_CO6),
.I4(CLBLM_L_X8Y150_SLICE_X11Y150_BQ),
.I5(CLBLM_R_X5Y152_SLICE_X6Y152_BQ),
.O5(CLBLM_L_X10Y148_SLICE_X12Y148_DO5),
.O6(CLBLM_L_X10Y148_SLICE_X12Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h332230200f0f0000)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_CLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I3(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y148_SLICE_X12Y148_CO5),
.O6(CLBLM_L_X10Y148_SLICE_X12Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2e2c0aaaaaa00)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_BLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y151_SLICE_X12Y151_AQ),
.I3(CLBLM_L_X10Y147_SLICE_X12Y147_DQ),
.I4(CLBLM_R_X5Y152_SLICE_X6Y152_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y148_SLICE_X12Y148_BO5),
.O6(CLBLM_L_X10Y148_SLICE_X12Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aaf0aa00aaf0)
  ) CLBLM_L_X10Y148_SLICE_X12Y148_ALUT (
.I0(CLBLM_L_X8Y148_SLICE_X11Y148_B5Q),
.I1(1'b1),
.I2(CLBLM_L_X10Y148_SLICE_X12Y148_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y148_SLICE_X12Y148_AO5),
.O6(CLBLM_L_X10Y148_SLICE_X12Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y148_SLICE_X13Y148_AO6),
.Q(CLBLM_L_X10Y148_SLICE_X13Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y148_SLICE_X13Y148_BO6),
.Q(CLBLM_L_X10Y148_SLICE_X13Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y148_SLICE_X13Y148_CO6),
.Q(CLBLM_L_X10Y148_SLICE_X13Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000080000000)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_DLUT (
.I0(CLBLM_L_X10Y148_SLICE_X13Y148_BQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X11Y152_SLICE_X15Y152_DQ),
.I3(CLBLM_L_X10Y155_SLICE_X12Y155_BQ),
.I4(CLBLM_L_X10Y148_SLICE_X13Y148_AQ),
.I5(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.O5(CLBLM_L_X10Y148_SLICE_X13Y148_DO5),
.O6(CLBLM_L_X10Y148_SLICE_X13Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccf0ccfaccf0)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_CLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_L_X12Y146_SLICE_X16Y146_CQ),
.I2(CLBLM_L_X10Y150_SLICE_X13Y150_DO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y148_SLICE_X13Y148_CQ),
.I5(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.O5(CLBLM_L_X10Y148_SLICE_X13Y148_CO5),
.O6(CLBLM_L_X10Y148_SLICE_X13Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haabe0014aaee0044)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y148_SLICE_X13Y148_BQ),
.I2(CLBLM_L_X10Y148_SLICE_X12Y148_CO5),
.I3(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I4(CLBLM_R_X13Y153_SLICE_X18Y153_C5Q),
.I5(CLBLM_L_X10Y155_SLICE_X12Y155_BQ),
.O5(CLBLM_L_X10Y148_SLICE_X13Y148_BO5),
.O6(CLBLM_L_X10Y148_SLICE_X13Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccee0022ccde0012)
  ) CLBLM_L_X10Y148_SLICE_X13Y148_ALUT (
.I0(CLBLM_L_X10Y148_SLICE_X13Y148_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y148_SLICE_X12Y148_CO5),
.I3(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I4(CLBLM_L_X12Y149_SLICE_X17Y149_AQ),
.I5(CLBLM_L_X8Y149_SLICE_X11Y149_DO6),
.O5(CLBLM_L_X10Y148_SLICE_X13Y148_AO5),
.O6(CLBLM_L_X10Y148_SLICE_X13Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y149_SLICE_X12Y149_CO5),
.Q(CLBLM_L_X10Y149_SLICE_X12Y149_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y149_SLICE_X12Y149_AO6),
.Q(CLBLM_L_X10Y149_SLICE_X12Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y149_SLICE_X12Y149_BO6),
.Q(CLBLM_L_X10Y149_SLICE_X12Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y149_SLICE_X12Y149_CO6),
.Q(CLBLM_L_X10Y149_SLICE_X12Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0e4e4f0000000)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y150_SLICE_X5Y150_DQ),
.I2(CLBLM_L_X10Y151_SLICE_X13Y151_B5Q),
.I3(CLBLM_L_X8Y153_SLICE_X10Y153_A5Q),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y149_SLICE_X12Y149_DO5),
.O6(CLBLM_L_X10Y149_SLICE_X12Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4e4fa50aa00)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y149_SLICE_X13Y149_BQ),
.I2(CLBLM_L_X10Y152_SLICE_X12Y152_BQ),
.I3(CLBLM_L_X10Y151_SLICE_X12Y151_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y149_SLICE_X12Y149_CO5),
.O6(CLBLM_L_X10Y149_SLICE_X12Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf077f0fff0fff0ff)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_BLUT (
.I0(CLBLM_L_X10Y151_SLICE_X13Y151_B5Q),
.I1(CLBLM_L_X10Y149_SLICE_X12Y149_BQ),
.I2(CLBLM_L_X10Y149_SLICE_X12Y149_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X8Y153_SLICE_X10Y153_A5Q),
.O5(CLBLM_L_X10Y149_SLICE_X12Y149_BO5),
.O6(CLBLM_L_X10Y149_SLICE_X12Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0bbf0bbf011f0bb)
  ) CLBLM_L_X10Y149_SLICE_X12Y149_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLL_L_X4Y150_SLICE_X5Y150_C5Q),
.I2(CLBLM_L_X12Y157_SLICE_X17Y157_A5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y151_SLICE_X5Y151_CQ),
.I5(CLBLM_L_X8Y148_SLICE_X11Y148_BQ),
.O5(CLBLM_L_X10Y149_SLICE_X12Y149_AO5),
.O6(CLBLM_L_X10Y149_SLICE_X12Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y149_SLICE_X13Y149_BO6),
.Q(CLBLM_L_X10Y149_SLICE_X13Y149_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X10Y149_SLICE_X13Y149_AO6),
.Q(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y150_SLICE_X15Y150_AO6),
.Q(CLBLM_L_X10Y149_SLICE_X13Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000050005)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_DLUT (
.I0(CLBLM_R_X11Y146_SLICE_X14Y146_BQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y153_SLICE_X9Y153_AQ),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_AQ),
.I4(1'b1),
.I5(CLBLM_L_X8Y149_SLICE_X11Y149_BQ),
.O5(CLBLM_L_X10Y149_SLICE_X13Y149_DO5),
.O6(CLBLM_L_X10Y149_SLICE_X13Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000f0e0e0)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_CLUT (
.I0(CLBLL_L_X4Y153_SLICE_X4Y153_BO6),
.I1(CLBLM_R_X13Y155_SLICE_X19Y155_AO6),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X10Y147_SLICE_X13Y147_CQ),
.I4(CLBLM_L_X10Y149_SLICE_X13Y149_DO6),
.I5(CLBLM_L_X12Y151_SLICE_X16Y151_BQ),
.O5(CLBLM_L_X10Y149_SLICE_X13Y149_CO5),
.O6(CLBLM_L_X10Y149_SLICE_X13Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aafc00fc00fc)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_BLUT (
.I0(CLBLM_R_X11Y152_SLICE_X14Y152_CQ),
.I1(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y149_SLICE_X15Y149_BO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y149_SLICE_X13Y149_BO5),
.O6(CLBLM_L_X10Y149_SLICE_X13Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff001010ff001010)
  ) CLBLM_L_X10Y149_SLICE_X13Y149_ALUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.I3(CLBLM_R_X11Y148_SLICE_X14Y148_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y149_SLICE_X13Y149_AO5),
.O6(CLBLM_L_X10Y149_SLICE_X13Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y150_SLICE_X12Y150_AO5),
.Q(CLBLM_L_X10Y150_SLICE_X12Y150_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y150_SLICE_X12Y150_AO6),
.Q(CLBLM_L_X10Y150_SLICE_X12Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y153_SLICE_X13Y153_BO6),
.Q(CLBLM_L_X10Y150_SLICE_X12Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y149_SLICE_X12Y149_DO6),
.Q(CLBLM_L_X10Y150_SLICE_X12Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_DLUT (
.I0(CLBLM_L_X10Y148_SLICE_X12Y148_AQ),
.I1(CLBLM_L_X8Y151_SLICE_X10Y151_BQ),
.I2(CLBLM_L_X10Y151_SLICE_X12Y151_DQ),
.I3(CLBLM_R_X11Y148_SLICE_X14Y148_BQ),
.I4(CLBLM_R_X13Y152_SLICE_X18Y152_A5Q),
.I5(CLBLM_L_X10Y150_SLICE_X12Y150_AQ),
.O5(CLBLM_L_X10Y150_SLICE_X12Y150_DO5),
.O6(CLBLM_L_X10Y150_SLICE_X12Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000200fdff)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_CLUT (
.I0(CLBLM_L_X8Y147_SLICE_X10Y147_CQ),
.I1(CLBLM_L_X8Y150_SLICE_X10Y150_BQ),
.I2(CLBLM_L_X8Y152_SLICE_X10Y152_BQ),
.I3(CLBLM_R_X7Y151_SLICE_X8Y151_CQ),
.I4(CLBLM_R_X13Y152_SLICE_X18Y152_A5Q),
.I5(CLBLM_R_X5Y147_SLICE_X7Y147_BQ),
.O5(CLBLM_L_X10Y150_SLICE_X12Y150_CO5),
.O6(CLBLM_L_X10Y150_SLICE_X12Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f1e0f0feeffeeff)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_BLUT (
.I0(CLBLM_L_X8Y152_SLICE_X10Y152_BQ),
.I1(CLBLM_L_X8Y150_SLICE_X10Y150_BQ),
.I2(CLBLM_L_X10Y150_SLICE_X12Y150_AQ),
.I3(CLBLM_R_X7Y151_SLICE_X8Y151_CQ),
.I4(CLBLM_L_X8Y147_SLICE_X10Y147_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y150_SLICE_X12Y150_BO5),
.O6(CLBLM_L_X10Y150_SLICE_X12Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0f00ff00aaaa)
  ) CLBLM_L_X10Y150_SLICE_X12Y150_ALUT (
.I0(CLBLM_L_X10Y149_SLICE_X12Y149_AQ),
.I1(CLBLM_R_X11Y156_SLICE_X15Y156_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y150_SLICE_X12Y150_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y150_SLICE_X12Y150_AO5),
.O6(CLBLM_L_X10Y150_SLICE_X12Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y150_SLICE_X13Y150_BO5),
.Q(CLBLM_L_X10Y150_SLICE_X13Y150_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y150_SLICE_X13Y150_CO5),
.Q(CLBLM_L_X10Y150_SLICE_X13Y150_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y150_SLICE_X13Y150_AO6),
.Q(CLBLM_L_X10Y150_SLICE_X13Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y150_SLICE_X13Y150_BO6),
.Q(CLBLM_L_X10Y150_SLICE_X13Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y150_SLICE_X13Y150_CO6),
.Q(CLBLM_L_X10Y150_SLICE_X13Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0404000400040004)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_DLUT (
.I0(CLBLM_R_X7Y149_SLICE_X8Y149_DO5),
.I1(CLBLM_R_X7Y154_SLICE_X8Y154_AO5),
.I2(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I3(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y150_SLICE_X9Y150_AO6),
.O5(CLBLM_L_X10Y150_SLICE_X13Y150_DO5),
.O6(CLBLM_L_X10Y150_SLICE_X13Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff000aaccaacc)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_CLUT (
.I0(CLBLM_L_X10Y147_SLICE_X13Y147_AQ),
.I1(CLBLM_L_X10Y150_SLICE_X12Y150_BQ),
.I2(CLBLM_R_X7Y152_SLICE_X9Y152_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y153_SLICE_X12Y153_DO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y150_SLICE_X13Y150_CO5),
.O6(CLBLM_L_X10Y150_SLICE_X13Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aaccf0bbf0bb)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_BLUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_CQ),
.I1(RIOB33_X105Y119_IOB_X1Y119_I),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y150_SLICE_X13Y150_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y150_SLICE_X13Y150_BO5),
.O6(CLBLM_L_X10Y150_SLICE_X13Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaaafaa05000500)
  ) CLBLM_L_X10Y150_SLICE_X13Y150_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X12Y151_SLICE_X16Y151_BQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y147_SLICE_X9Y147_CQ),
.O5(CLBLM_L_X10Y150_SLICE_X13Y150_AO5),
.O6(CLBLM_L_X10Y150_SLICE_X13Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y151_SLICE_X12Y151_AO6),
.Q(CLBLM_L_X10Y151_SLICE_X12Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y151_SLICE_X12Y151_BO6),
.Q(CLBLM_L_X10Y151_SLICE_X12Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y151_SLICE_X12Y151_CO6),
.Q(CLBLM_L_X10Y151_SLICE_X12Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y151_SLICE_X12Y151_DO6),
.Q(CLBLM_L_X10Y151_SLICE_X12Y151_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaf0aa00aa00)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_DLUT (
.I0(CLBLM_R_X5Y150_SLICE_X6Y150_AQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y151_SLICE_X12Y151_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y151_SLICE_X12Y151_DO5),
.O6(CLBLM_L_X10Y151_SLICE_X12Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf000f0ccf0cc)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y151_SLICE_X12Y151_CQ),
.I2(CLBLM_R_X11Y151_SLICE_X14Y151_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X10Y151_SLICE_X12Y151_CO5),
.O6(CLBLM_L_X10Y151_SLICE_X12Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5e4a0e4a0e4a0e4)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y151_SLICE_X14Y151_AQ),
.I2(CLBLM_L_X8Y147_SLICE_X10Y147_CQ),
.I3(CLBLM_R_X11Y149_SLICE_X15Y149_DO6),
.I4(CLBLM_L_X10Y151_SLICE_X12Y151_BQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y151_SLICE_X12Y151_BO5),
.O6(CLBLM_L_X10Y151_SLICE_X12Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffccd80000ccd8)
  ) CLBLM_L_X10Y151_SLICE_X12Y151_ALUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I1(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.I2(CLBLM_L_X10Y151_SLICE_X12Y151_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y153_SLICE_X11Y153_BQ),
.O5(CLBLM_L_X10Y151_SLICE_X12Y151_AO5),
.O6(CLBLM_L_X10Y151_SLICE_X12Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y151_SLICE_X13Y151_BO5),
.Q(CLBLM_L_X10Y151_SLICE_X13Y151_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y151_SLICE_X13Y151_AO6),
.Q(CLBLM_L_X10Y151_SLICE_X13Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y151_SLICE_X13Y151_BO6),
.Q(CLBLM_L_X10Y151_SLICE_X13Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y151_SLICE_X13Y151_CO6),
.Q(CLBLM_L_X10Y151_SLICE_X13Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff9a0000ffaa0000)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_DLUT (
.I0(CLBLM_L_X10Y154_SLICE_X13Y154_C5Q),
.I1(CLBLM_L_X8Y152_SLICE_X10Y152_BQ),
.I2(CLBLM_L_X8Y152_SLICE_X11Y152_BO6),
.I3(CLBLM_L_X10Y158_SLICE_X13Y158_BQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_L_X8Y150_SLICE_X10Y150_BQ),
.O5(CLBLM_L_X10Y151_SLICE_X13Y151_DO5),
.O6(CLBLM_L_X10Y151_SLICE_X13Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f033003300)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_CLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X10Y154_SLICE_X13Y154_CQ),
.I3(CLBLM_L_X10Y158_SLICE_X13Y158_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y151_SLICE_X13Y151_CO5),
.O6(CLBLM_L_X10Y151_SLICE_X13Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf033f000ffaa00aa)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_BLUT (
.I0(CLBLM_L_X8Y153_SLICE_X10Y153_A5Q),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y148_SLICE_X8Y148_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y151_SLICE_X14Y151_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y151_SLICE_X13Y151_BO5),
.O6(CLBLM_L_X10Y151_SLICE_X13Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffa00faffc800c8)
  ) CLBLM_L_X10Y151_SLICE_X13Y151_ALUT (
.I0(CLBLM_L_X10Y151_SLICE_X13Y151_DO6),
.I1(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I2(CLBLM_L_X10Y151_SLICE_X13Y151_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y149_SLICE_X14Y149_BQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X10Y151_SLICE_X13Y151_AO5),
.O6(CLBLM_L_X10Y151_SLICE_X13Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y152_SLICE_X12Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y152_SLICE_X12Y152_AO6),
.Q(CLBLM_L_X10Y152_SLICE_X12Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y152_SLICE_X12Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y152_SLICE_X12Y152_BO6),
.Q(CLBLM_L_X10Y152_SLICE_X12Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa080000fa000000)
  ) CLBLM_L_X10Y152_SLICE_X12Y152_DLUT (
.I0(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.I1(CLBLM_R_X3Y156_SLICE_X2Y156_DO6),
.I2(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I3(CLBLM_L_X10Y152_SLICE_X13Y152_BO6),
.I4(CLBLM_L_X10Y149_SLICE_X13Y149_BO5),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y152_SLICE_X12Y152_DO5),
.O6(CLBLM_L_X10Y152_SLICE_X12Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffa0e400005555)
  ) CLBLM_L_X10Y152_SLICE_X12Y152_CLUT (
.I0(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.I1(CLBLL_L_X4Y154_SLICE_X4Y154_BO6),
.I2(CLBLM_L_X10Y152_SLICE_X13Y152_BO5),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y152_SLICE_X12Y152_CO5),
.O6(CLBLM_L_X10Y152_SLICE_X12Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf505f505f000f000)
  ) CLBLM_L_X10Y152_SLICE_X12Y152_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y153_SLICE_X9Y153_BQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y149_SLICE_X15Y149_A5Q),
.O5(CLBLM_L_X10Y152_SLICE_X12Y152_BO5),
.O6(CLBLM_L_X10Y152_SLICE_X12Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf101f101f404f404)
  ) CLBLM_L_X10Y152_SLICE_X12Y152_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y153_SLICE_X12Y153_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y149_SLICE_X12Y149_C5Q),
.I4(1'b1),
.I5(CLBLM_L_X10Y152_SLICE_X13Y152_BO6),
.O5(CLBLM_L_X10Y152_SLICE_X12Y152_AO5),
.O6(CLBLM_L_X10Y152_SLICE_X12Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y152_SLICE_X13Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y152_SLICE_X13Y152_AO6),
.Q(CLBLM_L_X10Y152_SLICE_X13Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c040c0c0f0f0)
  ) CLBLM_L_X10Y152_SLICE_X13Y152_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X11Y152_SLICE_X14Y152_DO5),
.I2(CLBLM_L_X10Y149_SLICE_X13Y149_BO5),
.I3(CLBLL_L_X4Y154_SLICE_X4Y154_BO6),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I5(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.O5(CLBLM_L_X10Y152_SLICE_X13Y152_DO5),
.O6(CLBLM_L_X10Y152_SLICE_X13Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h44000000f0000000)
  ) CLBLM_L_X10Y152_SLICE_X13Y152_CLUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X10Y148_SLICE_X13Y148_AQ),
.I3(CLBLM_L_X10Y155_SLICE_X12Y155_BQ),
.I4(CLBLM_L_X10Y148_SLICE_X13Y148_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y152_SLICE_X13Y152_CO5),
.O6(CLBLM_L_X10Y152_SLICE_X13Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc8c8c8c8cccccc00)
  ) CLBLM_L_X10Y152_SLICE_X13Y152_BLUT (
.I0(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X10Y152_SLICE_X13Y152_AQ),
.I3(CLBLM_R_X5Y147_SLICE_X7Y147_BQ),
.I4(CLBLM_L_X12Y151_SLICE_X17Y151_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y152_SLICE_X13Y152_BO5),
.O6(CLBLM_L_X10Y152_SLICE_X13Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc4ffc8c4c4c8c8)
  ) CLBLM_L_X10Y152_SLICE_X13Y152_ALUT (
.I0(CLBLM_L_X8Y152_SLICE_X11Y152_DO6),
.I1(CLBLM_L_X10Y149_SLICE_X13Y149_BO5),
.I2(CLBLM_L_X10Y152_SLICE_X13Y152_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y149_SLICE_X13Y149_CO6),
.I5(CLBLM_L_X10Y153_SLICE_X13Y153_CQ),
.O5(CLBLM_L_X10Y152_SLICE_X13Y152_AO5),
.O6(CLBLM_L_X10Y152_SLICE_X13Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y153_SLICE_X12Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y153_SLICE_X12Y153_AO6),
.Q(CLBLM_L_X10Y153_SLICE_X12Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y153_SLICE_X12Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y153_SLICE_X12Y153_BO6),
.Q(CLBLM_L_X10Y153_SLICE_X12Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0609060990609060)
  ) CLBLM_L_X10Y153_SLICE_X12Y153_DLUT (
.I0(CLBLM_L_X10Y152_SLICE_X12Y152_AQ),
.I1(CLBLL_L_X4Y153_SLICE_X5Y153_AQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y153_SLICE_X12Y153_BQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y150_SLICE_X13Y150_CQ),
.O5(CLBLM_L_X10Y153_SLICE_X12Y153_DO5),
.O6(CLBLM_L_X10Y153_SLICE_X12Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0040000000000000)
  ) CLBLM_L_X10Y153_SLICE_X12Y153_CLUT (
.I0(CLBLM_R_X13Y149_SLICE_X18Y149_A5Q),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X10Y154_SLICE_X12Y154_DQ),
.I3(CLBLM_R_X11Y149_SLICE_X15Y149_A5Q),
.I4(CLBLM_R_X11Y153_SLICE_X15Y153_AQ),
.I5(CLBLM_R_X7Y154_SLICE_X8Y154_AO5),
.O5(CLBLM_L_X10Y153_SLICE_X12Y153_CO5),
.O6(CLBLM_L_X10Y153_SLICE_X12Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hababaeae01010404)
  ) CLBLM_L_X10Y153_SLICE_X12Y153_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y152_SLICE_X14Y152_DO5),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(1'b1),
.I4(CLBLM_R_X5Y150_SLICE_X6Y150_AQ),
.I5(CLBLM_L_X12Y154_SLICE_X17Y154_A5Q),
.O5(CLBLM_L_X10Y153_SLICE_X12Y153_BO5),
.O6(CLBLM_L_X10Y153_SLICE_X12Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaee0044faee5044)
  ) CLBLM_L_X10Y153_SLICE_X12Y153_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y155_SLICE_X12Y155_AQ),
.I2(CLBLM_L_X10Y153_SLICE_X12Y153_AQ),
.I3(CLBLM_R_X7Y155_SLICE_X8Y155_CO6),
.I4(CLBLM_L_X10Y147_SLICE_X12Y147_DQ),
.I5(CLBLM_R_X7Y158_SLICE_X8Y158_CO5),
.O5(CLBLM_L_X10Y153_SLICE_X12Y153_AO5),
.O6(CLBLM_L_X10Y153_SLICE_X12Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y153_SLICE_X13Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y153_SLICE_X13Y153_AO6),
.Q(CLBLM_L_X10Y153_SLICE_X13Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y153_SLICE_X13Y153_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y153_SLICE_X13Y153_CO6),
.Q(CLBLM_L_X10Y153_SLICE_X13Y153_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y153_SLICE_X13Y153_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y153_SLICE_X13Y153_DO6),
.Q(CLBLM_L_X10Y153_SLICE_X13Y153_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000cccc5a5a)
  ) CLBLM_L_X10Y153_SLICE_X13Y153_DLUT (
.I0(CLBLM_L_X10Y156_SLICE_X12Y156_AQ),
.I1(CLBLM_L_X10Y151_SLICE_X13Y151_CQ),
.I2(CLBLM_L_X12Y153_SLICE_X16Y153_BO5),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X10Y153_SLICE_X13Y153_DO5),
.O6(CLBLM_L_X10Y153_SLICE_X13Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f5f5f000050500)
  ) CLBLM_L_X10Y153_SLICE_X13Y153_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y154_SLICE_X14Y154_CQ),
.I4(CLBLM_L_X10Y153_SLICE_X13Y153_BO5),
.I5(CLBLM_R_X7Y153_SLICE_X9Y153_AQ),
.O5(CLBLM_L_X10Y153_SLICE_X13Y153_CO5),
.O6(CLBLM_L_X10Y153_SLICE_X13Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ec20aaaaa0a0)
  ) CLBLM_L_X10Y153_SLICE_X13Y153_BLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y153_SLICE_X14Y153_AQ),
.I3(CLBLL_L_X4Y155_SLICE_X4Y155_AQ),
.I4(CLBLM_L_X10Y151_SLICE_X13Y151_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y153_SLICE_X13Y153_BO5),
.O6(CLBLM_L_X10Y153_SLICE_X13Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeeeefa44444450)
  ) CLBLM_L_X10Y153_SLICE_X13Y153_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y153_SLICE_X6Y153_AQ),
.I2(CLBLM_L_X10Y153_SLICE_X13Y153_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I5(CLBLM_R_X11Y157_SLICE_X14Y157_CQ),
.O5(CLBLM_L_X10Y153_SLICE_X13Y153_AO5),
.O6(CLBLM_L_X10Y153_SLICE_X13Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y154_SLICE_X12Y154_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y154_SLICE_X12Y154_BO6),
.Q(CLBLM_L_X10Y154_SLICE_X12Y154_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y154_SLICE_X12Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y154_SLICE_X12Y154_AO6),
.Q(CLBLM_L_X10Y154_SLICE_X12Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y154_SLICE_X12Y154_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y154_SLICE_X12Y154_CO6),
.Q(CLBLM_L_X10Y154_SLICE_X12Y154_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y154_SLICE_X12Y154_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y154_SLICE_X12Y154_DO6),
.Q(CLBLM_L_X10Y154_SLICE_X12Y154_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff451000004510)
  ) CLBLM_L_X10Y154_SLICE_X12Y154_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y154_SLICE_X13Y154_AO5),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X8Y155_SLICE_X11Y155_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y154_SLICE_X12Y154_CQ),
.O5(CLBLM_L_X10Y154_SLICE_X12Y154_DO5),
.O6(CLBLM_L_X10Y154_SLICE_X12Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ffffff00aaaa)
  ) CLBLM_L_X10Y154_SLICE_X12Y154_CLUT (
.I0(CLBLM_R_X11Y159_SLICE_X15Y159_CO6),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X4Y150_SLICE_X5Y150_C5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y153_SLICE_X11Y153_BQ),
.O5(CLBLM_L_X10Y154_SLICE_X12Y154_CO5),
.O6(CLBLM_L_X10Y154_SLICE_X12Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44aa000f0f0000)
  ) CLBLM_L_X10Y154_SLICE_X12Y154_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y154_SLICE_X12Y154_A5Q),
.I2(CLBLM_R_X7Y153_SLICE_X8Y153_AQ),
.I3(CLBLM_R_X11Y153_SLICE_X14Y153_AQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y154_SLICE_X12Y154_BO5),
.O6(CLBLM_L_X10Y154_SLICE_X12Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888d8d8d8d8)
  ) CLBLM_L_X10Y154_SLICE_X12Y154_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y154_SLICE_X14Y154_AQ),
.I2(CLBLM_L_X10Y154_SLICE_X12Y154_AQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y156_SLICE_X12Y156_AQ),
.I5(CLBLM_R_X7Y153_SLICE_X9Y153_CO6),
.O5(CLBLM_L_X10Y154_SLICE_X12Y154_AO5),
.O6(CLBLM_L_X10Y154_SLICE_X12Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y154_SLICE_X13Y154_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y154_SLICE_X13Y154_CO5),
.Q(CLBLM_L_X10Y154_SLICE_X13Y154_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y154_SLICE_X13Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y154_SLICE_X13Y154_AO6),
.Q(CLBLM_L_X10Y154_SLICE_X13Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y154_SLICE_X13Y154_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y154_SLICE_X13Y154_BO6),
.Q(CLBLM_L_X10Y154_SLICE_X13Y154_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y154_SLICE_X13Y154_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y154_SLICE_X13Y154_CO6),
.Q(CLBLM_L_X10Y154_SLICE_X13Y154_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y154_SLICE_X13Y154_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y154_SLICE_X13Y154_DO6),
.Q(CLBLM_L_X10Y154_SLICE_X13Y154_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcffa800fc00a8)
  ) CLBLM_L_X10Y154_SLICE_X13Y154_DLUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I1(CLBLM_R_X7Y152_SLICE_X9Y152_CO6),
.I2(CLBLM_L_X10Y154_SLICE_X13Y154_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X5Y152_SLICE_X6Y152_AQ),
.O5(CLBLM_L_X10Y154_SLICE_X13Y154_DO5),
.O6(CLBLM_L_X10Y154_SLICE_X13Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0afa0aa3a3a0a0)
  ) CLBLM_L_X10Y154_SLICE_X13Y154_CLUT (
.I0(CLBLM_L_X12Y154_SLICE_X17Y154_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y154_SLICE_X10Y154_C5Q),
.I4(CLBLM_L_X10Y154_SLICE_X13Y154_C5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y154_SLICE_X13Y154_CO5),
.O6(CLBLM_L_X10Y154_SLICE_X13Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff300030ff300030)
  ) CLBLM_L_X10Y154_SLICE_X13Y154_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y154_SLICE_X10Y154_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y154_SLICE_X13Y154_BO5),
.O6(CLBLM_L_X10Y154_SLICE_X13Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaacca000000f0f)
  ) CLBLM_L_X10Y154_SLICE_X13Y154_ALUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_L_X10Y154_SLICE_X13Y154_BQ),
.I2(CLBLM_R_X11Y153_SLICE_X15Y153_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X10Y154_SLICE_X13Y154_AO5),
.O6(CLBLM_L_X10Y154_SLICE_X13Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y155_SLICE_X12Y155_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y155_SLICE_X12Y155_AO6),
.Q(CLBLM_L_X10Y155_SLICE_X12Y155_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y155_SLICE_X12Y155_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y155_SLICE_X12Y155_BO6),
.Q(CLBLM_L_X10Y155_SLICE_X12Y155_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y155_SLICE_X12Y155_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y155_SLICE_X12Y155_CO6),
.Q(CLBLM_L_X10Y155_SLICE_X12Y155_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffeeffee)
  ) CLBLM_L_X10Y155_SLICE_X12Y155_DLUT (
.I0(CLBLM_L_X10Y154_SLICE_X12Y154_A5Q),
.I1(CLBLM_L_X10Y155_SLICE_X13Y155_AQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y158_SLICE_X10Y158_BQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y154_SLICE_X13Y154_C5Q),
.O5(CLBLM_L_X10Y155_SLICE_X12Y155_DO5),
.O6(CLBLM_L_X10Y155_SLICE_X12Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff05ff5000050050)
  ) CLBLM_L_X10Y155_SLICE_X12Y155_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(CLBLM_L_X10Y148_SLICE_X12Y148_BO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y156_SLICE_X13Y156_BQ),
.I5(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.O5(CLBLM_L_X10Y155_SLICE_X12Y155_CO5),
.O6(CLBLM_L_X10Y155_SLICE_X12Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaafcfcf3fc)
  ) CLBLM_L_X10Y155_SLICE_X12Y155_BLUT (
.I0(CLBLM_L_X10Y155_SLICE_X12Y155_CQ),
.I1(CLBLM_L_X10Y155_SLICE_X12Y155_BQ),
.I2(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y155_SLICE_X12Y155_BO5),
.O6(CLBLM_L_X10Y155_SLICE_X12Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa3300f3c0)
  ) CLBLM_L_X10Y155_SLICE_X12Y155_ALUT (
.I0(CLBLM_R_X11Y146_SLICE_X14Y146_DQ),
.I1(CLBLM_R_X7Y155_SLICE_X8Y155_CO6),
.I2(CLBLM_L_X10Y155_SLICE_X12Y155_AQ),
.I3(CLBLM_R_X7Y157_SLICE_X9Y157_AQ),
.I4(CLBLM_R_X7Y158_SLICE_X8Y158_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X10Y155_SLICE_X12Y155_AO5),
.O6(CLBLM_L_X10Y155_SLICE_X12Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y155_SLICE_X13Y155_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y155_SLICE_X13Y155_AO5),
.Q(CLBLM_L_X10Y155_SLICE_X13Y155_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y155_SLICE_X13Y155_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y155_SLICE_X13Y155_AO6),
.Q(CLBLM_L_X10Y155_SLICE_X13Y155_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y155_SLICE_X13Y155_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y155_SLICE_X13Y155_BO6),
.Q(CLBLM_L_X10Y155_SLICE_X13Y155_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff2fffffffff)
  ) CLBLM_L_X10Y155_SLICE_X13Y155_DLUT (
.I0(CLBLM_L_X10Y155_SLICE_X13Y155_BQ),
.I1(CLBLM_R_X7Y154_SLICE_X8Y154_AO5),
.I2(CLBLM_L_X10Y156_SLICE_X13Y156_AO5),
.I3(CLBLM_L_X10Y156_SLICE_X13Y156_CO6),
.I4(CLBLM_R_X11Y153_SLICE_X14Y153_DO6),
.I5(CLBLM_L_X10Y152_SLICE_X13Y152_CO5),
.O5(CLBLM_L_X10Y155_SLICE_X13Y155_DO5),
.O6(CLBLM_L_X10Y155_SLICE_X13Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffeeffea)
  ) CLBLM_L_X10Y155_SLICE_X13Y155_CLUT (
.I0(CLBLM_L_X8Y152_SLICE_X11Y152_AO6),
.I1(CLBLM_R_X7Y153_SLICE_X9Y153_CO6),
.I2(CLBLM_R_X11Y152_SLICE_X14Y152_AQ),
.I3(CLBLM_L_X8Y156_SLICE_X11Y156_DO6),
.I4(CLBLM_L_X8Y153_SLICE_X11Y153_CQ),
.I5(CLBLM_L_X10Y155_SLICE_X13Y155_DO6),
.O5(CLBLM_L_X10Y155_SLICE_X13Y155_CO5),
.O6(CLBLM_L_X10Y155_SLICE_X13Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaccaaffaac0)
  ) CLBLM_L_X10Y155_SLICE_X13Y155_BLUT (
.I0(CLBLM_R_X5Y157_SLICE_X7Y157_AQ),
.I1(CLBLM_L_X10Y155_SLICE_X13Y155_BQ),
.I2(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y150_SLICE_X13Y150_DO6),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X10Y155_SLICE_X13Y155_BO5),
.O6(CLBLM_L_X10Y155_SLICE_X13Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he2e2c0c0bb88bb88)
  ) CLBLM_L_X10Y155_SLICE_X13Y155_ALUT (
.I0(CLBLM_L_X10Y155_SLICE_X13Y155_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_AQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y155_SLICE_X13Y155_AO5),
.O6(CLBLM_L_X10Y155_SLICE_X13Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y156_SLICE_X12Y156_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y156_SLICE_X12Y156_AO6),
.Q(CLBLM_L_X10Y156_SLICE_X12Y156_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffff7)
  ) CLBLM_L_X10Y156_SLICE_X12Y156_DLUT (
.I0(CLBLM_L_X8Y153_SLICE_X11Y153_CQ),
.I1(CLBLM_L_X12Y149_SLICE_X16Y149_CQ),
.I2(CLBLM_R_X13Y150_SLICE_X18Y150_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_L_X10Y156_SLICE_X12Y156_DO5),
.O6(CLBLM_L_X10Y156_SLICE_X12Y156_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000200)
  ) CLBLM_L_X10Y156_SLICE_X12Y156_CLUT (
.I0(CLBLM_L_X8Y155_SLICE_X11Y155_CQ),
.I1(CLBLM_L_X8Y156_SLICE_X10Y156_CQ),
.I2(CLBLM_L_X10Y154_SLICE_X12Y154_DQ),
.I3(CLBLM_L_X12Y158_SLICE_X16Y158_A5Q),
.I4(CLBLM_L_X10Y153_SLICE_X13Y153_DQ),
.I5(CLBLM_L_X8Y155_SLICE_X11Y155_BQ),
.O5(CLBLM_L_X10Y156_SLICE_X12Y156_CO5),
.O6(CLBLM_L_X10Y156_SLICE_X12Y156_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001000000000000)
  ) CLBLM_L_X10Y156_SLICE_X12Y156_BLUT (
.I0(CLBLM_L_X10Y156_SLICE_X12Y156_DO6),
.I1(CLBLM_L_X10Y156_SLICE_X13Y156_DO6),
.I2(CLBLM_L_X10Y156_SLICE_X12Y156_AQ),
.I3(CLBLM_L_X10Y153_SLICE_X13Y153_CQ),
.I4(CLBLM_L_X10Y156_SLICE_X12Y156_CO6),
.I5(CLBLM_L_X10Y155_SLICE_X12Y155_CQ),
.O5(CLBLM_L_X10Y156_SLICE_X12Y156_BO5),
.O6(CLBLM_L_X10Y156_SLICE_X12Y156_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff050005ff0a000a)
  ) CLBLM_L_X10Y156_SLICE_X12Y156_ALUT (
.I0(CLBLM_R_X11Y154_SLICE_X15Y154_CO5),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y159_SLICE_X8Y159_AQ),
.I5(CLBLM_L_X10Y155_SLICE_X12Y155_CQ),
.O5(CLBLM_L_X10Y156_SLICE_X12Y156_AO5),
.O6(CLBLM_L_X10Y156_SLICE_X12Y156_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y156_SLICE_X13Y156_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y156_SLICE_X13Y156_BO6),
.Q(CLBLM_L_X10Y156_SLICE_X13Y156_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffdddd)
  ) CLBLM_L_X10Y156_SLICE_X13Y156_DLUT (
.I0(CLBLM_L_X10Y156_SLICE_X13Y156_BQ),
.I1(CLBLM_R_X13Y151_SLICE_X18Y151_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X13Y155_SLICE_X18Y155_BQ),
.I5(CLBLM_R_X11Y154_SLICE_X14Y154_CQ),
.O5(CLBLM_L_X10Y156_SLICE_X13Y156_DO5),
.O6(CLBLM_L_X10Y156_SLICE_X13Y156_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff7fff7fff7f7f7f)
  ) CLBLM_L_X10Y156_SLICE_X13Y156_CLUT (
.I0(CLBLM_L_X10Y157_SLICE_X12Y157_BQ),
.I1(CLBLM_L_X12Y157_SLICE_X16Y157_CQ),
.I2(CLBLM_R_X11Y156_SLICE_X15Y156_AQ),
.I3(CLBLM_R_X7Y148_SLICE_X8Y148_AQ),
.I4(CLBLM_L_X8Y158_SLICE_X10Y158_AQ),
.I5(CLBLM_R_X7Y148_SLICE_X8Y148_BQ),
.O5(CLBLM_L_X10Y156_SLICE_X13Y156_CO5),
.O6(CLBLM_L_X10Y156_SLICE_X13Y156_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8d888d88888d888d)
  ) CLBLM_L_X10Y156_SLICE_X13Y156_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y158_SLICE_X11Y158_AQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y153_SLICE_X13Y153_CQ),
.I4(1'b1),
.I5(CLBLM_L_X12Y152_SLICE_X16Y152_AO5),
.O5(CLBLM_L_X10Y156_SLICE_X13Y156_BO5),
.O6(CLBLM_L_X10Y156_SLICE_X13Y156_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033003333cc33cc)
  ) CLBLM_L_X10Y156_SLICE_X13Y156_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y148_SLICE_X8Y148_BQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y148_SLICE_X8Y148_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y156_SLICE_X13Y156_AO5),
.O6(CLBLM_L_X10Y156_SLICE_X13Y156_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y157_SLICE_X12Y157_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y157_SLICE_X12Y157_AO6),
.Q(CLBLM_L_X10Y157_SLICE_X12Y157_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y157_SLICE_X12Y157_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y157_SLICE_X12Y157_BO6),
.Q(CLBLM_L_X10Y157_SLICE_X12Y157_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff000037f7)
  ) CLBLM_L_X10Y157_SLICE_X12Y157_DLUT (
.I0(CLBLM_L_X10Y157_SLICE_X12Y157_CO5),
.I1(CLBLM_L_X8Y156_SLICE_X11Y156_AQ),
.I2(CLBLM_L_X10Y158_SLICE_X12Y158_BQ),
.I3(CLBLM_L_X10Y157_SLICE_X12Y157_CO6),
.I4(CLBLM_L_X8Y157_SLICE_X11Y157_DO6),
.I5(CLBLM_L_X8Y156_SLICE_X11Y156_DO6),
.O5(CLBLM_L_X10Y157_SLICE_X12Y157_DO5),
.O6(CLBLM_L_X10Y157_SLICE_X12Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33003300000f000f)
  ) CLBLM_L_X10Y157_SLICE_X12Y157_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y156_SLICE_X13Y156_CO6),
.I2(CLBLM_L_X10Y157_SLICE_X13Y157_DO6),
.I3(CLBLM_R_X11Y156_SLICE_X14Y156_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y157_SLICE_X12Y157_CO5),
.O6(CLBLM_L_X10Y157_SLICE_X12Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeffee00ee00ee)
  ) CLBLM_L_X10Y157_SLICE_X12Y157_BLUT (
.I0(CLBLM_L_X10Y159_SLICE_X12Y159_CO6),
.I1(CLBLM_L_X10Y157_SLICE_X13Y157_BO6),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y157_SLICE_X9Y157_DQ),
.O5(CLBLM_L_X10Y157_SLICE_X12Y157_BO5),
.O6(CLBLM_L_X10Y157_SLICE_X12Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0f000fff000000)
  ) CLBLM_L_X10Y157_SLICE_X12Y157_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y155_SLICE_X12Y155_AQ),
.I5(CLBLM_L_X10Y150_SLICE_X12Y150_CQ),
.O5(CLBLM_L_X10Y157_SLICE_X12Y157_AO5),
.O6(CLBLM_L_X10Y157_SLICE_X12Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffff57)
  ) CLBLM_L_X10Y157_SLICE_X13Y157_DLUT (
.I0(CLBLM_R_X7Y148_SLICE_X8Y148_AQ),
.I1(CLBLM_R_X7Y148_SLICE_X8Y148_BQ),
.I2(CLBLM_L_X8Y158_SLICE_X10Y158_AQ),
.I3(CLBLM_L_X12Y157_SLICE_X16Y157_CQ),
.I4(CLBLM_R_X11Y156_SLICE_X15Y156_AQ),
.I5(CLBLM_L_X10Y157_SLICE_X12Y157_BQ),
.O5(CLBLM_L_X10Y157_SLICE_X13Y157_DO5),
.O6(CLBLM_L_X10Y157_SLICE_X13Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a5a5a9a5a9a5a9)
  ) CLBLM_L_X10Y157_SLICE_X13Y157_CLUT (
.I0(CLBLM_R_X11Y156_SLICE_X14Y156_BQ),
.I1(CLBLM_L_X10Y155_SLICE_X12Y155_AQ),
.I2(CLBLM_L_X8Y157_SLICE_X11Y157_DO6),
.I3(CLBLM_L_X8Y156_SLICE_X11Y156_DO6),
.I4(CLBLM_L_X10Y157_SLICE_X13Y157_DO6),
.I5(CLBLM_L_X10Y156_SLICE_X13Y156_CO6),
.O5(CLBLM_L_X10Y157_SLICE_X13Y157_CO5),
.O6(CLBLM_L_X10Y157_SLICE_X13Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h50a050a010e050a0)
  ) CLBLM_L_X10Y157_SLICE_X13Y157_BLUT (
.I0(CLBLM_L_X8Y157_SLICE_X11Y157_DO6),
.I1(CLBLM_R_X7Y157_SLICE_X9Y157_AQ),
.I2(CLBLM_L_X10Y159_SLICE_X12Y159_DO6),
.I3(CLBLM_L_X10Y157_SLICE_X12Y157_BQ),
.I4(CLBLM_L_X10Y157_SLICE_X13Y157_AO6),
.I5(CLBLM_L_X8Y156_SLICE_X11Y156_DO6),
.O5(CLBLM_L_X10Y157_SLICE_X13Y157_BO5),
.O6(CLBLM_L_X10Y157_SLICE_X13Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h10f00e0011ff11ff)
  ) CLBLM_L_X10Y157_SLICE_X13Y157_ALUT (
.I0(CLBLM_L_X8Y158_SLICE_X10Y158_AQ),
.I1(CLBLM_R_X7Y148_SLICE_X8Y148_BQ),
.I2(CLBLM_R_X11Y156_SLICE_X15Y156_AQ),
.I3(CLBLM_R_X7Y148_SLICE_X8Y148_AQ),
.I4(CLBLM_L_X12Y157_SLICE_X16Y157_CQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y157_SLICE_X13Y157_AO5),
.O6(CLBLM_L_X10Y157_SLICE_X13Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y158_SLICE_X12Y158_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y158_SLICE_X12Y158_AO6),
.Q(CLBLM_L_X10Y158_SLICE_X12Y158_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y158_SLICE_X12Y158_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y158_SLICE_X12Y158_BO6),
.Q(CLBLM_L_X10Y158_SLICE_X12Y158_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y158_SLICE_X12Y158_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y158_SLICE_X12Y158_DO5),
.O6(CLBLM_L_X10Y158_SLICE_X12Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0f0f0f0c0f0d0f)
  ) CLBLM_L_X10Y158_SLICE_X12Y158_CLUT (
.I0(CLBLM_R_X11Y156_SLICE_X14Y156_BQ),
.I1(CLBLM_L_X8Y156_SLICE_X11Y156_DO6),
.I2(CLBLM_L_X8Y157_SLICE_X11Y157_DO6),
.I3(CLBLM_L_X10Y153_SLICE_X12Y153_AQ),
.I4(CLBLM_L_X10Y157_SLICE_X12Y157_CO5),
.I5(CLBLM_L_X10Y156_SLICE_X13Y156_CO6),
.O5(CLBLM_L_X10Y158_SLICE_X12Y158_CO5),
.O6(CLBLM_L_X10Y158_SLICE_X12Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffea00eaffba00ba)
  ) CLBLM_L_X10Y158_SLICE_X12Y158_BLUT (
.I0(CLBLM_L_X10Y159_SLICE_X12Y159_CO6),
.I1(CLBLM_L_X10Y158_SLICE_X12Y158_BQ),
.I2(CLBLM_L_X10Y159_SLICE_X12Y159_DO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y153_SLICE_X15Y153_AQ),
.I5(CLBLM_L_X10Y158_SLICE_X12Y158_CO6),
.O5(CLBLM_L_X10Y158_SLICE_X12Y158_BO5),
.O6(CLBLM_L_X10Y158_SLICE_X12Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heefceecceefceecc)
  ) CLBLM_L_X10Y158_SLICE_X12Y158_ALUT (
.I0(CLBLM_L_X10Y146_SLICE_X12Y146_BQ),
.I1(CLBLM_L_X10Y156_SLICE_X12Y156_BO6),
.I2(CLBLM_L_X10Y158_SLICE_X12Y158_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y158_SLICE_X12Y158_AO5),
.O6(CLBLM_L_X10Y158_SLICE_X12Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y158_SLICE_X13Y158_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y158_SLICE_X13Y158_AO6),
.Q(CLBLM_L_X10Y158_SLICE_X13Y158_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X10Y158_SLICE_X13Y158_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X10Y158_SLICE_X13Y158_BO6),
.Q(CLBLM_L_X10Y158_SLICE_X13Y158_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y158_SLICE_X13Y158_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y158_SLICE_X13Y158_DO5),
.O6(CLBLM_L_X10Y158_SLICE_X13Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3030c0c0303060c0)
  ) CLBLM_L_X10Y158_SLICE_X13Y158_CLUT (
.I0(CLBLM_L_X10Y159_SLICE_X13Y159_AO6),
.I1(CLBLM_R_X11Y160_SLICE_X14Y160_AQ),
.I2(CLBLM_L_X10Y159_SLICE_X12Y159_DO6),
.I3(CLBLM_L_X8Y157_SLICE_X10Y157_BQ),
.I4(CLBLM_L_X8Y157_SLICE_X11Y157_DO6),
.I5(CLBLM_L_X8Y156_SLICE_X11Y156_DO6),
.O5(CLBLM_L_X10Y158_SLICE_X13Y158_CO5),
.O6(CLBLM_L_X10Y158_SLICE_X13Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hecec2020ecec2020)
  ) CLBLM_L_X10Y158_SLICE_X13Y158_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y152_SLICE_X17Y152_AQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y158_SLICE_X12Y158_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y158_SLICE_X13Y158_BO5),
.O6(CLBLM_L_X10Y158_SLICE_X13Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa33aaffaa30)
  ) CLBLM_L_X10Y158_SLICE_X13Y158_ALUT (
.I0(CLBLM_L_X8Y157_SLICE_X10Y157_CQ),
.I1(CLBLM_R_X11Y159_SLICE_X15Y159_DO5),
.I2(CLBLM_L_X10Y158_SLICE_X13Y158_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y158_SLICE_X15Y158_BO6),
.I5(CLBLM_R_X11Y157_SLICE_X14Y157_CQ),
.O5(CLBLM_L_X10Y158_SLICE_X13Y158_AO5),
.O6(CLBLM_L_X10Y158_SLICE_X13Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff030000ffcf)
  ) CLBLM_L_X10Y159_SLICE_X12Y159_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y159_SLICE_X14Y159_DQ),
.I2(CLBLM_L_X10Y159_SLICE_X13Y159_BO5),
.I3(CLBLM_L_X8Y156_SLICE_X11Y156_DO6),
.I4(CLBLM_R_X7Y158_SLICE_X8Y158_CO5),
.I5(CLBLM_L_X10Y159_SLICE_X12Y159_BO6),
.O5(CLBLM_L_X10Y159_SLICE_X12Y159_DO5),
.O6(CLBLM_L_X10Y159_SLICE_X12Y159_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000fc00000030)
  ) CLBLM_L_X10Y159_SLICE_X12Y159_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y159_SLICE_X14Y159_DQ),
.I2(CLBLM_L_X10Y159_SLICE_X13Y159_BO5),
.I3(CLBLM_L_X8Y156_SLICE_X11Y156_DO6),
.I4(CLBLM_L_X8Y159_SLICE_X10Y159_BO6),
.I5(CLBLM_L_X10Y159_SLICE_X12Y159_BO6),
.O5(CLBLM_L_X10Y159_SLICE_X12Y159_CO5),
.O6(CLBLM_L_X10Y159_SLICE_X12Y159_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000000000000000)
  ) CLBLM_L_X10Y159_SLICE_X12Y159_BLUT (
.I0(CLBLM_R_X11Y160_SLICE_X14Y160_AQ),
.I1(CLBLM_L_X10Y156_SLICE_X13Y156_CO6),
.I2(CLBLM_R_X11Y156_SLICE_X14Y156_BQ),
.I3(CLBLM_R_X11Y155_SLICE_X14Y155_CQ),
.I4(CLBLM_L_X10Y158_SLICE_X12Y158_BQ),
.I5(CLBLM_R_X11Y159_SLICE_X15Y159_BQ),
.O5(CLBLM_L_X10Y159_SLICE_X12Y159_BO5),
.O6(CLBLM_L_X10Y159_SLICE_X12Y159_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000e4444444)
  ) CLBLM_L_X10Y159_SLICE_X12Y159_ALUT (
.I0(CLBLM_R_X11Y159_SLICE_X14Y159_DQ),
.I1(CLBLM_L_X10Y159_SLICE_X13Y159_BO5),
.I2(CLBLM_R_X11Y160_SLICE_X14Y160_AQ),
.I3(CLBLM_L_X10Y159_SLICE_X13Y159_AO5),
.I4(CLBLM_R_X11Y159_SLICE_X15Y159_BQ),
.I5(CLBLM_L_X8Y156_SLICE_X11Y156_DO6),
.O5(CLBLM_L_X10Y159_SLICE_X12Y159_AO5),
.O6(CLBLM_L_X10Y159_SLICE_X12Y159_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ddfd0000dfff)
  ) CLBLM_L_X10Y159_SLICE_X13Y159_DLUT (
.I0(CLBLM_L_X8Y158_SLICE_X11Y158_AQ),
.I1(CLBLM_L_X8Y156_SLICE_X11Y156_DO6),
.I2(CLBLM_R_X11Y160_SLICE_X14Y160_AQ),
.I3(CLBLM_L_X10Y159_SLICE_X13Y159_AO5),
.I4(CLBLM_L_X8Y157_SLICE_X11Y157_DO6),
.I5(CLBLM_L_X10Y159_SLICE_X13Y159_BO6),
.O5(CLBLM_L_X10Y159_SLICE_X13Y159_DO5),
.O6(CLBLM_L_X10Y159_SLICE_X13Y159_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00fc3f0f00f87)
  ) CLBLM_L_X10Y159_SLICE_X13Y159_CLUT (
.I0(CLBLM_L_X10Y159_SLICE_X13Y159_AO5),
.I1(CLBLM_L_X8Y157_SLICE_X10Y157_BQ),
.I2(CLBLM_R_X11Y160_SLICE_X14Y160_AQ),
.I3(CLBLM_L_X8Y156_SLICE_X11Y156_DO6),
.I4(CLBLM_L_X8Y157_SLICE_X11Y157_DO6),
.I5(CLBLM_L_X10Y159_SLICE_X13Y159_BO6),
.O5(CLBLM_L_X10Y159_SLICE_X13Y159_CO5),
.O6(CLBLM_L_X10Y159_SLICE_X13Y159_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1010101000000010)
  ) CLBLM_L_X10Y159_SLICE_X13Y159_BLUT (
.I0(CLBLM_L_X10Y158_SLICE_X12Y158_BQ),
.I1(CLBLM_R_X11Y155_SLICE_X14Y155_CQ),
.I2(CLBLM_L_X10Y157_SLICE_X12Y157_CO5),
.I3(CLBLM_R_X11Y159_SLICE_X15Y159_BQ),
.I4(CLBLM_R_X11Y160_SLICE_X14Y160_AQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y159_SLICE_X13Y159_BO5),
.O6(CLBLM_L_X10Y159_SLICE_X13Y159_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1098101000880000)
  ) CLBLM_L_X10Y159_SLICE_X13Y159_ALUT (
.I0(CLBLM_L_X10Y158_SLICE_X12Y158_BQ),
.I1(CLBLM_R_X11Y155_SLICE_X14Y155_CQ),
.I2(CLBLM_L_X10Y157_SLICE_X12Y157_CO5),
.I3(CLBLM_L_X10Y156_SLICE_X13Y156_CO6),
.I4(CLBLM_R_X11Y156_SLICE_X14Y156_BQ),
.I5(1'b1),
.O5(CLBLM_L_X10Y159_SLICE_X13Y159_AO5),
.O6(CLBLM_L_X10Y159_SLICE_X13Y159_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y163_SLICE_X12Y163_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y163_SLICE_X12Y163_DO5),
.O6(CLBLM_L_X10Y163_SLICE_X12Y163_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y163_SLICE_X12Y163_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y163_SLICE_X12Y163_CO5),
.O6(CLBLM_L_X10Y163_SLICE_X12Y163_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y163_SLICE_X12Y163_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y163_SLICE_X12Y163_BO5),
.O6(CLBLM_L_X10Y163_SLICE_X12Y163_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y163_SLICE_X12Y163_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y163_SLICE_X12Y163_AO5),
.O6(CLBLM_L_X10Y163_SLICE_X12Y163_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y163_SLICE_X13Y163_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y163_SLICE_X13Y163_DO5),
.O6(CLBLM_L_X10Y163_SLICE_X13Y163_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y163_SLICE_X13Y163_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y163_SLICE_X13Y163_CO5),
.O6(CLBLM_L_X10Y163_SLICE_X13Y163_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y163_SLICE_X13Y163_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y163_SLICE_X13Y163_BO5),
.O6(CLBLM_L_X10Y163_SLICE_X13Y163_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffffffff)
  ) CLBLM_L_X10Y163_SLICE_X13Y163_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X10Y155_SLICE_X13Y155_A5Q),
.O5(CLBLM_L_X10Y163_SLICE_X13Y163_AO5),
.O6(CLBLM_L_X10Y163_SLICE_X13Y163_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y146_SLICE_X16Y146_AO6),
.Q(CLBLM_L_X12Y146_SLICE_X16Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y146_SLICE_X16Y146_BO6),
.Q(CLBLM_L_X12Y146_SLICE_X16Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y146_SLICE_X16Y146_CO6),
.Q(CLBLM_L_X12Y146_SLICE_X16Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y146_SLICE_X16Y146_DO6),
.Q(CLBLM_L_X12Y146_SLICE_X16Y146_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00ff55aa00fa50)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_L_X12Y146_SLICE_X16Y146_DQ),
.I3(CLBLM_L_X8Y146_SLICE_X11Y146_CQ),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.I5(CLBLM_R_X11Y150_SLICE_X14Y150_AQ),
.O5(CLBLM_L_X12Y146_SLICE_X16Y146_DO5),
.O6(CLBLM_L_X12Y146_SLICE_X16Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafefe00005454)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y146_SLICE_X16Y146_CQ),
.I2(CLBLM_L_X12Y146_SLICE_X16Y146_DQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.I5(CLBLM_L_X12Y146_SLICE_X16Y146_AQ),
.O5(CLBLM_L_X12Y146_SLICE_X16Y146_CO5),
.O6(CLBLM_L_X12Y146_SLICE_X16Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0f0c00000f0c)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y146_SLICE_X16Y146_BQ),
.I2(CLBLM_R_X7Y146_SLICE_X8Y146_DO6),
.I3(CLBLM_L_X12Y146_SLICE_X16Y146_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y153_SLICE_X16Y153_AQ),
.O5(CLBLM_L_X12Y146_SLICE_X16Y146_BO5),
.O6(CLBLM_L_X12Y146_SLICE_X16Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00ffcccc00f0)
  ) CLBLM_L_X12Y146_SLICE_X16Y146_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y146_SLICE_X16Y146_BQ),
.I2(CLBLM_L_X12Y146_SLICE_X16Y146_AQ),
.I3(CLBLM_R_X7Y146_SLICE_X9Y146_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y147_SLICE_X13Y147_BQ),
.O5(CLBLM_L_X12Y146_SLICE_X16Y146_AO5),
.O6(CLBLM_L_X12Y146_SLICE_X16Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y146_SLICE_X17Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y146_SLICE_X17Y146_DO5),
.O6(CLBLM_L_X12Y146_SLICE_X17Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y146_SLICE_X17Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y146_SLICE_X17Y146_CO5),
.O6(CLBLM_L_X12Y146_SLICE_X17Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y146_SLICE_X17Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y146_SLICE_X17Y146_BO5),
.O6(CLBLM_L_X12Y146_SLICE_X17Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000a0f0000080c0)
  ) CLBLM_L_X12Y146_SLICE_X17Y146_ALUT (
.I0(CLBLM_R_X11Y146_SLICE_X15Y146_DO5),
.I1(CLBLM_R_X7Y148_SLICE_X9Y148_CO5),
.I2(CLBLM_L_X10Y145_SLICE_X13Y145_CQ),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_BQ),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_BO6),
.I5(CLBLM_R_X7Y146_SLICE_X9Y146_BO6),
.O5(CLBLM_L_X12Y146_SLICE_X17Y146_AO5),
.O6(CLBLM_L_X12Y146_SLICE_X17Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y147_SLICE_X16Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y147_SLICE_X16Y147_AO6),
.Q(CLBLM_L_X12Y147_SLICE_X16Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_L_X12Y147_SLICE_X16Y147_DLUT (
.I0(CLBLM_R_X11Y150_SLICE_X14Y150_AQ),
.I1(CLBLM_L_X10Y147_SLICE_X12Y147_CQ),
.I2(CLBLM_L_X12Y146_SLICE_X16Y146_DQ),
.I3(CLBLM_R_X13Y153_SLICE_X19Y153_CQ),
.I4(CLBLM_L_X12Y153_SLICE_X17Y153_CQ),
.I5(CLBLM_L_X10Y145_SLICE_X12Y145_BQ),
.O5(CLBLM_L_X12Y147_SLICE_X16Y147_DO5),
.O6(CLBLM_L_X12Y147_SLICE_X16Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033003312121111)
  ) CLBLM_L_X12Y147_SLICE_X16Y147_CLUT (
.I0(CLBLM_L_X12Y153_SLICE_X17Y153_CQ),
.I1(CLBLM_L_X12Y147_SLICE_X16Y147_AQ),
.I2(CLBLM_R_X13Y147_SLICE_X18Y147_AO5),
.I3(CLBLM_L_X8Y148_SLICE_X11Y148_B5Q),
.I4(CLBLM_R_X13Y147_SLICE_X18Y147_BO5),
.I5(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.O5(CLBLM_L_X12Y147_SLICE_X16Y147_CO5),
.O6(CLBLM_L_X12Y147_SLICE_X16Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h20002000fbff0400)
  ) CLBLM_L_X12Y147_SLICE_X16Y147_BLUT (
.I0(CLBLM_L_X10Y146_SLICE_X12Y146_C5Q),
.I1(CLBLM_L_X10Y145_SLICE_X13Y145_BQ),
.I2(CLBLM_L_X10Y146_SLICE_X12Y146_CQ),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_CQ),
.I4(CLBLM_R_X11Y150_SLICE_X14Y150_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y147_SLICE_X16Y147_BO5),
.O6(CLBLM_L_X12Y147_SLICE_X16Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00fd31fd31)
  ) CLBLM_L_X12Y147_SLICE_X16Y147_ALUT (
.I0(RIOB33_X105Y141_IOB_X1Y142_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.I3(CLBLM_L_X10Y150_SLICE_X12Y150_A5Q),
.I4(1'b1),
.I5(CLBLM_L_X12Y147_SLICE_X16Y147_CO6),
.O5(CLBLM_L_X12Y147_SLICE_X16Y147_AO5),
.O6(CLBLM_L_X12Y147_SLICE_X16Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c553c3c3caa)
  ) CLBLM_L_X12Y147_SLICE_X17Y147_DLUT (
.I0(CLBLM_R_X13Y147_SLICE_X18Y147_BO6),
.I1(CLBLM_R_X11Y152_SLICE_X14Y152_BQ),
.I2(CLBLM_L_X12Y154_SLICE_X16Y154_A5Q),
.I3(CLBLM_R_X3Y154_SLICE_X2Y154_AO6),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_BO6),
.I5(CLBLM_R_X13Y147_SLICE_X18Y147_DO6),
.O5(CLBLM_L_X12Y147_SLICE_X17Y147_DO5),
.O6(CLBLM_L_X12Y147_SLICE_X17Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffde00120012ffde)
  ) CLBLM_L_X12Y147_SLICE_X17Y147_CLUT (
.I0(CLBLM_R_X13Y147_SLICE_X18Y147_AO6),
.I1(CLBLM_R_X7Y146_SLICE_X8Y146_BO6),
.I2(CLBLM_L_X12Y147_SLICE_X16Y147_BO5),
.I3(CLBLM_R_X3Y154_SLICE_X2Y154_AO6),
.I4(CLBLM_L_X12Y149_SLICE_X16Y149_B5Q),
.I5(CLBLM_L_X10Y149_SLICE_X12Y149_CQ),
.O5(CLBLM_L_X12Y147_SLICE_X17Y147_CO5),
.O6(CLBLM_L_X12Y147_SLICE_X17Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4e4e1b1b4e0f1b0f)
  ) CLBLM_L_X12Y147_SLICE_X17Y147_BLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_BO6),
.I1(CLBLM_L_X12Y147_SLICE_X16Y147_BO6),
.I2(CLBLM_L_X10Y150_SLICE_X13Y150_C5Q),
.I3(CLBLM_R_X7Y148_SLICE_X9Y148_CO5),
.I4(CLBLM_R_X11Y153_SLICE_X15Y153_DQ),
.I5(CLBLM_R_X7Y146_SLICE_X9Y146_BO6),
.O5(CLBLM_L_X12Y147_SLICE_X17Y147_BO5),
.O6(CLBLM_L_X12Y147_SLICE_X17Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996966996696996)
  ) CLBLM_L_X12Y147_SLICE_X17Y147_ALUT (
.I0(CLBLM_L_X12Y147_SLICE_X17Y147_DO6),
.I1(CLBLM_R_X11Y147_SLICE_X15Y147_AO6),
.I2(CLBLM_L_X12Y148_SLICE_X17Y148_DO6),
.I3(CLBLM_L_X12Y147_SLICE_X17Y147_BO6),
.I4(CLBLM_L_X12Y148_SLICE_X16Y148_CO6),
.I5(CLBLM_L_X12Y147_SLICE_X17Y147_CO6),
.O5(CLBLM_L_X12Y147_SLICE_X17Y147_AO5),
.O6(CLBLM_L_X12Y147_SLICE_X17Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3c3c3c3f3c3f3c)
  ) CLBLM_L_X12Y148_SLICE_X16Y148_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y149_SLICE_X19Y149_CQ),
.I2(CLBLM_R_X13Y149_SLICE_X18Y149_AQ),
.I3(CLBLM_L_X12Y147_SLICE_X16Y147_DO6),
.I4(1'b1),
.I5(CLBLM_L_X12Y148_SLICE_X16Y148_BO6),
.O5(CLBLM_L_X12Y148_SLICE_X16Y148_DO5),
.O6(CLBLM_L_X12Y148_SLICE_X16Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055aaff0050afff)
  ) CLBLM_L_X12Y148_SLICE_X16Y148_CLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_BO6),
.I1(1'b1),
.I2(CLBLM_R_X7Y146_SLICE_X9Y146_BO6),
.I3(CLBLM_L_X12Y148_SLICE_X16Y148_AO5),
.I4(CLBLM_L_X8Y148_SLICE_X11Y148_B5Q),
.I5(CLBLM_R_X7Y148_SLICE_X9Y148_CO5),
.O5(CLBLM_L_X12Y148_SLICE_X16Y148_CO5),
.O6(CLBLM_L_X12Y148_SLICE_X16Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffd)
  ) CLBLM_L_X12Y148_SLICE_X16Y148_BLUT (
.I0(CLBLM_L_X12Y149_SLICE_X17Y149_BO5),
.I1(CLBLM_L_X12Y146_SLICE_X16Y146_BQ),
.I2(CLBLM_L_X12Y149_SLICE_X17Y149_AQ),
.I3(CLBLM_L_X10Y145_SLICE_X12Y145_CQ),
.I4(CLBLM_R_X13Y149_SLICE_X18Y149_BQ),
.I5(CLBLM_L_X12Y146_SLICE_X16Y146_CQ),
.O5(CLBLM_L_X12Y148_SLICE_X16Y148_BO5),
.O6(CLBLM_L_X12Y148_SLICE_X16Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff5fff5cccccc6c)
  ) CLBLM_L_X12Y148_SLICE_X16Y148_ALUT (
.I0(CLBLM_L_X10Y146_SLICE_X12Y146_C5Q),
.I1(CLBLM_L_X12Y153_SLICE_X17Y153_CQ),
.I2(CLBLM_L_X10Y145_SLICE_X13Y145_CQ),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_BQ),
.I4(CLBLM_L_X10Y146_SLICE_X12Y146_CQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y148_SLICE_X16Y148_AO5),
.O6(CLBLM_L_X12Y148_SLICE_X16Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44ee44ff00)
  ) CLBLM_L_X12Y148_SLICE_X17Y148_DLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_BO6),
.I1(CLBLM_L_X12Y149_SLICE_X17Y149_CO5),
.I2(1'b1),
.I3(CLBLM_L_X12Y157_SLICE_X17Y157_A5Q),
.I4(CLBLM_R_X7Y146_SLICE_X9Y146_BO6),
.I5(CLBLM_R_X7Y148_SLICE_X9Y148_CO5),
.O5(CLBLM_L_X12Y148_SLICE_X17Y148_DO5),
.O6(CLBLM_L_X12Y148_SLICE_X17Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000a000b000f000f)
  ) CLBLM_L_X12Y148_SLICE_X17Y148_CLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_BO6),
.I1(CLBLM_R_X7Y148_SLICE_X9Y148_CO5),
.I2(CLBLM_R_X7Y153_SLICE_X8Y153_DO6),
.I3(CLBLM_R_X13Y152_SLICE_X18Y152_DO6),
.I4(CLBLM_R_X7Y146_SLICE_X9Y146_BO6),
.I5(CLBLM_L_X12Y146_SLICE_X16Y146_BQ),
.O5(CLBLM_L_X12Y148_SLICE_X17Y148_CO5),
.O6(CLBLM_L_X12Y148_SLICE_X17Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555455005504)
  ) CLBLM_L_X12Y148_SLICE_X17Y148_BLUT (
.I0(CLBLM_R_X13Y148_SLICE_X18Y148_AO5),
.I1(CLBLM_L_X12Y149_SLICE_X17Y149_CO5),
.I2(CLBLM_R_X3Y154_SLICE_X2Y154_AO6),
.I3(CLBLM_L_X12Y150_SLICE_X17Y150_BQ),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_BO6),
.I5(CLBLM_L_X12Y157_SLICE_X17Y157_A5Q),
.O5(CLBLM_L_X12Y148_SLICE_X17Y148_BO5),
.O6(CLBLM_L_X12Y148_SLICE_X17Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000050505554)
  ) CLBLM_L_X12Y148_SLICE_X17Y148_ALUT (
.I0(CLBLM_R_X13Y149_SLICE_X19Y149_A5Q),
.I1(CLBLM_R_X11Y148_SLICE_X15Y148_CO6),
.I2(CLBLM_R_X13Y149_SLICE_X18Y149_A5Q),
.I3(CLBLM_L_X12Y148_SLICE_X17Y148_BO6),
.I4(CLBLM_R_X11Y148_SLICE_X15Y148_DO6),
.I5(CLBLM_L_X12Y148_SLICE_X17Y148_CO6),
.O5(CLBLM_L_X12Y148_SLICE_X17Y148_AO5),
.O6(CLBLM_L_X12Y148_SLICE_X17Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y149_SLICE_X16Y149_BO5),
.Q(CLBLM_L_X12Y149_SLICE_X16Y149_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y149_SLICE_X16Y149_AO6),
.Q(CLBLM_L_X12Y149_SLICE_X16Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y149_SLICE_X16Y149_BO6),
.Q(CLBLM_L_X12Y149_SLICE_X16Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y149_SLICE_X16Y149_CO6),
.Q(CLBLM_L_X12Y149_SLICE_X16Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y149_SLICE_X16Y149_DO6),
.Q(CLBLM_L_X12Y149_SLICE_X16Y149_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aa00ee44)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y151_SLICE_X16Y151_BQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y144_SLICE_X15Y144_A5Q),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X11Y151_SLICE_X15Y151_CO6),
.O5(CLBLM_L_X12Y149_SLICE_X16Y149_DO5),
.O6(CLBLM_L_X12Y149_SLICE_X16Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000aaea0040)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y151_SLICE_X16Y151_BQ),
.I2(CLBLM_L_X12Y150_SLICE_X16Y150_BQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y146_SLICE_X14Y146_BQ),
.I5(CLBLM_R_X11Y151_SLICE_X15Y151_CO6),
.O5(CLBLM_L_X12Y149_SLICE_X16Y149_CO5),
.O6(CLBLM_L_X12Y149_SLICE_X16Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfc0cfc0fafa0a0a)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_BLUT (
.I0(CLBLM_L_X12Y150_SLICE_X16Y150_A5Q),
.I1(CLBLM_R_X13Y149_SLICE_X18Y149_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(CLBLM_R_X5Y149_SLICE_X7Y149_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y149_SLICE_X16Y149_BO5),
.O6(CLBLM_L_X12Y149_SLICE_X16Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc00ee22ec20)
  ) CLBLM_L_X12Y149_SLICE_X16Y149_ALUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y149_SLICE_X16Y149_AQ),
.I3(CLBLM_L_X12Y150_SLICE_X16Y150_BQ),
.I4(CLBLM_L_X12Y147_SLICE_X16Y147_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X12Y149_SLICE_X16Y149_AO5),
.O6(CLBLM_L_X12Y149_SLICE_X16Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y149_SLICE_X17Y149_BO6),
.Q(CLBLM_L_X12Y149_SLICE_X17Y149_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X12Y149_SLICE_X17Y149_AO6),
.Q(CLBLM_L_X12Y149_SLICE_X17Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f2f0f2f0f0f0fa)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_DLUT (
.I0(CLBLM_L_X12Y146_SLICE_X17Y146_AO6),
.I1(CLBLM_L_X12Y157_SLICE_X17Y157_A5Q),
.I2(CLBLM_R_X13Y149_SLICE_X19Y149_AQ),
.I3(CLBLM_R_X11Y155_SLICE_X15Y155_BO6),
.I4(CLBLM_L_X12Y149_SLICE_X17Y149_CO5),
.I5(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.O5(CLBLM_L_X12Y149_SLICE_X17Y149_DO5),
.O6(CLBLM_L_X12Y149_SLICE_X17Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfffcffaaa6aaaa)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_CLUT (
.I0(CLBLM_L_X10Y145_SLICE_X12Y145_BQ),
.I1(CLBLM_L_X10Y145_SLICE_X13Y145_CQ),
.I2(CLBLM_L_X10Y146_SLICE_X12Y146_C5Q),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_BQ),
.I4(CLBLM_L_X10Y146_SLICE_X12Y146_CQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y149_SLICE_X17Y149_CO5),
.O6(CLBLM_L_X12Y149_SLICE_X17Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f000ee11111111)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_BLUT (
.I0(CLBLM_R_X11Y153_SLICE_X15Y153_DQ),
.I1(CLBLM_L_X12Y149_SLICE_X17Y149_A5Q),
.I2(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y149_SLICE_X17Y149_BO5),
.O6(CLBLM_L_X12Y149_SLICE_X17Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aafcaa00aafc)
  ) CLBLM_L_X12Y149_SLICE_X17Y149_ALUT (
.I0(CLBLM_L_X12Y157_SLICE_X17Y157_CQ),
.I1(CLBLM_L_X12Y146_SLICE_X16Y146_BQ),
.I2(CLBLM_L_X12Y149_SLICE_X17Y149_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_DO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y149_SLICE_X17Y149_AO5),
.O6(CLBLM_L_X12Y149_SLICE_X17Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y150_SLICE_X16Y150_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y154_SLICE_X15Y154_CO6),
.Q(CLBLM_L_X12Y150_SLICE_X16Y150_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y150_SLICE_X16Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y150_SLICE_X16Y150_AO6),
.Q(CLBLM_L_X12Y150_SLICE_X16Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y150_SLICE_X16Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y150_SLICE_X16Y150_BO6),
.Q(CLBLM_L_X12Y150_SLICE_X16Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y150_SLICE_X16Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y150_SLICE_X16Y150_CO6),
.Q(CLBLM_L_X12Y150_SLICE_X16Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f1100000fee)
  ) CLBLM_L_X12Y150_SLICE_X16Y150_DLUT (
.I0(CLBLM_L_X10Y146_SLICE_X12Y146_CQ),
.I1(CLBLM_L_X12Y149_SLICE_X17Y149_CO6),
.I2(CLBLM_L_X8Y155_SLICE_X10Y155_BQ),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.I4(CLBLM_L_X12Y150_SLICE_X16Y150_CQ),
.I5(CLBLM_L_X12Y149_SLICE_X17Y149_A5Q),
.O5(CLBLM_L_X12Y150_SLICE_X16Y150_DO5),
.O6(CLBLM_L_X12Y150_SLICE_X16Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00fd31cc00fd31)
  ) CLBLM_L_X12Y150_SLICE_X16Y150_CLUT (
.I0(RIOB33_X105Y141_IOB_X1Y142_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.I3(CLBLM_L_X8Y153_SLICE_X11Y153_CQ),
.I4(CLBLM_L_X12Y150_SLICE_X16Y150_DO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y150_SLICE_X16Y150_CO5),
.O6(CLBLM_L_X12Y150_SLICE_X16Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0faa00aa0caa00)
  ) CLBLM_L_X12Y150_SLICE_X16Y150_BLUT (
.I0(CLBLM_L_X12Y152_SLICE_X16Y152_CQ),
.I1(CLBLM_L_X12Y150_SLICE_X16Y150_BQ),
.I2(CLBLM_L_X12Y149_SLICE_X16Y149_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X12Y149_SLICE_X16Y149_DQ),
.O5(CLBLM_L_X12Y150_SLICE_X16Y150_BO5),
.O6(CLBLM_L_X12Y150_SLICE_X16Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccf0ccaacca0)
  ) CLBLM_L_X12Y150_SLICE_X16Y150_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X13Y149_SLICE_X18Y149_BQ),
.I2(CLBLM_L_X12Y150_SLICE_X16Y150_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y150_SLICE_X9Y150_BO6),
.I5(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.O5(CLBLM_L_X12Y150_SLICE_X16Y150_AO5),
.O6(CLBLM_L_X12Y150_SLICE_X16Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y150_SLICE_X17Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y150_SLICE_X17Y150_AO6),
.Q(CLBLM_L_X12Y150_SLICE_X17Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y150_SLICE_X17Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y150_SLICE_X17Y150_BO6),
.Q(CLBLM_L_X12Y150_SLICE_X17Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000505f5c53)
  ) CLBLM_L_X12Y150_SLICE_X17Y150_DLUT (
.I0(CLBLM_R_X11Y152_SLICE_X14Y152_BQ),
.I1(CLBLM_L_X10Y146_SLICE_X12Y146_CQ),
.I2(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.I3(CLBLM_L_X12Y146_SLICE_X16Y146_DQ),
.I4(CLBLM_L_X12Y149_SLICE_X17Y149_CO6),
.I5(CLBLM_R_X13Y150_SLICE_X18Y150_CQ),
.O5(CLBLM_L_X12Y150_SLICE_X17Y150_DO5),
.O6(CLBLM_L_X12Y150_SLICE_X17Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0213130202130213)
  ) CLBLM_L_X12Y150_SLICE_X17Y150_CLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.I1(CLBLM_L_X12Y155_SLICE_X17Y155_CQ),
.I2(CLBLM_L_X12Y154_SLICE_X16Y154_A5Q),
.I3(CLBLM_R_X13Y153_SLICE_X19Y153_CQ),
.I4(CLBLM_L_X12Y148_SLICE_X16Y148_AO6),
.I5(CLBLM_L_X10Y146_SLICE_X12Y146_CQ),
.O5(CLBLM_L_X12Y150_SLICE_X17Y150_CO5),
.O6(CLBLM_L_X12Y150_SLICE_X17Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000af8caf8c)
  ) CLBLM_L_X12Y150_SLICE_X17Y150_BLUT (
.I0(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.I1(CLBLM_L_X12Y150_SLICE_X17Y150_BQ),
.I2(RIOB33_X105Y141_IOB_X1Y142_I),
.I3(CLBLM_L_X12Y148_SLICE_X17Y148_DO6),
.I4(CLBLM_R_X7Y149_SLICE_X9Y149_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y150_SLICE_X17Y150_BO5),
.O6(CLBLM_L_X12Y150_SLICE_X17Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000033723372)
  ) CLBLM_L_X12Y150_SLICE_X17Y150_ALUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I1(CLBLM_L_X10Y150_SLICE_X12Y150_BO6),
.I2(CLBLM_L_X12Y150_SLICE_X17Y150_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X12Y154_SLICE_X17Y154_DQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y150_SLICE_X17Y150_AO5),
.O6(CLBLM_L_X12Y150_SLICE_X17Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y151_SLICE_X16Y151_CO5),
.Q(CLBLM_L_X12Y151_SLICE_X16Y151_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y151_SLICE_X16Y151_AO6),
.Q(CLBLM_L_X12Y151_SLICE_X16Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y151_SLICE_X16Y151_BO6),
.Q(CLBLM_L_X12Y151_SLICE_X16Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y151_SLICE_X16Y151_CO6),
.Q(CLBLM_L_X12Y151_SLICE_X16Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff6f6f6f6)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_DLUT (
.I0(CLBLM_R_X13Y150_SLICE_X19Y150_AQ),
.I1(CLBLM_L_X12Y153_SLICE_X16Y153_AQ),
.I2(CLBLM_R_X11Y150_SLICE_X15Y150_DO6),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X11Y151_SLICE_X14Y151_DO6),
.O5(CLBLM_L_X12Y151_SLICE_X16Y151_DO5),
.O6(CLBLM_L_X12Y151_SLICE_X16Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8b8b8ff33cc00)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_CLUT (
.I0(CLBLM_R_X13Y153_SLICE_X18Y153_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(CLBLM_L_X12Y150_SLICE_X17Y150_BQ),
.I4(CLBLM_R_X11Y151_SLICE_X15Y151_A5Q),
.I5(1'b1),
.O5(CLBLM_L_X12Y151_SLICE_X16Y151_CO5),
.O6(CLBLM_L_X12Y151_SLICE_X16Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaabbeea00011440)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y151_SLICE_X16Y151_BQ),
.I2(CLBLM_L_X12Y151_SLICE_X17Y151_DO6),
.I3(CLBLM_L_X12Y152_SLICE_X16Y152_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X10Y154_SLICE_X13Y154_C5Q),
.O5(CLBLM_L_X12Y151_SLICE_X16Y151_BO5),
.O6(CLBLM_L_X12Y151_SLICE_X16Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffeccdc33320010)
  ) CLBLM_L_X12Y151_SLICE_X16Y151_ALUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y151_SLICE_X16Y151_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_L_X12Y149_SLICE_X16Y149_AQ),
.I5(CLBLM_R_X11Y157_SLICE_X14Y157_BQ),
.O5(CLBLM_L_X12Y151_SLICE_X16Y151_AO5),
.O6(CLBLM_L_X12Y151_SLICE_X16Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y151_SLICE_X17Y151_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y151_SLICE_X17Y151_AO5),
.Q(CLBLM_L_X12Y151_SLICE_X17Y151_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y151_SLICE_X17Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y151_SLICE_X17Y151_AO6),
.Q(CLBLM_L_X12Y151_SLICE_X17Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y151_SLICE_X17Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y151_SLICE_X17Y151_BO6),
.Q(CLBLM_L_X12Y151_SLICE_X17Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc33cc33dd22dd22)
  ) CLBLM_L_X12Y151_SLICE_X17Y151_DLUT (
.I0(CLBLM_R_X11Y151_SLICE_X15Y151_CO6),
.I1(CLBLM_L_X10Y154_SLICE_X13Y154_BQ),
.I2(1'b1),
.I3(CLBLM_L_X12Y151_SLICE_X17Y151_BQ),
.I4(1'b1),
.I5(CLBLM_L_X12Y151_SLICE_X16Y151_BQ),
.O5(CLBLM_L_X12Y151_SLICE_X17Y151_DO5),
.O6(CLBLM_L_X12Y151_SLICE_X17Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6f6f6f6ff6f6f6f6)
  ) CLBLM_L_X12Y151_SLICE_X17Y151_CLUT (
.I0(CLBLM_R_X11Y149_SLICE_X14Y149_BQ),
.I1(CLBLM_R_X13Y153_SLICE_X19Y153_AQ),
.I2(CLBLM_R_X13Y151_SLICE_X18Y151_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X12Y151_SLICE_X16Y151_AQ),
.O5(CLBLM_L_X12Y151_SLICE_X17Y151_CO5),
.O6(CLBLM_L_X12Y151_SLICE_X17Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0c0c00000c0c)
  ) CLBLM_L_X12Y151_SLICE_X17Y151_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y152_SLICE_X16Y152_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y154_SLICE_X16Y154_A5Q),
.O5(CLBLM_L_X12Y151_SLICE_X17Y151_BO5),
.O6(CLBLM_L_X12Y151_SLICE_X17Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aacccc00ccf0)
  ) CLBLM_L_X12Y151_SLICE_X17Y151_ALUT (
.I0(CLBLM_L_X12Y155_SLICE_X17Y155_CQ),
.I1(CLBLM_L_X12Y151_SLICE_X17Y151_BQ),
.I2(CLBLM_R_X5Y152_SLICE_X6Y152_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y151_SLICE_X17Y151_AO5),
.O6(CLBLM_L_X12Y151_SLICE_X17Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y152_SLICE_X16Y152_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y153_SLICE_X17Y153_DO6),
.Q(CLBLM_L_X12Y152_SLICE_X16Y152_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y152_SLICE_X16Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y152_SLICE_X16Y152_AO6),
.Q(CLBLM_L_X12Y152_SLICE_X16Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y152_SLICE_X16Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y152_SLICE_X16Y152_BO6),
.Q(CLBLM_L_X12Y152_SLICE_X16Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y152_SLICE_X16Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y152_SLICE_X16Y152_CO6),
.Q(CLBLM_L_X12Y152_SLICE_X16Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000f00000003000f)
  ) CLBLM_L_X12Y152_SLICE_X16Y152_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y155_SLICE_X16Y155_AO5),
.I2(CLBLM_L_X12Y152_SLICE_X17Y152_DO6),
.I3(CLBLM_L_X12Y151_SLICE_X16Y151_DO6),
.I4(CLBLM_R_X7Y154_SLICE_X9Y154_DO6),
.I5(CLBLM_R_X13Y152_SLICE_X19Y152_CO6),
.O5(CLBLM_L_X12Y152_SLICE_X16Y152_DO5),
.O6(CLBLM_L_X12Y152_SLICE_X16Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffc8ff00ffc8)
  ) CLBLM_L_X12Y152_SLICE_X16Y152_CLUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I1(CLBLM_L_X12Y152_SLICE_X16Y152_CQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_L_X8Y152_SLICE_X11Y152_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X13Y156_SLICE_X18Y156_AQ),
.O5(CLBLM_L_X12Y152_SLICE_X16Y152_CO5),
.O6(CLBLM_L_X12Y152_SLICE_X16Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44aa00aa00)
  ) CLBLM_L_X12Y152_SLICE_X16Y152_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y150_SLICE_X13Y150_AQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y152_SLICE_X15Y152_AQ),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X12Y152_SLICE_X16Y152_BO5),
.O6(CLBLM_L_X12Y152_SLICE_X16Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8b8b8880f0f0fff)
  ) CLBLM_L_X12Y152_SLICE_X16Y152_ALUT (
.I0(CLBLM_R_X11Y152_SLICE_X15Y152_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X12Y152_SLICE_X16Y152_CQ),
.I4(CLBLM_R_X5Y151_SLICE_X6Y151_CQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y152_SLICE_X16Y152_AO5),
.O6(CLBLM_L_X12Y152_SLICE_X16Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y152_SLICE_X17Y152_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y152_SLICE_X17Y152_BO6),
.Q(CLBLM_L_X12Y152_SLICE_X17Y152_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y152_SLICE_X17Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y152_SLICE_X17Y152_AO6),
.Q(CLBLM_L_X12Y152_SLICE_X17Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hddeeffffffffddee)
  ) CLBLM_L_X12Y152_SLICE_X17Y152_DLUT (
.I0(CLBLM_R_X13Y153_SLICE_X18Y153_AQ),
.I1(CLBLM_L_X12Y151_SLICE_X17Y151_CO6),
.I2(1'b1),
.I3(CLBLM_R_X11Y153_SLICE_X15Y153_CQ),
.I4(CLBLM_R_X11Y152_SLICE_X15Y152_CQ),
.I5(CLBLM_L_X10Y153_SLICE_X13Y153_AQ),
.O5(CLBLM_L_X12Y152_SLICE_X17Y152_DO5),
.O6(CLBLM_L_X12Y152_SLICE_X17Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_L_X12Y152_SLICE_X17Y152_CLUT (
.I0(CLBLM_R_X13Y151_SLICE_X18Y151_BQ),
.I1(CLBLM_R_X11Y153_SLICE_X15Y153_CQ),
.I2(CLBLM_R_X11Y152_SLICE_X15Y152_CQ),
.I3(CLBLM_R_X11Y152_SLICE_X15Y152_BQ),
.I4(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I5(CLBLM_L_X12Y153_SLICE_X17Y153_BQ),
.O5(CLBLM_L_X12Y152_SLICE_X17Y152_CO5),
.O6(CLBLM_L_X12Y152_SLICE_X17Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0cca0f0f0a0a0)
  ) CLBLM_L_X12Y152_SLICE_X17Y152_BLUT (
.I0(CLBLM_L_X12Y151_SLICE_X17Y151_AQ),
.I1(CLBLL_L_X4Y147_SLICE_X5Y147_AQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y152_SLICE_X14Y152_CQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y152_SLICE_X17Y152_BO5),
.O6(CLBLM_L_X12Y152_SLICE_X17Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0fcc0fcc00cc00)
  ) CLBLM_L_X12Y152_SLICE_X17Y152_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y152_SLICE_X18Y152_AQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y151_SLICE_X8Y151_DQ),
.O5(CLBLM_L_X12Y152_SLICE_X17Y152_AO5),
.O6(CLBLM_L_X12Y152_SLICE_X17Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y153_SLICE_X16Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y153_SLICE_X16Y153_AO6),
.Q(CLBLM_L_X12Y153_SLICE_X16Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffb)
  ) CLBLM_L_X12Y153_SLICE_X16Y153_DLUT (
.I0(CLBLM_L_X10Y155_SLICE_X12Y155_AQ),
.I1(CLBLM_R_X13Y153_SLICE_X18Y153_CQ),
.I2(CLBLM_L_X12Y153_SLICE_X17Y153_CQ),
.I3(CLBLM_L_X12Y153_SLICE_X16Y153_CO6),
.I4(CLBLM_R_X7Y152_SLICE_X9Y152_AQ),
.I5(CLBLM_R_X13Y149_SLICE_X18Y149_A5Q),
.O5(CLBLM_L_X12Y153_SLICE_X16Y153_DO5),
.O6(CLBLM_L_X12Y153_SLICE_X16Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbfffafffb3ffa0ff)
  ) CLBLM_L_X12Y153_SLICE_X16Y153_CLUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(CLBLM_L_X8Y153_SLICE_X10Y153_A5Q),
.I4(RIOB33_X105Y141_IOB_X1Y142_I),
.I5(RIOB33_X105Y127_IOB_X1Y128_I),
.O5(CLBLM_L_X12Y153_SLICE_X16Y153_CO5),
.O6(CLBLM_L_X12Y153_SLICE_X16Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50ea40f0f0c0c0)
  ) CLBLM_L_X12Y153_SLICE_X16Y153_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y151_SLICE_X8Y151_DQ),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X12Y153_SLICE_X17Y153_BQ),
.I4(CLBLM_L_X8Y149_SLICE_X11Y149_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y153_SLICE_X16Y153_BO5),
.O6(CLBLM_L_X12Y153_SLICE_X16Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc0ffaa00c000aa)
  ) CLBLM_L_X12Y153_SLICE_X16Y153_ALUT (
.I0(CLBLM_R_X11Y153_SLICE_X15Y153_CQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X12Y153_SLICE_X16Y153_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y149_SLICE_X15Y149_DO6),
.I5(CLBLL_L_X4Y153_SLICE_X5Y153_AQ),
.O5(CLBLM_L_X12Y153_SLICE_X16Y153_AO5),
.O6(CLBLM_L_X12Y153_SLICE_X16Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y153_SLICE_X17Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y153_SLICE_X17Y153_AO6),
.Q(CLBLM_L_X12Y153_SLICE_X17Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y153_SLICE_X17Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y153_SLICE_X17Y153_BO6),
.Q(CLBLM_L_X12Y153_SLICE_X17Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y153_SLICE_X17Y153_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y153_SLICE_X17Y153_CO6),
.Q(CLBLM_L_X12Y153_SLICE_X17Y153_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaca0a0ffcc0000)
  ) CLBLM_L_X12Y153_SLICE_X17Y153_DLUT (
.I0(CLBLM_R_X13Y150_SLICE_X18Y150_CQ),
.I1(CLBLM_L_X10Y158_SLICE_X13Y158_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X13Y153_SLICE_X18Y153_DQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y153_SLICE_X17Y153_DO5),
.O6(CLBLM_L_X12Y153_SLICE_X17Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0055554444)
  ) CLBLM_L_X12Y153_SLICE_X17Y153_CLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.I1(CLBLM_L_X10Y145_SLICE_X12Y145_CQ),
.I2(1'b1),
.I3(CLBLM_R_X13Y153_SLICE_X18Y153_DQ),
.I4(CLBLM_L_X12Y153_SLICE_X17Y153_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y153_SLICE_X17Y153_CO5),
.O6(CLBLM_L_X12Y153_SLICE_X17Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00caca0a0a)
  ) CLBLM_L_X12Y153_SLICE_X17Y153_BLUT (
.I0(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I1(CLBLM_L_X12Y153_SLICE_X17Y153_BQ),
.I2(CLBLM_R_X11Y149_SLICE_X15Y149_DO6),
.I3(CLBLM_L_X10Y157_SLICE_X12Y157_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y153_SLICE_X17Y153_BO5),
.O6(CLBLM_L_X12Y153_SLICE_X17Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffcccfcffecccec)
  ) CLBLM_L_X12Y153_SLICE_X17Y153_ALUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I1(CLBLM_L_X10Y152_SLICE_X12Y152_DO6),
.I2(CLBLM_L_X12Y153_SLICE_X17Y153_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y150_SLICE_X5Y150_D5Q),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_L_X12Y153_SLICE_X17Y153_AO5),
.O6(CLBLM_L_X12Y153_SLICE_X17Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y154_SLICE_X16Y154_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y154_SLICE_X16Y154_CO6),
.Q(CLBLM_L_X12Y154_SLICE_X16Y154_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y154_SLICE_X16Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y154_SLICE_X16Y154_AO6),
.Q(CLBLM_L_X12Y154_SLICE_X16Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y154_SLICE_X16Y154_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y154_SLICE_X16Y154_BO6),
.Q(CLBLM_L_X12Y154_SLICE_X16Y154_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h15550000efafffff)
  ) CLBLM_L_X12Y154_SLICE_X16Y154_DLUT (
.I0(CLBLM_R_X11Y149_SLICE_X15Y149_DO6),
.I1(CLBLM_L_X12Y154_SLICE_X16Y154_AQ),
.I2(CLBLM_R_X11Y154_SLICE_X15Y154_BQ),
.I3(CLBLM_L_X12Y154_SLICE_X16Y154_BQ),
.I4(CLBLM_R_X13Y155_SLICE_X18Y155_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y154_SLICE_X16Y154_DO5),
.O6(CLBLM_L_X12Y154_SLICE_X16Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaa03000300)
  ) CLBLM_L_X12Y154_SLICE_X16Y154_CLUT (
.I0(CLBLM_L_X12Y152_SLICE_X16Y152_AQ),
.I1(CLBLM_L_X12Y154_SLICE_X17Y154_A5Q),
.I2(CLBLM_L_X12Y155_SLICE_X17Y155_AQ),
.I3(CLBLM_L_X8Y153_SLICE_X11Y153_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y154_SLICE_X16Y154_CO5),
.O6(CLBLM_L_X12Y154_SLICE_X16Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaa0acccc00aa)
  ) CLBLM_L_X12Y154_SLICE_X16Y154_BLUT (
.I0(CLBLM_L_X10Y154_SLICE_X12Y154_BO5),
.I1(CLBLM_R_X7Y152_SLICE_X8Y152_A5Q),
.I2(CLBLM_R_X13Y155_SLICE_X18Y155_AQ),
.I3(CLBLM_L_X12Y154_SLICE_X16Y154_DO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y154_SLICE_X16Y154_BQ),
.O5(CLBLM_L_X12Y154_SLICE_X16Y154_BO5),
.O6(CLBLM_L_X12Y154_SLICE_X16Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccca0aacccca0a0)
  ) CLBLM_L_X12Y154_SLICE_X16Y154_ALUT (
.I0(CLBLM_L_X10Y154_SLICE_X12Y154_BO5),
.I1(CLBLM_R_X13Y154_SLICE_X18Y154_BQ),
.I2(CLBLM_L_X12Y154_SLICE_X16Y154_AQ),
.I3(CLBLM_L_X12Y154_SLICE_X16Y154_DO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y154_SLICE_X16Y154_BQ),
.O5(CLBLM_L_X12Y154_SLICE_X16Y154_AO5),
.O6(CLBLM_L_X12Y154_SLICE_X16Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y154_SLICE_X17Y154_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y154_SLICE_X17Y154_CO6),
.Q(CLBLM_L_X12Y154_SLICE_X17Y154_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y154_SLICE_X17Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y154_SLICE_X17Y154_AO6),
.Q(CLBLM_L_X12Y154_SLICE_X17Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y154_SLICE_X17Y154_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y154_SLICE_X17Y154_BO6),
.Q(CLBLM_L_X12Y154_SLICE_X17Y154_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y154_SLICE_X17Y154_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y154_SLICE_X17Y154_DO6),
.Q(CLBLM_L_X12Y154_SLICE_X17Y154_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaaf0ffffaac0)
  ) CLBLM_L_X12Y154_SLICE_X17Y154_DLUT (
.I0(CLBLM_L_X12Y157_SLICE_X16Y157_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_L_X12Y154_SLICE_X17Y154_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y148_SLICE_X12Y148_DO6),
.I5(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.O5(CLBLM_L_X12Y154_SLICE_X17Y154_DO5),
.O6(CLBLM_L_X12Y154_SLICE_X17Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa3ac00cc00cc)
  ) CLBLM_L_X12Y154_SLICE_X17Y154_CLUT (
.I0(CLBLM_R_X13Y152_SLICE_X18Y152_A5Q),
.I1(CLBLM_L_X8Y153_SLICE_X11Y153_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y154_SLICE_X17Y154_A5Q),
.I4(CLBLM_R_X11Y158_SLICE_X15Y158_BO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y154_SLICE_X17Y154_CO5),
.O6(CLBLM_L_X12Y154_SLICE_X17Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff140014ff040004)
  ) CLBLM_L_X12Y154_SLICE_X17Y154_BLUT (
.I0(CLBLM_R_X11Y158_SLICE_X15Y158_BO6),
.I1(CLBLM_L_X12Y154_SLICE_X17Y154_BQ),
.I2(CLBLM_L_X12Y154_SLICE_X16Y154_CO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X13Y152_SLICE_X18Y152_CQ),
.I5(CLBLM_R_X11Y155_SLICE_X15Y155_AQ),
.O5(CLBLM_L_X12Y154_SLICE_X17Y154_BO5),
.O6(CLBLM_L_X12Y154_SLICE_X17Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00fffff700f7)
  ) CLBLM_L_X12Y154_SLICE_X17Y154_ALUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLL_L_X4Y158_SLICE_X4Y158_AO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y154_SLICE_X13Y154_AQ),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLM_L_X12Y154_SLICE_X17Y154_AO5),
.O6(CLBLM_L_X12Y154_SLICE_X17Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y155_SLICE_X16Y155_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X12Y151_SLICE_X16Y151_CQ),
.Q(CLBLM_L_X12Y155_SLICE_X16Y155_AQ),
.R(CLBLM_R_X13Y155_SLICE_X18Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aa9a00000000)
  ) CLBLM_L_X12Y155_SLICE_X16Y155_DLUT (
.I0(CLBLM_R_X11Y154_SLICE_X15Y154_BQ),
.I1(CLBLM_R_X11Y149_SLICE_X15Y149_DO6),
.I2(CLBLM_R_X13Y155_SLICE_X18Y155_AQ),
.I3(CLBLM_L_X12Y155_SLICE_X16Y155_AO5),
.I4(CLBLM_R_X7Y153_SLICE_X8Y153_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_L_X12Y155_SLICE_X16Y155_DO5),
.O6(CLBLM_L_X12Y155_SLICE_X16Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff7fffffff)
  ) CLBLM_L_X12Y155_SLICE_X16Y155_CLUT (
.I0(CLBLM_L_X12Y154_SLICE_X16Y154_BQ),
.I1(CLBLM_R_X11Y154_SLICE_X15Y154_BQ),
.I2(CLBLM_R_X13Y155_SLICE_X18Y155_AQ),
.I3(CLBLM_L_X12Y154_SLICE_X16Y154_AQ),
.I4(CLBLM_R_X11Y149_SLICE_X15Y149_DO6),
.I5(CLBLM_L_X12Y152_SLICE_X16Y152_DO6),
.O5(CLBLM_L_X12Y155_SLICE_X16Y155_CO5),
.O6(CLBLM_L_X12Y155_SLICE_X16Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000030000000100)
  ) CLBLM_L_X12Y155_SLICE_X16Y155_BLUT (
.I0(CLBLM_R_X11Y155_SLICE_X15Y155_AQ),
.I1(CLBLM_L_X12Y154_SLICE_X17Y154_BQ),
.I2(CLBLM_L_X12Y154_SLICE_X17Y154_A5Q),
.I3(CLBLM_L_X8Y153_SLICE_X11Y153_BQ),
.I4(CLBLM_L_X12Y155_SLICE_X17Y155_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y155_SLICE_X16Y155_BO5),
.O6(CLBLM_L_X12Y155_SLICE_X16Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heaaaaaaac0000000)
  ) CLBLM_L_X12Y155_SLICE_X16Y155_ALUT (
.I0(CLBLM_R_X11Y149_SLICE_X15Y149_DO6),
.I1(CLBLM_R_X11Y154_SLICE_X15Y154_BQ),
.I2(CLBLM_R_X13Y155_SLICE_X18Y155_AQ),
.I3(CLBLM_L_X12Y154_SLICE_X16Y154_AQ),
.I4(CLBLM_L_X12Y154_SLICE_X16Y154_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y155_SLICE_X16Y155_AO5),
.O6(CLBLM_L_X12Y155_SLICE_X16Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y155_SLICE_X17Y155_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y155_SLICE_X17Y155_AO6),
.Q(CLBLM_L_X12Y155_SLICE_X17Y155_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y155_SLICE_X17Y155_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y155_SLICE_X17Y155_BO6),
.Q(CLBLM_L_X12Y155_SLICE_X17Y155_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y155_SLICE_X17Y155_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y155_SLICE_X17Y155_CO6),
.Q(CLBLM_L_X12Y155_SLICE_X17Y155_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffcc0000fafa)
  ) CLBLM_L_X12Y155_SLICE_X17Y155_DLUT (
.I0(CLBLM_R_X7Y154_SLICE_X8Y154_AQ),
.I1(CLBLM_R_X11Y155_SLICE_X14Y155_DQ),
.I2(CLBLM_L_X12Y154_SLICE_X17Y154_DQ),
.I3(CLBLM_L_X10Y148_SLICE_X13Y148_CQ),
.I4(CLBLM_L_X10Y150_SLICE_X13Y150_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y155_SLICE_X17Y155_DO5),
.O6(CLBLM_L_X12Y155_SLICE_X17Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff000000afaf)
  ) CLBLM_L_X12Y155_SLICE_X17Y155_CLUT (
.I0(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.I1(1'b1),
.I2(RIOB33_X105Y141_IOB_X1Y142_I),
.I3(CLBLM_L_X8Y156_SLICE_X10Y156_BQ),
.I4(CLBLM_L_X12Y150_SLICE_X17Y150_CO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y155_SLICE_X17Y155_CO5),
.O6(CLBLM_L_X12Y155_SLICE_X17Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aafcaa00aa00)
  ) CLBLM_L_X12Y155_SLICE_X17Y155_BLUT (
.I0(CLBLM_R_X11Y156_SLICE_X14Y156_AQ),
.I1(CLBLM_L_X12Y155_SLICE_X17Y155_BQ),
.I2(CLBLM_L_X12Y155_SLICE_X17Y155_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.O5(CLBLM_L_X12Y155_SLICE_X17Y155_BO5),
.O6(CLBLM_L_X12Y155_SLICE_X17Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000cddc0110)
  ) CLBLM_L_X12Y155_SLICE_X17Y155_ALUT (
.I0(CLBLM_R_X11Y158_SLICE_X15Y158_BO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y155_SLICE_X17Y155_AQ),
.I3(CLBLM_L_X12Y154_SLICE_X17Y154_CO5),
.I4(CLBLM_L_X12Y155_SLICE_X16Y155_AQ),
.I5(CLBLM_L_X12Y155_SLICE_X16Y155_BO5),
.O5(CLBLM_L_X12Y155_SLICE_X17Y155_AO5),
.O6(CLBLM_L_X12Y155_SLICE_X17Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y156_SLICE_X16Y156_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X7Y155_SLICE_X8Y155_AQ),
.Q(CLBLM_L_X12Y156_SLICE_X16Y156_AQ),
.R(CLBLM_R_X13Y155_SLICE_X18Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y156_SLICE_X16Y156_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X11Y146_SLICE_X15Y146_BQ),
.Q(CLBLM_L_X12Y156_SLICE_X16Y156_BQ),
.R(CLBLM_R_X13Y155_SLICE_X18Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0054005555015500)
  ) CLBLM_L_X12Y156_SLICE_X16Y156_DLUT (
.I0(CLBLM_R_X11Y159_SLICE_X15Y159_CO5),
.I1(CLBLM_R_X13Y156_SLICE_X18Y156_CO6),
.I2(CLBLM_L_X12Y158_SLICE_X16Y158_BO5),
.I3(CLBLM_R_X11Y158_SLICE_X15Y158_DO6),
.I4(CLBLM_R_X11Y156_SLICE_X14Y156_AQ),
.I5(CLBLM_R_X11Y157_SLICE_X15Y157_BQ),
.O5(CLBLM_L_X12Y156_SLICE_X16Y156_DO5),
.O6(CLBLM_L_X12Y156_SLICE_X16Y156_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333303300312)
  ) CLBLM_L_X12Y156_SLICE_X16Y156_CLUT (
.I0(CLBLM_L_X10Y158_SLICE_X13Y158_AQ),
.I1(CLBLM_R_X11Y159_SLICE_X15Y159_CO5),
.I2(CLBLM_L_X8Y154_SLICE_X10Y154_AQ),
.I3(CLBLM_R_X11Y158_SLICE_X15Y158_DO6),
.I4(CLBLM_L_X12Y158_SLICE_X16Y158_BO5),
.I5(CLBLM_R_X11Y158_SLICE_X14Y158_DO5),
.O5(CLBLM_L_X12Y156_SLICE_X16Y156_CO5),
.O6(CLBLM_L_X12Y156_SLICE_X16Y156_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffeffff)
  ) CLBLM_L_X12Y156_SLICE_X16Y156_BLUT (
.I0(CLBLM_R_X11Y151_SLICE_X15Y151_CO6),
.I1(CLBLL_L_X4Y156_SLICE_X4Y156_BO6),
.I2(CLBLM_L_X12Y156_SLICE_X17Y156_DO6),
.I3(CLBLM_L_X12Y157_SLICE_X16Y157_DO5),
.I4(CLBLM_R_X13Y150_SLICE_X18Y150_AQ),
.I5(CLBLM_R_X11Y157_SLICE_X15Y157_CO6),
.O5(CLBLM_L_X12Y156_SLICE_X16Y156_BO5),
.O6(CLBLM_L_X12Y156_SLICE_X16Y156_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffff7f3f4f0)
  ) CLBLM_L_X12Y156_SLICE_X16Y156_ALUT (
.I0(CLBLM_R_X11Y158_SLICE_X15Y158_BO6),
.I1(CLBLM_R_X11Y159_SLICE_X15Y159_DO5),
.I2(CLBLM_L_X12Y156_SLICE_X16Y156_BO6),
.I3(CLBLM_R_X11Y158_SLICE_X15Y158_AQ),
.I4(CLBLM_L_X10Y158_SLICE_X13Y158_AQ),
.I5(CLBLM_L_X10Y157_SLICE_X12Y157_DO6),
.O5(CLBLM_L_X12Y156_SLICE_X16Y156_AO5),
.O6(CLBLM_L_X12Y156_SLICE_X16Y156_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y156_SLICE_X17Y156_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y156_SLICE_X17Y156_AO6),
.Q(CLBLM_L_X12Y156_SLICE_X17Y156_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y156_SLICE_X17Y156_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y156_SLICE_X17Y156_BO6),
.Q(CLBLM_L_X12Y156_SLICE_X17Y156_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffeffffffff)
  ) CLBLM_L_X12Y156_SLICE_X17Y156_DLUT (
.I0(CLBLM_R_X11Y152_SLICE_X15Y152_BQ),
.I1(CLBLM_L_X10Y153_SLICE_X12Y153_AQ),
.I2(CLBLM_L_X12Y157_SLICE_X16Y157_CQ),
.I3(CLBLM_L_X12Y159_SLICE_X17Y159_CO6),
.I4(CLBLM_R_X13Y151_SLICE_X19Y151_AO6),
.I5(CLBLM_R_X13Y149_SLICE_X18Y149_A5Q),
.O5(CLBLM_L_X12Y156_SLICE_X17Y156_DO5),
.O6(CLBLM_L_X12Y156_SLICE_X17Y156_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00fffb04f708)
  ) CLBLM_L_X12Y156_SLICE_X17Y156_CLUT (
.I0(CLBLM_L_X8Y154_SLICE_X10Y154_AQ),
.I1(CLBLM_R_X11Y158_SLICE_X15Y158_AQ),
.I2(CLBLM_L_X12Y158_SLICE_X16Y158_BO5),
.I3(CLBLM_L_X12Y156_SLICE_X17Y156_AQ),
.I4(CLBLM_L_X12Y158_SLICE_X16Y158_CO5),
.I5(CLBLM_R_X11Y158_SLICE_X15Y158_DO6),
.O5(CLBLM_L_X12Y156_SLICE_X17Y156_CO5),
.O6(CLBLM_L_X12Y156_SLICE_X17Y156_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0afa0acacafa0)
  ) CLBLM_L_X12Y156_SLICE_X17Y156_BLUT (
.I0(CLBLM_R_X11Y149_SLICE_X14Y149_DQ),
.I1(CLBLM_L_X12Y156_SLICE_X17Y156_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y158_SLICE_X15Y158_AQ),
.I4(CLBLM_R_X11Y159_SLICE_X15Y159_DO5),
.I5(CLBLM_R_X11Y158_SLICE_X15Y158_BO6),
.O5(CLBLM_L_X12Y156_SLICE_X17Y156_BO5),
.O6(CLBLM_L_X12Y156_SLICE_X17Y156_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000ff0ff000fc0c)
  ) CLBLM_L_X12Y156_SLICE_X17Y156_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y158_SLICE_X14Y158_DO5),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X13Y150_SLICE_X18Y150_AQ),
.I4(CLBLM_R_X11Y159_SLICE_X15Y159_CO5),
.I5(CLBLM_L_X12Y156_SLICE_X17Y156_CO6),
.O5(CLBLM_L_X12Y156_SLICE_X17Y156_AO5),
.O6(CLBLM_L_X12Y156_SLICE_X17Y156_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y157_SLICE_X16Y157_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y153_SLICE_X16Y153_BO6),
.Q(CLBLM_L_X12Y157_SLICE_X16Y157_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y157_SLICE_X16Y157_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y157_SLICE_X16Y157_AO6),
.Q(CLBLM_L_X12Y157_SLICE_X16Y157_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y157_SLICE_X16Y157_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y157_SLICE_X16Y157_BO6),
.Q(CLBLM_L_X12Y157_SLICE_X16Y157_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y157_SLICE_X16Y157_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y157_SLICE_X16Y157_CO6),
.Q(CLBLM_L_X12Y157_SLICE_X16Y157_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00f000f000aaccaa)
  ) CLBLM_L_X12Y157_SLICE_X16Y157_DLUT (
.I0(CLBLM_R_X11Y156_SLICE_X14Y156_AQ),
.I1(CLBLM_R_X11Y158_SLICE_X14Y158_BQ),
.I2(CLBLM_R_X11Y157_SLICE_X14Y157_CQ),
.I3(CLBLM_R_X11Y159_SLICE_X15Y159_DO5),
.I4(CLBLM_R_X11Y158_SLICE_X15Y158_BO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y157_SLICE_X16Y157_DO5),
.O6(CLBLM_L_X12Y157_SLICE_X16Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaafff0fff0)
  ) CLBLM_L_X12Y157_SLICE_X16Y157_CLUT (
.I0(CLBLM_R_X11Y151_SLICE_X15Y151_BQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y159_SLICE_X12Y159_CO6),
.I3(CLBLM_R_X11Y157_SLICE_X15Y157_DO6),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y157_SLICE_X16Y157_CO5),
.O6(CLBLM_L_X12Y157_SLICE_X16Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0f5e4f5a0a0e4a0)
  ) CLBLM_L_X12Y157_SLICE_X16Y157_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y157_SLICE_X16Y157_BQ),
.I2(CLBLM_R_X11Y155_SLICE_X14Y155_DQ),
.I3(CLBLM_R_X11Y159_SLICE_X15Y159_DO5),
.I4(CLBLM_R_X11Y158_SLICE_X15Y158_BO6),
.I5(CLBLM_L_X12Y157_SLICE_X17Y157_CQ),
.O5(CLBLM_L_X12Y157_SLICE_X16Y157_BO5),
.O6(CLBLM_L_X12Y157_SLICE_X16Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff5200ff0052)
  ) CLBLM_L_X12Y157_SLICE_X16Y157_ALUT (
.I0(CLBLM_L_X12Y155_SLICE_X16Y155_BO5),
.I1(CLBLM_L_X12Y158_SLICE_X16Y158_BO6),
.I2(CLBLM_L_X12Y157_SLICE_X16Y157_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y158_SLICE_X15Y158_BO6),
.I5(CLBLL_L_X4Y148_SLICE_X4Y148_AQ),
.O5(CLBLM_L_X12Y157_SLICE_X16Y157_AO5),
.O6(CLBLM_L_X12Y157_SLICE_X16Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y157_SLICE_X17Y157_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y157_SLICE_X18Y157_AO6),
.Q(CLBLM_L_X12Y157_SLICE_X17Y157_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y157_SLICE_X17Y157_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y157_SLICE_X17Y157_AO6),
.Q(CLBLM_L_X12Y157_SLICE_X17Y157_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y157_SLICE_X17Y157_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y157_SLICE_X17Y157_BO6),
.Q(CLBLM_L_X12Y157_SLICE_X17Y157_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y157_SLICE_X17Y157_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y157_SLICE_X17Y157_CO6),
.Q(CLBLM_L_X12Y157_SLICE_X17Y157_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f03030f0f0f0f)
  ) CLBLM_L_X12Y157_SLICE_X17Y157_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y157_SLICE_X17Y157_CQ),
.I2(CLBLM_R_X11Y158_SLICE_X15Y158_DO6),
.I3(1'b1),
.I4(CLBLM_L_X12Y158_SLICE_X16Y158_BO5),
.I5(CLBLM_L_X12Y159_SLICE_X17Y159_BO6),
.O5(CLBLM_L_X12Y157_SLICE_X17Y157_DO5),
.O6(CLBLM_L_X12Y157_SLICE_X17Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0cff0c00)
  ) CLBLM_L_X12Y157_SLICE_X17Y157_CLUT (
.I0(CLBLM_R_X7Y157_SLICE_X9Y157_CQ),
.I1(CLBLM_L_X12Y157_SLICE_X17Y157_CQ),
.I2(CLBLM_R_X11Y158_SLICE_X15Y158_BO6),
.I3(CLBLM_R_X11Y159_SLICE_X15Y159_DO5),
.I4(CLBLM_L_X12Y156_SLICE_X17Y156_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_L_X12Y157_SLICE_X17Y157_CO5),
.O6(CLBLM_L_X12Y157_SLICE_X17Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0fff09000f0009)
  ) CLBLM_L_X12Y157_SLICE_X17Y157_BLUT (
.I0(CLBLM_R_X13Y157_SLICE_X18Y157_BO6),
.I1(CLBLM_L_X12Y157_SLICE_X17Y157_BQ),
.I2(CLBLM_R_X11Y159_SLICE_X15Y159_CO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y158_SLICE_X14Y158_DO5),
.I5(CLBLM_L_X12Y157_SLICE_X16Y157_CQ),
.O5(CLBLM_L_X12Y157_SLICE_X17Y157_BO5),
.O6(CLBLM_L_X12Y157_SLICE_X17Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f3f3f3f3f3d1)
  ) CLBLM_L_X12Y157_SLICE_X17Y157_ALUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X12Y157_SLICE_X16Y157_A5Q),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLL_L_X4Y158_SLICE_X4Y158_AO6),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLM_L_X12Y157_SLICE_X17Y157_AO5),
.O6(CLBLM_L_X12Y157_SLICE_X17Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y158_SLICE_X16Y158_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y159_SLICE_X16Y159_AO6),
.Q(CLBLM_L_X12Y158_SLICE_X16Y158_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y158_SLICE_X16Y158_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y158_SLICE_X16Y158_AO6),
.Q(CLBLM_L_X12Y158_SLICE_X16Y158_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h92009200ff009200)
  ) CLBLM_L_X12Y158_SLICE_X16Y158_DLUT (
.I0(CLBLM_L_X12Y158_SLICE_X17Y158_AQ),
.I1(CLBLM_L_X12Y158_SLICE_X16Y158_AQ),
.I2(CLBLM_R_X11Y159_SLICE_X15Y159_AQ),
.I3(CLBLM_L_X12Y159_SLICE_X17Y159_AO6),
.I4(CLBLM_L_X12Y159_SLICE_X16Y159_BO5),
.I5(CLBLM_R_X11Y159_SLICE_X14Y159_AQ),
.O5(CLBLM_L_X12Y158_SLICE_X16Y158_DO5),
.O6(CLBLM_L_X12Y158_SLICE_X16Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h838bc3cff0c0f0c0)
  ) CLBLM_L_X12Y158_SLICE_X16Y158_CLUT (
.I0(CLBLM_R_X11Y157_SLICE_X15Y157_AQ),
.I1(CLBLM_L_X12Y158_SLICE_X16Y158_AQ),
.I2(CLBLM_R_X11Y159_SLICE_X15Y159_AQ),
.I3(CLBLM_L_X12Y158_SLICE_X17Y158_AQ),
.I4(CLBLM_R_X11Y159_SLICE_X14Y159_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y158_SLICE_X16Y158_CO5),
.O6(CLBLM_L_X12Y158_SLICE_X16Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000333305ff07ff)
  ) CLBLM_L_X12Y158_SLICE_X16Y158_BLUT (
.I0(CLBLM_L_X12Y157_SLICE_X16Y157_AQ),
.I1(CLBLM_R_X11Y159_SLICE_X15Y159_AQ),
.I2(CLBLM_L_X12Y159_SLICE_X16Y159_BO5),
.I3(CLBLM_L_X12Y155_SLICE_X16Y155_BO5),
.I4(CLBLM_L_X12Y158_SLICE_X17Y158_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y158_SLICE_X16Y158_BO5),
.O6(CLBLM_L_X12Y158_SLICE_X16Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbaba1010abba0110)
  ) CLBLM_L_X12Y158_SLICE_X16Y158_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_L_X12Y158_SLICE_X16Y158_AQ),
.I3(CLBLM_L_X12Y159_SLICE_X17Y159_AO6),
.I4(CLBLM_L_X12Y157_SLICE_X17Y157_AQ),
.I5(CLBLM_L_X12Y158_SLICE_X16Y158_CO6),
.O5(CLBLM_L_X12Y158_SLICE_X16Y158_AO5),
.O6(CLBLM_L_X12Y158_SLICE_X16Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y158_SLICE_X17Y158_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y158_SLICE_X17Y158_AO6),
.Q(CLBLM_L_X12Y158_SLICE_X17Y158_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y158_SLICE_X17Y158_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_L_X12Y158_SLICE_X17Y158_BO6),
.Q(CLBLM_L_X12Y158_SLICE_X17Y158_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaff0000aaff7777)
  ) CLBLM_L_X12Y158_SLICE_X17Y158_DLUT (
.I0(CLBLM_L_X12Y158_SLICE_X16Y158_AQ),
.I1(CLBLM_L_X12Y158_SLICE_X17Y158_AQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y159_SLICE_X15Y159_AQ),
.I4(CLBLM_L_X12Y157_SLICE_X16Y157_AQ),
.I5(CLBLM_R_X11Y159_SLICE_X14Y159_BQ),
.O5(CLBLM_L_X12Y158_SLICE_X17Y158_DO5),
.O6(CLBLM_L_X12Y158_SLICE_X17Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf733fb33ff33f333)
  ) CLBLM_L_X12Y158_SLICE_X17Y158_CLUT (
.I0(CLBLM_L_X12Y152_SLICE_X17Y152_A5Q),
.I1(CLBLM_L_X12Y159_SLICE_X17Y159_CO6),
.I2(CLBLM_R_X11Y158_SLICE_X15Y158_CO6),
.I3(CLBLM_L_X12Y158_SLICE_X17Y158_BQ),
.I4(CLBLM_L_X12Y158_SLICE_X17Y158_DO6),
.I5(CLBLM_R_X11Y159_SLICE_X14Y159_AQ),
.O5(CLBLM_L_X12Y158_SLICE_X17Y158_CO5),
.O6(CLBLM_L_X12Y158_SLICE_X17Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcf3303fccc3000)
  ) CLBLM_L_X12Y158_SLICE_X17Y158_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y158_SLICE_X15Y158_BO6),
.I3(CLBLM_R_X5Y148_SLICE_X6Y148_CO6),
.I4(CLBLM_R_X13Y158_SLICE_X18Y158_AQ),
.I5(CLBLM_L_X12Y158_SLICE_X17Y158_CO6),
.O5(CLBLM_L_X12Y158_SLICE_X17Y158_BO5),
.O6(CLBLM_L_X12Y158_SLICE_X17Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbfe1154aaaa0000)
  ) CLBLM_L_X12Y158_SLICE_X17Y158_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y158_SLICE_X16Y158_DO6),
.I2(CLBLM_R_X11Y158_SLICE_X15Y158_BO6),
.I3(CLBLM_L_X12Y158_SLICE_X17Y158_AQ),
.I4(CLBLM_R_X13Y155_SLICE_X18Y155_AQ),
.I5(RIOB33_X105Y121_IOB_X1Y121_I),
.O5(CLBLM_L_X12Y158_SLICE_X17Y158_AO5),
.O6(CLBLM_L_X12Y158_SLICE_X17Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y159_SLICE_X16Y159_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X12Y158_SLICE_X17Y158_AQ),
.Q(CLBLM_L_X12Y159_SLICE_X16Y159_AQ),
.R(CLBLM_R_X13Y155_SLICE_X18Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_L_X12Y159_SLICE_X16Y159_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_L_X10Y150_SLICE_X12Y150_CQ),
.Q(CLBLM_L_X12Y159_SLICE_X16Y159_BQ),
.R(CLBLM_R_X13Y155_SLICE_X18Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y159_SLICE_X16Y159_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y159_SLICE_X16Y159_DO5),
.O6(CLBLM_L_X12Y159_SLICE_X16Y159_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5555f0ff000f)
  ) CLBLM_L_X12Y159_SLICE_X16Y159_CLUT (
.I0(RIOB33_X105Y143_IOB_X1Y143_I),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y152_SLICE_X3Y152_AO5),
.I4(CLBLM_L_X12Y159_SLICE_X16Y159_BQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y159_SLICE_X16Y159_CO5),
.O6(CLBLM_L_X12Y159_SLICE_X16Y159_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000008000008888)
  ) CLBLM_L_X12Y159_SLICE_X16Y159_BLUT (
.I0(CLBLM_L_X12Y158_SLICE_X16Y158_AQ),
.I1(CLBLM_R_X11Y159_SLICE_X14Y159_BQ),
.I2(CLBLM_L_X12Y159_SLICE_X17Y159_AO6),
.I3(CLBLM_R_X11Y159_SLICE_X14Y159_AQ),
.I4(CLBLM_R_X11Y157_SLICE_X15Y157_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y159_SLICE_X16Y159_BO5),
.O6(CLBLM_L_X12Y159_SLICE_X16Y159_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f0aaf3f3f3f3)
  ) CLBLM_L_X12Y159_SLICE_X16Y159_ALUT (
.I0(CLBLM_L_X8Y153_SLICE_X11Y153_CQ),
.I1(RIOB33_X105Y143_IOB_X1Y143_I),
.I2(CLBLM_L_X12Y159_SLICE_X16Y159_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_L_X12Y159_SLICE_X16Y159_AO5),
.O6(CLBLM_L_X12Y159_SLICE_X16Y159_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y159_SLICE_X17Y159_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y159_SLICE_X17Y159_DO5),
.O6(CLBLM_L_X12Y159_SLICE_X17Y159_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffcfffffffcf)
  ) CLBLM_L_X12Y159_SLICE_X17Y159_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y159_SLICE_X14Y159_AQ),
.I2(CLBLM_L_X12Y158_SLICE_X17Y158_AQ),
.I3(CLBLM_R_X11Y159_SLICE_X15Y159_AQ),
.I4(CLBLM_L_X12Y158_SLICE_X16Y158_AQ),
.I5(1'b1),
.O5(CLBLM_L_X12Y159_SLICE_X17Y159_CO5),
.O6(CLBLM_L_X12Y159_SLICE_X17Y159_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00400302c0c00000)
  ) CLBLM_L_X12Y159_SLICE_X17Y159_BLUT (
.I0(CLBLM_L_X12Y158_SLICE_X16Y158_AQ),
.I1(CLBLM_L_X12Y157_SLICE_X17Y157_BQ),
.I2(CLBLM_L_X12Y156_SLICE_X17Y156_AQ),
.I3(CLBLM_L_X12Y158_SLICE_X17Y158_AQ),
.I4(CLBLM_L_X8Y154_SLICE_X10Y154_AQ),
.I5(CLBLM_R_X11Y159_SLICE_X15Y159_AQ),
.O5(CLBLM_L_X12Y159_SLICE_X17Y159_BO5),
.O6(CLBLM_L_X12Y159_SLICE_X17Y159_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3330030033300300)
  ) CLBLM_L_X12Y159_SLICE_X17Y159_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y158_SLICE_X16Y158_BO5),
.I2(CLBLM_R_X13Y158_SLICE_X18Y158_AQ),
.I3(CLBLM_R_X13Y159_SLICE_X18Y159_AO6),
.I4(CLBLM_R_X13Y159_SLICE_X18Y159_BO6),
.I5(1'b1),
.O5(CLBLM_L_X12Y159_SLICE_X17Y159_AO5),
.O6(CLBLM_L_X12Y159_SLICE_X17Y159_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y156_SLICE_X22Y156_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y156_SLICE_X22Y156_DO5),
.O6(CLBLM_L_X16Y156_SLICE_X22Y156_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y156_SLICE_X22Y156_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y156_SLICE_X22Y156_CO5),
.O6(CLBLM_L_X16Y156_SLICE_X22Y156_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y156_SLICE_X22Y156_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y156_SLICE_X22Y156_BO5),
.O6(CLBLM_L_X16Y156_SLICE_X22Y156_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff5fff5fffffff0)
  ) CLBLM_L_X16Y156_SLICE_X22Y156_ALUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(1'b1),
.I2(RIOB33_X105Y129_IOB_X1Y129_I),
.I3(RIOB33_X105Y129_IOB_X1Y130_I),
.I4(RIOB33_X105Y127_IOB_X1Y128_I),
.I5(1'b1),
.O5(CLBLM_L_X16Y156_SLICE_X22Y156_AO5),
.O6(CLBLM_L_X16Y156_SLICE_X22Y156_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y156_SLICE_X23Y156_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y156_SLICE_X23Y156_DO5),
.O6(CLBLM_L_X16Y156_SLICE_X23Y156_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y156_SLICE_X23Y156_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y156_SLICE_X23Y156_CO5),
.O6(CLBLM_L_X16Y156_SLICE_X23Y156_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y156_SLICE_X23Y156_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y156_SLICE_X23Y156_BO5),
.O6(CLBLM_L_X16Y156_SLICE_X23Y156_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X16Y156_SLICE_X23Y156_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X16Y156_SLICE_X23Y156_AO5),
.O6(CLBLM_L_X16Y156_SLICE_X23Y156_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X2Y142_DO5),
.O6(CLBLM_R_X3Y142_SLICE_X2Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X2Y142_CO5),
.O6(CLBLM_R_X3Y142_SLICE_X2Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X2Y142_BO5),
.O6(CLBLM_R_X3Y142_SLICE_X2Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y142_SLICE_X2Y142_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y142_SLICE_X2Y142_AO5),
.O6(CLBLM_R_X3Y142_SLICE_X2Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa55555555)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_DLUT (
.I0(CLBLM_R_X3Y152_SLICE_X3Y152_AO5),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X4Y148_SLICE_X4Y148_CO6),
.O5(CLBLM_R_X3Y142_SLICE_X3Y142_DO5),
.O6(CLBLM_R_X3Y142_SLICE_X3Y142_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f5f0f5f0f5f)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_CLUT (
.I0(CLBLM_R_X3Y142_SLICE_X3Y142_AO6),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLL_L_X4Y147_SLICE_X4Y147_AO6),
.I4(LIOB33_X0Y53_IOB_X0Y53_I),
.I5(CLBLL_L_X4Y154_SLICE_X4Y154_BO6),
.O5(CLBLM_R_X3Y142_SLICE_X3Y142_CO5),
.O6(CLBLM_R_X3Y142_SLICE_X3Y142_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000040ccccccccc)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_BLUT (
.I0(LIOB33_X0Y53_IOB_X0Y53_I),
.I1(CLBLL_L_X4Y148_SLICE_X4Y148_CO6),
.I2(CLBLL_L_X4Y147_SLICE_X4Y147_AO6),
.I3(CLBLL_L_X4Y154_SLICE_X4Y154_BO6),
.I4(CLBLM_R_X3Y142_SLICE_X3Y142_AO6),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X3Y142_SLICE_X3Y142_BO5),
.O6(CLBLM_R_X3Y142_SLICE_X3Y142_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaeaa00000c00)
  ) CLBLM_R_X3Y142_SLICE_X3Y142_ALUT (
.I0(LIOB33_X0Y51_IOB_X0Y51_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLL_L_X4Y151_SLICE_X4Y151_CQ),
.I3(CLBLL_L_X4Y152_SLICE_X4Y152_AQ),
.I4(CLBLL_L_X4Y153_SLICE_X4Y153_AO6),
.I5(CLBLM_R_X3Y156_SLICE_X2Y156_DO6),
.O5(CLBLM_R_X3Y142_SLICE_X3Y142_AO5),
.O6(CLBLM_R_X3Y142_SLICE_X3Y142_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y150_SLICE_X2Y150_BO6),
.Q(CLBLM_R_X3Y150_SLICE_X2Y150_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y150_SLICE_X2Y150_AO6),
.Q(CLBLM_R_X3Y150_SLICE_X2Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fffffff5fffffff)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_DLUT (
.I0(CLBLM_L_X8Y147_SLICE_X11Y147_CO6),
.I1(1'b1),
.I2(CLBLM_R_X3Y150_SLICE_X2Y150_AQ),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_CQ),
.I4(CLBLM_R_X3Y150_SLICE_X2Y150_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y150_SLICE_X2Y150_DO5),
.O6(CLBLM_R_X3Y150_SLICE_X2Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0301000002000000)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLM_R_X3Y152_SLICE_X2Y152_AO5),
.I2(CLBLL_L_X4Y157_SLICE_X4Y157_CO6),
.I3(LIOB33_X0Y57_IOB_X0Y58_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_R_X3Y151_SLICE_X2Y151_BQ),
.O5(CLBLM_R_X3Y150_SLICE_X2Y150_CO5),
.O6(CLBLM_R_X3Y150_SLICE_X2Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf202f8083333ffff)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_BLUT (
.I0(CLBLL_L_X4Y149_SLICE_X4Y149_DO6),
.I1(CLBLM_R_X3Y150_SLICE_X2Y150_A5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X3Y151_SLICE_X2Y151_BQ),
.I4(CLBLM_L_X8Y147_SLICE_X11Y147_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y150_SLICE_X2Y150_BO5),
.O6(CLBLM_R_X3Y150_SLICE_X2Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hedcc2100fccc3000)
  ) CLBLM_R_X3Y150_SLICE_X2Y150_ALUT (
.I0(CLBLM_R_X3Y150_SLICE_X2Y150_BO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X3Y150_SLICE_X2Y150_AQ),
.I3(CLBLL_L_X4Y149_SLICE_X4Y149_DO6),
.I4(CLBLM_L_X12Y153_SLICE_X17Y153_CQ),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_CQ),
.O5(CLBLM_R_X3Y150_SLICE_X2Y150_AO5),
.O6(CLBLM_R_X3Y150_SLICE_X2Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y150_SLICE_X3Y150_AO6),
.Q(CLBLM_R_X3Y150_SLICE_X3Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y150_SLICE_X3Y150_BO6),
.Q(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y150_SLICE_X3Y150_CO6),
.Q(CLBLM_R_X3Y150_SLICE_X3Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y150_SLICE_X3Y150_DO5),
.O6(CLBLM_R_X3Y150_SLICE_X3Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffc3000000c300)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_CQ),
.I2(CLBLM_R_X3Y150_SLICE_X2Y150_BO5),
.I3(CLBLL_L_X4Y149_SLICE_X4Y149_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y149_SLICE_X4Y149_AQ),
.O5(CLBLM_R_X3Y150_SLICE_X3Y150_CO5),
.O6(CLBLM_R_X3Y150_SLICE_X3Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff880088ff220022)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_BLUT (
.I0(CLBLL_L_X4Y149_SLICE_X5Y149_CO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y148_SLICE_X12Y148_AQ),
.I5(CLBLM_R_X3Y151_SLICE_X3Y151_AO5),
.O5(CLBLM_R_X3Y150_SLICE_X3Y150_BO5),
.O6(CLBLM_R_X3Y150_SLICE_X3Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00a0a0ff002828)
  ) CLBLM_R_X3Y150_SLICE_X3Y150_ALUT (
.I0(CLBLL_L_X4Y149_SLICE_X5Y149_CO6),
.I1(CLBLM_R_X3Y150_SLICE_X3Y150_BQ),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_AQ),
.I3(CLBLM_R_X11Y154_SLICE_X15Y154_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X3Y151_SLICE_X3Y151_AO5),
.O5(CLBLM_R_X3Y150_SLICE_X3Y150_AO5),
.O6(CLBLM_R_X3Y150_SLICE_X3Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y151_SLICE_X2Y151_AO6),
.Q(CLBLM_R_X3Y151_SLICE_X2Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y151_SLICE_X2Y151_BO6),
.Q(CLBLM_R_X3Y151_SLICE_X2Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h30ba30baffff30ba)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_DLUT (
.I0(CLBLM_R_X3Y150_SLICE_X2Y150_AQ),
.I1(CLBLL_L_X2Y154_SLICE_X1Y154_AO5),
.I2(LIOB33_X0Y57_IOB_X0Y57_I),
.I3(CLBLM_R_X3Y151_SLICE_X2Y151_CO6),
.I4(LIOB33_X0Y61_IOB_X0Y62_I),
.I5(CLBLL_L_X2Y153_SLICE_X1Y153_AO5),
.O5(CLBLM_R_X3Y151_SLICE_X2Y151_DO5),
.O6(CLBLM_R_X3Y151_SLICE_X2Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffbffffffffb)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_CLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(CLBLL_L_X4Y157_SLICE_X4Y157_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y151_SLICE_X2Y151_CO5),
.O6(CLBLM_R_X3Y151_SLICE_X2Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaac000aaaac0f0)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_BLUT (
.I0(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.I1(CLBLM_R_X3Y151_SLICE_X2Y151_BQ),
.I2(CLBLL_L_X4Y149_SLICE_X4Y149_DO6),
.I3(CLBLM_R_X3Y150_SLICE_X2Y150_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X3Y151_SLICE_X2Y151_AO5),
.O5(CLBLM_R_X3Y151_SLICE_X2Y151_BO5),
.O6(CLBLM_R_X3Y151_SLICE_X2Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heaaa0000c0000000)
  ) CLBLM_R_X3Y151_SLICE_X2Y151_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y151_SLICE_X2Y151_BQ),
.I2(CLBLM_R_X3Y150_SLICE_X3Y150_CQ),
.I3(CLBLM_R_X3Y150_SLICE_X2Y150_A5Q),
.I4(CLBLM_R_X3Y150_SLICE_X2Y150_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y151_SLICE_X2Y151_AO5),
.O6(CLBLM_R_X3Y151_SLICE_X2Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X3Y151_SLICE_X3Y151_AO6),
.Q(CLBLM_R_X3Y151_SLICE_X3Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y151_SLICE_X3Y151_DO5),
.O6(CLBLM_R_X3Y151_SLICE_X3Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff0fffffffc)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y150_SLICE_X7Y150_CQ),
.I2(CLBLM_R_X3Y152_SLICE_X2Y152_CO6),
.I3(CLBLM_R_X3Y150_SLICE_X2Y150_CO6),
.I4(CLBLM_R_X3Y152_SLICE_X3Y152_DO6),
.I5(CLBLM_R_X3Y151_SLICE_X2Y151_CO5),
.O5(CLBLM_R_X3Y151_SLICE_X3Y151_CO5),
.O6(CLBLM_R_X3Y151_SLICE_X3Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbfffbfff0ff0000)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_BLUT (
.I0(RIOB33_X105Y127_IOB_X1Y128_I),
.I1(CLBLM_R_X3Y152_SLICE_X3Y152_AO5),
.I2(RIOB33_X105Y129_IOB_X1Y129_I),
.I3(RIOB33_X105Y137_IOB_X1Y137_I),
.I4(CLBLL_L_X4Y151_SLICE_X4Y151_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y151_SLICE_X3Y151_BO5),
.O6(CLBLM_R_X3Y151_SLICE_X3Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00ebc3cfcfcfcf)
  ) CLBLM_R_X3Y151_SLICE_X3Y151_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y155_SLICE_X16Y155_CO6),
.I2(CLBLM_R_X3Y151_SLICE_X3Y151_AQ),
.I3(CLBLM_R_X5Y151_SLICE_X6Y151_C5Q),
.I4(CLBLL_L_X4Y150_SLICE_X4Y150_DO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y151_SLICE_X3Y151_AO5),
.O6(CLBLM_R_X3Y151_SLICE_X3Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9999666666669999)
  ) CLBLM_R_X3Y152_SLICE_X2Y152_DLUT (
.I0(CLBLL_L_X4Y153_SLICE_X4Y153_AO6),
.I1(CLBLL_L_X4Y154_SLICE_X4Y154_BO6),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y156_SLICE_X2Y156_DO6),
.I5(CLBLM_R_X3Y155_SLICE_X2Y155_BO6),
.O5(CLBLM_R_X3Y152_SLICE_X2Y152_DO5),
.O6(CLBLM_R_X3Y152_SLICE_X2Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h222f2222000f0000)
  ) CLBLM_R_X3Y152_SLICE_X2Y152_CLUT (
.I0(RIOB33_X105Y117_IOB_X1Y117_I),
.I1(CLBLM_R_X3Y158_SLICE_X2Y158_AO5),
.I2(CLBLL_L_X4Y157_SLICE_X4Y157_CO6),
.I3(CLBLL_L_X2Y155_SLICE_X1Y155_CO6),
.I4(LIOB33_X0Y63_IOB_X0Y63_I),
.I5(CLBLM_R_X3Y156_SLICE_X3Y156_AO6),
.O5(CLBLM_R_X3Y152_SLICE_X2Y152_CO5),
.O6(CLBLM_R_X3Y152_SLICE_X2Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfdf0055cfcf0000)
  ) CLBLM_R_X3Y152_SLICE_X2Y152_BLUT (
.I0(CLBLL_L_X4Y157_SLICE_X4Y157_CO6),
.I1(RIOB33_X105Y129_IOB_X1Y129_I),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(CLBLL_L_X2Y155_SLICE_X1Y155_CO6),
.I4(CLBLL_L_X4Y151_SLICE_X4Y151_D5Q),
.I5(LIOB33_X0Y67_IOB_X0Y68_I),
.O5(CLBLM_R_X3Y152_SLICE_X2Y152_BO5),
.O6(CLBLM_R_X3Y152_SLICE_X2Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h77ff77ffccffccff)
  ) CLBLM_R_X3Y152_SLICE_X2Y152_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(1'b1),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y152_SLICE_X2Y152_AO5),
.O6(CLBLM_R_X3Y152_SLICE_X2Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000abaa0300)
  ) CLBLM_R_X3Y152_SLICE_X3Y152_DLUT (
.I0(CLBLM_R_X3Y152_SLICE_X3Y152_AO6),
.I1(CLBLM_R_X3Y152_SLICE_X2Y152_AO6),
.I2(CLBLL_L_X4Y157_SLICE_X4Y157_CO6),
.I3(CLBLL_L_X4Y149_SLICE_X4Y149_AQ),
.I4(CLBLL_L_X4Y151_SLICE_X4Y151_DQ),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X3Y152_SLICE_X3Y152_DO5),
.O6(CLBLM_R_X3Y152_SLICE_X3Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f2f00000022)
  ) CLBLM_R_X3Y152_SLICE_X3Y152_CLUT (
.I0(CLBLL_L_X4Y155_SLICE_X4Y155_BQ),
.I1(CLBLM_R_X3Y152_SLICE_X2Y152_AO6),
.I2(CLBLL_L_X2Y155_SLICE_X1Y155_CO5),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(CLBLL_L_X4Y157_SLICE_X4Y157_CO6),
.I5(CLBLM_R_X3Y150_SLICE_X3Y150_CQ),
.O5(CLBLM_R_X3Y152_SLICE_X3Y152_CO5),
.O6(CLBLM_R_X3Y152_SLICE_X3Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc33c3cc30000aaaa)
  ) CLBLM_R_X3Y152_SLICE_X3Y152_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLL_L_X4Y154_SLICE_X5Y154_BO6),
.I2(CLBLM_R_X5Y155_SLICE_X6Y155_DO6),
.I3(CLBLL_L_X4Y153_SLICE_X4Y153_BO6),
.I4(CLBLL_L_X4Y154_SLICE_X5Y154_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y152_SLICE_X3Y152_BO5),
.O6(CLBLM_R_X3Y152_SLICE_X3Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5555c33cc936)
  ) CLBLM_R_X3Y152_SLICE_X3Y152_ALUT (
.I0(RIOB33_X105Y137_IOB_X1Y137_I),
.I1(CLBLM_R_X3Y152_SLICE_X2Y152_DO6),
.I2(CLBLL_L_X4Y158_SLICE_X5Y158_AQ),
.I3(CLBLM_R_X3Y152_SLICE_X3Y152_BO6),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y152_SLICE_X3Y152_AO5),
.O6(CLBLM_R_X3Y152_SLICE_X3Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haeaeaeaeffaeffae)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_DLUT (
.I0(CLBLM_R_X3Y152_SLICE_X2Y152_BO6),
.I1(CLBLM_L_X8Y154_SLICE_X11Y154_AQ),
.I2(CLBLM_R_X3Y153_SLICE_X3Y153_AO6),
.I3(CLBLL_L_X4Y152_SLICE_X5Y152_CQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y151_SLICE_X2Y151_CO6),
.O5(CLBLM_R_X3Y153_SLICE_X2Y153_DO5),
.O6(CLBLM_R_X3Y153_SLICE_X2Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffdfff)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_CLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(CLBLM_R_X3Y158_SLICE_X2Y158_AO5),
.I5(RIOB33_X105Y133_IOB_X1Y134_I),
.O5(CLBLM_R_X3Y153_SLICE_X2Y153_CO5),
.O6(CLBLM_R_X3Y153_SLICE_X2Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h404040404040ff40)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_BLUT (
.I0(CLBLM_R_X3Y158_SLICE_X2Y158_AO5),
.I1(CLBLM_R_X3Y156_SLICE_X3Y156_AO6),
.I2(RIOB33_X105Y115_IOB_X1Y115_I),
.I3(LIOB33_X0Y55_IOB_X0Y55_I),
.I4(CLBLL_L_X4Y157_SLICE_X4Y157_CO6),
.I5(CLBLM_R_X3Y153_SLICE_X2Y153_AO5),
.O5(CLBLM_R_X3Y153_SLICE_X2Y153_BO5),
.O6(CLBLM_R_X3Y153_SLICE_X2Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbffffffcfffffff)
  ) CLBLM_R_X3Y153_SLICE_X2Y153_ALUT (
.I0(CLBLL_L_X4Y157_SLICE_X4Y157_CO6),
.I1(RIOB33_X105Y133_IOB_X1Y133_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y153_SLICE_X2Y153_AO5),
.O6(CLBLM_R_X3Y153_SLICE_X2Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff50ff50ffffff50)
  ) CLBLM_R_X3Y153_SLICE_X3Y153_DLUT (
.I0(CLBLM_R_X3Y153_SLICE_X3Y153_AO6),
.I1(1'b1),
.I2(CLBLM_R_X11Y152_SLICE_X14Y152_AQ),
.I3(CLBLM_R_X3Y152_SLICE_X3Y152_CO6),
.I4(LIOB33_X0Y61_IOB_X0Y61_I),
.I5(CLBLL_L_X2Y153_SLICE_X1Y153_AO5),
.O5(CLBLM_R_X3Y153_SLICE_X3Y153_DO5),
.O6(CLBLM_R_X3Y153_SLICE_X3Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfffcfefcfcfcfe)
  ) CLBLM_R_X3Y153_SLICE_X3Y153_CLUT (
.I0(CLBLM_R_X5Y154_SLICE_X6Y154_AQ),
.I1(CLBLL_L_X2Y153_SLICE_X0Y153_AO6),
.I2(CLBLM_R_X3Y153_SLICE_X2Y153_BO6),
.I3(CLBLM_R_X3Y153_SLICE_X3Y153_AO5),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLM_R_X5Y153_SLICE_X7Y153_AQ),
.O5(CLBLM_R_X3Y153_SLICE_X3Y153_CO5),
.O6(CLBLM_R_X3Y153_SLICE_X3Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0303030300010203)
  ) CLBLM_R_X3Y153_SLICE_X3Y153_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLM_R_X3Y155_SLICE_X3Y155_DO6),
.I2(CLBLL_L_X2Y153_SLICE_X1Y153_BO6),
.I3(CLBLM_R_X5Y154_SLICE_X6Y154_AQ),
.I4(CLBLM_R_X5Y153_SLICE_X7Y153_AQ),
.I5(CLBLM_R_X3Y153_SLICE_X3Y153_AO5),
.O5(CLBLM_R_X3Y153_SLICE_X3Y153_BO5),
.O6(CLBLM_R_X3Y153_SLICE_X3Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffdffffffffffcf)
  ) CLBLM_R_X3Y153_SLICE_X3Y153_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLL_L_X4Y157_SLICE_X4Y157_CO5),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y153_SLICE_X3Y153_AO5),
.O6(CLBLM_R_X3Y153_SLICE_X3Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffa0ffffffec)
  ) CLBLM_R_X3Y154_SLICE_X2Y154_DLUT (
.I0(CLBLM_R_X3Y152_SLICE_X3Y152_AO6),
.I1(LIOB33_X0Y59_IOB_X0Y59_I),
.I2(CLBLL_L_X4Y155_SLICE_X5Y155_AQ),
.I3(CLBLM_R_X3Y154_SLICE_X2Y154_CO6),
.I4(CLBLM_R_X3Y155_SLICE_X2Y155_DO6),
.I5(CLBLL_L_X2Y153_SLICE_X1Y153_AO5),
.O5(CLBLM_R_X3Y154_SLICE_X2Y154_DO5),
.O6(CLBLM_R_X3Y154_SLICE_X2Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h05cd050500cc0000)
  ) CLBLM_R_X3Y154_SLICE_X2Y154_CLUT (
.I0(CLBLL_L_X4Y157_SLICE_X4Y157_CO6),
.I1(CLBLM_R_X3Y156_SLICE_X3Y156_AO6),
.I2(CLBLL_L_X2Y155_SLICE_X1Y155_CO5),
.I3(CLBLM_R_X3Y158_SLICE_X2Y158_AO5),
.I4(RIOB33_X105Y113_IOB_X1Y114_I),
.I5(CLBLM_R_X3Y150_SLICE_X2Y150_A5Q),
.O5(CLBLM_R_X3Y154_SLICE_X2Y154_CO5),
.O6(CLBLM_R_X3Y154_SLICE_X2Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff73ff00ff50)
  ) CLBLM_R_X3Y154_SLICE_X2Y154_BLUT (
.I0(CLBLL_L_X2Y155_SLICE_X1Y155_CO5),
.I1(CLBLL_L_X2Y155_SLICE_X1Y155_CO6),
.I2(CLBLL_L_X4Y152_SLICE_X5Y152_CQ),
.I3(CLBLM_R_X3Y151_SLICE_X3Y151_BO5),
.I4(CLBLL_L_X4Y157_SLICE_X4Y157_CO6),
.I5(LIOB33_X0Y67_IOB_X0Y68_I),
.O5(CLBLM_R_X3Y154_SLICE_X2Y154_BO5),
.O6(CLBLM_R_X3Y154_SLICE_X2Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000010000)
  ) CLBLM_R_X3Y154_SLICE_X2Y154_ALUT (
.I0(CLBLL_L_X4Y154_SLICE_X5Y154_CO6),
.I1(CLBLL_L_X4Y154_SLICE_X4Y154_AO6),
.I2(CLBLL_L_X4Y154_SLICE_X4Y154_BO6),
.I3(CLBLM_R_X3Y156_SLICE_X3Y156_BO6),
.I4(CLBLL_L_X4Y153_SLICE_X4Y153_AO6),
.I5(CLBLL_L_X4Y154_SLICE_X5Y154_BO6),
.O5(CLBLM_R_X3Y154_SLICE_X2Y154_AO5),
.O6(CLBLM_R_X3Y154_SLICE_X2Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffdfdffff)
  ) CLBLM_R_X3Y154_SLICE_X3Y154_DLUT (
.I0(CLBLM_R_X3Y154_SLICE_X3Y154_AO6),
.I1(CLBLL_L_X2Y155_SLICE_X1Y155_BO6),
.I2(CLBLM_R_X3Y157_SLICE_X2Y157_CO6),
.I3(1'b1),
.I4(CLBLL_L_X4Y156_SLICE_X4Y156_BO5),
.I5(CLBLL_L_X2Y154_SLICE_X1Y154_AO6),
.O5(CLBLM_R_X3Y154_SLICE_X3Y154_DO5),
.O6(CLBLM_R_X3Y154_SLICE_X3Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000001000)
  ) CLBLM_R_X3Y154_SLICE_X3Y154_CLUT (
.I0(CLBLM_R_X3Y155_SLICE_X2Y155_CO6),
.I1(CLBLM_R_X3Y155_SLICE_X2Y155_DO6),
.I2(CLBLL_L_X4Y156_SLICE_X4Y156_BO5),
.I3(CLBLM_R_X3Y153_SLICE_X3Y153_AO5),
.I4(CLBLL_L_X2Y155_SLICE_X1Y155_BO6),
.I5(CLBLL_L_X2Y154_SLICE_X1Y154_AO6),
.O5(CLBLM_R_X3Y154_SLICE_X3Y154_CO5),
.O6(CLBLM_R_X3Y154_SLICE_X3Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000020000)
  ) CLBLM_R_X3Y154_SLICE_X3Y154_BLUT (
.I0(CLBLL_L_X4Y156_SLICE_X4Y156_BO5),
.I1(CLBLM_R_X3Y155_SLICE_X2Y155_DO6),
.I2(CLBLM_R_X3Y157_SLICE_X2Y157_CO6),
.I3(CLBLL_L_X2Y154_SLICE_X1Y154_AO6),
.I4(CLBLM_R_X3Y154_SLICE_X3Y154_AO6),
.I5(CLBLL_L_X2Y155_SLICE_X1Y155_BO6),
.O5(CLBLM_R_X3Y154_SLICE_X3Y154_BO5),
.O6(CLBLM_R_X3Y154_SLICE_X3Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffbffffffffd)
  ) CLBLM_R_X3Y154_SLICE_X3Y154_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(CLBLL_L_X4Y157_SLICE_X4Y157_CO5),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y154_SLICE_X3Y154_AO5),
.O6(CLBLM_R_X3Y154_SLICE_X3Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0010000000000000)
  ) CLBLM_R_X3Y155_SLICE_X2Y155_DLUT (
.I0(RIOB33_X105Y129_IOB_X1Y130_I),
.I1(CLBLM_R_X3Y152_SLICE_X3Y152_AO6),
.I2(RIOB33_X105Y135_IOB_X1Y135_I),
.I3(RIOB33_X105Y131_IOB_X1Y131_I),
.I4(CLBLL_L_X4Y157_SLICE_X5Y157_AO6),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLM_R_X3Y155_SLICE_X2Y155_DO5),
.O6(CLBLM_R_X3Y155_SLICE_X2Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccdcccccccddcccd)
  ) CLBLM_R_X3Y155_SLICE_X2Y155_CLUT (
.I0(RIOB33_X105Y129_IOB_X1Y130_I),
.I1(CLBLM_R_X3Y152_SLICE_X3Y152_AO6),
.I2(RIOB33_X105Y135_IOB_X1Y135_I),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(CLBLL_L_X4Y157_SLICE_X5Y157_AO6),
.I5(CLBLL_L_X2Y155_SLICE_X1Y155_CO5),
.O5(CLBLM_R_X3Y155_SLICE_X2Y155_CO5),
.O6(CLBLM_R_X3Y155_SLICE_X2Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffabffabffffffab)
  ) CLBLM_R_X3Y155_SLICE_X2Y155_BLUT (
.I0(CLBLM_R_X3Y153_SLICE_X2Y153_DO6),
.I1(CLBLL_L_X2Y155_SLICE_X1Y155_DO6),
.I2(CLBLM_R_X3Y155_SLICE_X3Y155_CO6),
.I3(CLBLM_R_X3Y157_SLICE_X3Y157_DO6),
.I4(CLBLL_L_X4Y152_SLICE_X5Y152_AQ),
.I5(CLBLM_R_X3Y157_SLICE_X2Y157_AO5),
.O5(CLBLM_R_X3Y155_SLICE_X2Y155_BO5),
.O6(CLBLM_R_X3Y155_SLICE_X2Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0cac0cccccccc)
  ) CLBLM_R_X3Y155_SLICE_X2Y155_ALUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(CLBLL_L_X4Y155_SLICE_X5Y155_AQ),
.I2(RIOB33_X105Y129_IOB_X1Y129_I),
.I3(CLBLM_R_X3Y156_SLICE_X3Y156_AO6),
.I4(RIOB33_X105Y129_IOB_X1Y130_I),
.I5(RIOB33_X105Y137_IOB_X1Y137_I),
.O5(CLBLM_R_X3Y155_SLICE_X2Y155_AO5),
.O6(CLBLM_R_X3Y155_SLICE_X2Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000010)
  ) CLBLM_R_X3Y155_SLICE_X3Y155_DLUT (
.I0(CLBLM_R_X3Y157_SLICE_X2Y157_DO6),
.I1(CLBLM_R_X3Y155_SLICE_X2Y155_CO6),
.I2(CLBLL_L_X4Y156_SLICE_X4Y156_BO5),
.I3(CLBLL_L_X2Y155_SLICE_X1Y155_BO6),
.I4(CLBLM_R_X3Y156_SLICE_X3Y156_DO6),
.I5(CLBLL_L_X2Y154_SLICE_X1Y154_AO6),
.O5(CLBLM_R_X3Y155_SLICE_X3Y155_DO5),
.O6(CLBLM_R_X3Y155_SLICE_X3Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff75ffff)
  ) CLBLM_R_X3Y155_SLICE_X3Y155_CLUT (
.I0(CLBLM_R_X3Y154_SLICE_X3Y154_AO6),
.I1(CLBLL_L_X4Y157_SLICE_X4Y157_CO6),
.I2(CLBLL_L_X4Y157_SLICE_X5Y157_AO6),
.I3(CLBLM_R_X3Y152_SLICE_X3Y152_AO6),
.I4(CLBLL_L_X4Y156_SLICE_X4Y156_BO5),
.I5(CLBLL_L_X2Y154_SLICE_X1Y154_AO6),
.O5(CLBLM_R_X3Y155_SLICE_X3Y155_CO5),
.O6(CLBLM_R_X3Y155_SLICE_X3Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001000000000000)
  ) CLBLM_R_X3Y155_SLICE_X3Y155_BLUT (
.I0(CLBLL_L_X2Y155_SLICE_X1Y155_AO6),
.I1(CLBLL_L_X2Y154_SLICE_X1Y154_AO6),
.I2(CLBLM_R_X3Y155_SLICE_X2Y155_CO6),
.I3(CLBLM_R_X3Y155_SLICE_X2Y155_DO6),
.I4(CLBLL_L_X4Y156_SLICE_X4Y156_CO5),
.I5(CLBLL_L_X4Y156_SLICE_X4Y156_BO5),
.O5(CLBLM_R_X3Y155_SLICE_X3Y155_BO5),
.O6(CLBLM_R_X3Y155_SLICE_X3Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000400000)
  ) CLBLM_R_X3Y155_SLICE_X3Y155_ALUT (
.I0(CLBLM_R_X3Y157_SLICE_X2Y157_CO6),
.I1(CLBLL_L_X4Y156_SLICE_X4Y156_BO5),
.I2(CLBLM_R_X3Y154_SLICE_X3Y154_AO6),
.I3(CLBLL_L_X2Y154_SLICE_X1Y154_AO6),
.I4(CLBLL_L_X4Y156_SLICE_X4Y156_CO5),
.I5(CLBLL_L_X2Y155_SLICE_X1Y155_BO6),
.O5(CLBLM_R_X3Y155_SLICE_X3Y155_AO5),
.O6(CLBLM_R_X3Y155_SLICE_X3Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X3Y156_SLICE_X2Y156_DLUT (
.I0(CLBLL_L_X4Y156_SLICE_X5Y156_AO6),
.I1(CLBLM_R_X3Y154_SLICE_X2Y154_DO6),
.I2(CLBLL_L_X2Y153_SLICE_X1Y153_DO6),
.I3(CLBLM_R_X7Y158_SLICE_X9Y158_DO6),
.I4(CLBLM_R_X3Y155_SLICE_X3Y155_DO6),
.I5(CLBLL_L_X4Y157_SLICE_X5Y157_BO6),
.O5(CLBLM_R_X3Y156_SLICE_X2Y156_DO5),
.O6(CLBLM_R_X3Y156_SLICE_X2Y156_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000002000000)
  ) CLBLM_R_X3Y156_SLICE_X2Y156_CLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLL_L_X4Y157_SLICE_X4Y157_CO6),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(LIOB33_X0Y69_IOB_X0Y70_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X3Y156_SLICE_X2Y156_CO5),
.O6(CLBLM_R_X3Y156_SLICE_X2Y156_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0400000000000000)
  ) CLBLM_R_X3Y156_SLICE_X2Y156_BLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(CLBLL_L_X4Y157_SLICE_X4Y157_CO6),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(LIOB33_X0Y59_IOB_X0Y59_I),
.I5(RIOB33_X105Y131_IOB_X1Y131_I),
.O5(CLBLM_R_X3Y156_SLICE_X2Y156_BO5),
.O6(CLBLM_R_X3Y156_SLICE_X2Y156_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X3Y156_SLICE_X2Y156_ALUT (
.I0(CLBLM_R_X3Y156_SLICE_X2Y156_BO6),
.I1(CLBLM_R_X3Y157_SLICE_X2Y157_BO6),
.I2(CLBLM_R_X3Y155_SLICE_X2Y155_AO6),
.I3(CLBLL_L_X4Y157_SLICE_X5Y157_BO6),
.I4(CLBLM_R_X3Y154_SLICE_X2Y154_CO6),
.I5(CLBLL_L_X2Y153_SLICE_X1Y153_CO6),
.O5(CLBLM_R_X3Y156_SLICE_X2Y156_AO5),
.O6(CLBLM_R_X3Y156_SLICE_X2Y156_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a000a000a000e04)
  ) CLBLM_R_X3Y156_SLICE_X3Y156_DLUT (
.I0(RIOB33_X105Y135_IOB_X1Y135_I),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(CLBLM_L_X16Y156_SLICE_X22Y156_AO6),
.I3(CLBLM_R_X3Y156_SLICE_X3Y156_AO6),
.I4(CLBLL_L_X4Y157_SLICE_X4Y157_AO6),
.I5(RIOB33_X105Y135_IOB_X1Y136_I),
.O5(CLBLM_R_X3Y156_SLICE_X3Y156_DO5),
.O6(CLBLM_R_X3Y156_SLICE_X3Y156_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffae)
  ) CLBLM_R_X3Y156_SLICE_X3Y156_CLUT (
.I0(CLBLM_R_X3Y157_SLICE_X3Y157_AO6),
.I1(CLBLL_L_X4Y152_SLICE_X5Y152_AQ),
.I2(CLBLM_R_X3Y157_SLICE_X2Y157_AO5),
.I3(CLBLL_L_X4Y156_SLICE_X4Y156_DO6),
.I4(CLBLM_R_X3Y157_SLICE_X3Y157_BO6),
.I5(CLBLM_R_X3Y154_SLICE_X2Y154_BO6),
.O5(CLBLM_R_X3Y156_SLICE_X3Y156_CO5),
.O6(CLBLM_R_X3Y156_SLICE_X3Y156_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X3Y156_SLICE_X3Y156_BLUT (
.I0(CLBLM_R_X3Y155_SLICE_X3Y155_DO6),
.I1(CLBLM_R_X3Y155_SLICE_X3Y155_BO6),
.I2(CLBLM_R_X3Y156_SLICE_X2Y156_AO6),
.I3(CLBLL_L_X4Y156_SLICE_X5Y156_AO6),
.I4(CLBLM_R_X3Y156_SLICE_X3Y156_CO6),
.I5(CLBLM_R_X7Y158_SLICE_X9Y158_DO6),
.O5(CLBLM_R_X3Y156_SLICE_X3Y156_BO5),
.O6(CLBLM_R_X3Y156_SLICE_X3Y156_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h10000000fffdfffd)
  ) CLBLM_R_X3Y156_SLICE_X3Y156_ALUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y156_SLICE_X3Y156_AO5),
.O6(CLBLM_R_X3Y156_SLICE_X3Y156_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000002010000000)
  ) CLBLM_R_X3Y157_SLICE_X2Y157_DLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(CLBLM_R_X3Y158_SLICE_X2Y158_AO5),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X3Y157_SLICE_X2Y157_DO5),
.O6(CLBLM_R_X3Y157_SLICE_X2Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haabaffffaaaaffff)
  ) CLBLM_R_X3Y157_SLICE_X2Y157_CLUT (
.I0(RIOB33_X105Y129_IOB_X1Y129_I),
.I1(CLBLL_L_X4Y157_SLICE_X4Y157_CO6),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y137_IOB_X1Y137_I),
.I5(RIOB33_X105Y131_IOB_X1Y132_I),
.O5(CLBLM_R_X3Y157_SLICE_X2Y157_CO5),
.O6(CLBLM_R_X3Y157_SLICE_X2Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000400000000000)
  ) CLBLM_R_X3Y157_SLICE_X2Y157_BLUT (
.I0(CLBLL_L_X4Y157_SLICE_X4Y157_CO6),
.I1(CLBLL_L_X4Y155_SLICE_X4Y155_AQ),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(RIOB33_X105Y133_IOB_X1Y134_I),
.O5(CLBLM_R_X3Y157_SLICE_X2Y157_BO5),
.O6(CLBLM_R_X3Y157_SLICE_X2Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff7fffff7fffffff)
  ) CLBLM_R_X3Y157_SLICE_X2Y157_ALUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_R_X3Y158_SLICE_X2Y158_AO6),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y133_IOB_X1Y133_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y157_SLICE_X2Y157_AO5),
.O6(CLBLM_R_X3Y157_SLICE_X2Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffddffccfffdfffc)
  ) CLBLM_R_X3Y157_SLICE_X3Y157_DLUT (
.I0(CLBLL_L_X4Y157_SLICE_X4Y157_BO6),
.I1(CLBLL_L_X4Y157_SLICE_X4Y157_DO6),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(CLBLM_R_X3Y157_SLICE_X3Y157_CO6),
.I4(CLBLM_R_X5Y157_SLICE_X7Y157_CQ),
.I5(CLBLM_R_X3Y157_SLICE_X2Y157_AO6),
.O5(CLBLM_R_X3Y157_SLICE_X3Y157_DO5),
.O6(CLBLM_R_X3Y157_SLICE_X3Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000400000)
  ) CLBLM_R_X3Y157_SLICE_X3Y157_CLUT (
.I0(RIOB33_X105Y133_IOB_X1Y133_I),
.I1(CLBLM_R_X5Y157_SLICE_X7Y157_BQ),
.I2(RIOB33_X105Y133_IOB_X1Y134_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLL_L_X4Y157_SLICE_X4Y157_CO5),
.O5(CLBLM_R_X3Y157_SLICE_X3Y157_CO5),
.O6(CLBLM_R_X3Y157_SLICE_X3Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h001b0011000a0000)
  ) CLBLM_R_X3Y157_SLICE_X3Y157_BLUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(CLBLL_L_X2Y155_SLICE_X1Y155_CO6),
.I2(CLBLL_L_X2Y155_SLICE_X1Y155_CO5),
.I3(CLBLM_R_X3Y158_SLICE_X2Y158_AO5),
.I4(CLBLM_L_X8Y152_SLICE_X10Y152_CQ),
.I5(CLBLM_R_X5Y157_SLICE_X7Y157_CQ),
.O5(CLBLM_R_X3Y157_SLICE_X3Y157_BO5),
.O6(CLBLM_R_X3Y157_SLICE_X3Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000050005c0c)
  ) CLBLM_R_X3Y157_SLICE_X3Y157_ALUT (
.I0(CLBLL_L_X2Y155_SLICE_X1Y155_CO6),
.I1(CLBLM_R_X5Y157_SLICE_X7Y157_BQ),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(CLBLL_L_X2Y155_SLICE_X1Y155_CO5),
.I5(CLBLM_R_X3Y158_SLICE_X2Y158_AO5),
.O5(CLBLM_R_X3Y157_SLICE_X3Y157_AO5),
.O6(CLBLM_R_X3Y157_SLICE_X3Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y158_SLICE_X2Y158_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y158_SLICE_X2Y158_DO5),
.O6(CLBLM_R_X3Y158_SLICE_X2Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y158_SLICE_X2Y158_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y158_SLICE_X2Y158_CO5),
.O6(CLBLM_R_X3Y158_SLICE_X2Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y158_SLICE_X2Y158_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y158_SLICE_X2Y158_BO5),
.O6(CLBLM_R_X3Y158_SLICE_X2Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000020ffffffcf)
  ) CLBLM_R_X3Y158_SLICE_X2Y158_ALUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(RIOB33_X105Y129_IOB_X1Y130_I),
.I2(RIOB33_X105Y137_IOB_X1Y137_I),
.I3(RIOB33_X105Y135_IOB_X1Y135_I),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y158_SLICE_X2Y158_AO5),
.O6(CLBLM_R_X3Y158_SLICE_X2Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y158_SLICE_X3Y158_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y158_SLICE_X3Y158_DO5),
.O6(CLBLM_R_X3Y158_SLICE_X3Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y158_SLICE_X3Y158_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y158_SLICE_X3Y158_CO5),
.O6(CLBLM_R_X3Y158_SLICE_X3Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y158_SLICE_X3Y158_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y158_SLICE_X3Y158_BO5),
.O6(CLBLM_R_X3Y158_SLICE_X3Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y158_SLICE_X3Y158_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y158_SLICE_X3Y158_AO5),
.O6(CLBLM_R_X3Y158_SLICE_X3Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X6Y144_AO6),
.Q(CLBLM_R_X5Y144_SLICE_X6Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y144_SLICE_X6Y144_BO6),
.Q(CLBLM_R_X5Y144_SLICE_X6Y144_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_DLUT (
.I0(CLBLM_R_X5Y146_SLICE_X6Y146_AQ),
.I1(CLBLM_R_X5Y146_SLICE_X6Y146_BQ),
.I2(CLBLM_R_X5Y144_SLICE_X6Y144_BQ),
.I3(CLBLM_R_X5Y146_SLICE_X6Y146_A5Q),
.I4(CLBLM_R_X7Y145_SLICE_X8Y145_AQ),
.I5(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.O5(CLBLM_R_X5Y144_SLICE_X6Y144_DO5),
.O6(CLBLM_R_X5Y144_SLICE_X6Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000088000000)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_CLUT (
.I0(CLBLM_R_X5Y146_SLICE_X6Y146_AQ),
.I1(CLBLM_R_X5Y146_SLICE_X6Y146_A5Q),
.I2(CLBLM_R_X5Y144_SLICE_X6Y144_BQ),
.I3(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I4(CLBLM_R_X7Y145_SLICE_X8Y145_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y144_SLICE_X6Y144_CO5),
.O6(CLBLM_R_X5Y144_SLICE_X6Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000220088)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y144_SLICE_X6Y144_BQ),
.I2(CLBLM_R_X5Y153_SLICE_X7Y153_AQ),
.I3(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I4(CLBLM_R_X5Y144_SLICE_X6Y144_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y144_SLICE_X6Y144_BO5),
.O6(CLBLM_R_X5Y144_SLICE_X6Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000000ff004848)
  ) CLBLM_R_X5Y144_SLICE_X6Y144_ALUT (
.I0(CLBLM_R_X5Y144_SLICE_X6Y144_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X5Y144_SLICE_X6Y144_AQ),
.I3(CLBLM_R_X11Y155_SLICE_X14Y155_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.O5(CLBLM_R_X5Y144_SLICE_X6Y144_AO5),
.O6(CLBLM_R_X5Y144_SLICE_X6Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y144_SLICE_X7Y144_DO5),
.O6(CLBLM_R_X5Y144_SLICE_X7Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y144_SLICE_X7Y144_CO5),
.O6(CLBLM_R_X5Y144_SLICE_X7Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y144_SLICE_X7Y144_BO5),
.O6(CLBLM_R_X5Y144_SLICE_X7Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y144_SLICE_X7Y144_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y144_SLICE_X7Y144_AO5),
.O6(CLBLM_R_X5Y144_SLICE_X7Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y146_SLICE_X6Y146_CO6),
.Q(CLBLM_R_X5Y146_SLICE_X6Y146_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y146_SLICE_X6Y146_AO6),
.Q(CLBLM_R_X5Y146_SLICE_X6Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y146_SLICE_X6Y146_BO6),
.Q(CLBLM_R_X5Y146_SLICE_X6Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y146_SLICE_X6Y146_DO5),
.O6(CLBLM_R_X5Y146_SLICE_X6Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0d1c0c011110000)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_CLUT (
.I0(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y152_SLICE_X8Y152_AQ),
.I3(CLBLM_R_X5Y146_SLICE_X6Y146_A5Q),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y146_SLICE_X6Y146_CO5),
.O6(CLBLM_R_X5Y146_SLICE_X6Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff2800000028)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y146_SLICE_X6Y146_BQ),
.I2(CLBLM_R_X5Y144_SLICE_X6Y144_CO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I5(CLBLM_L_X10Y149_SLICE_X13Y149_BQ),
.O5(CLBLM_R_X5Y146_SLICE_X6Y146_BO5),
.O6(CLBLM_R_X5Y146_SLICE_X6Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hde5acc00fcf0cc00)
  ) CLBLM_R_X5Y146_SLICE_X6Y146_ALUT (
.I0(CLBLM_R_X7Y145_SLICE_X8Y145_AQ),
.I1(CLBLM_R_X5Y147_SLICE_X6Y147_BQ),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y146_SLICE_X6Y146_CO5),
.I5(CLBLM_R_X5Y146_SLICE_X6Y146_A5Q),
.O5(CLBLM_R_X5Y146_SLICE_X6Y146_AO5),
.O6(CLBLM_R_X5Y146_SLICE_X6Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y146_SLICE_X7Y146_DO5),
.O6(CLBLM_R_X5Y146_SLICE_X7Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y146_SLICE_X7Y146_CO5),
.O6(CLBLM_R_X5Y146_SLICE_X7Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y146_SLICE_X7Y146_BO5),
.O6(CLBLM_R_X5Y146_SLICE_X7Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y146_SLICE_X7Y146_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y146_SLICE_X7Y146_AO5),
.O6(CLBLM_R_X5Y146_SLICE_X7Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X6Y147_AO6),
.Q(CLBLM_R_X5Y147_SLICE_X6Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X6Y147_BO6),
.Q(CLBLM_R_X5Y147_SLICE_X6Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y147_SLICE_X6Y147_DO5),
.O6(CLBLM_R_X5Y147_SLICE_X6Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y147_SLICE_X6Y147_CO5),
.O6(CLBLM_R_X5Y147_SLICE_X6Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0f000fff0c000c)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y147_SLICE_X6Y147_BQ),
.I2(CLBLL_L_X4Y147_SLICE_X4Y147_BO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y155_SLICE_X11Y155_BQ),
.I5(CLBLM_R_X5Y148_SLICE_X7Y148_A5Q),
.O5(CLBLM_R_X5Y147_SLICE_X6Y147_BO5),
.O6(CLBLM_R_X5Y147_SLICE_X6Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0aa0cccca0a0)
  ) CLBLM_R_X5Y147_SLICE_X6Y147_ALUT (
.I0(CLBLM_R_X7Y152_SLICE_X8Y152_BO5),
.I1(CLBLM_R_X5Y149_SLICE_X6Y149_AQ),
.I2(CLBLM_R_X5Y147_SLICE_X6Y147_AQ),
.I3(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y146_SLICE_X5Y146_AO5),
.O5(CLBLM_R_X5Y147_SLICE_X6Y147_AO5),
.O6(CLBLM_R_X5Y147_SLICE_X6Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X7Y147_CO5),
.Q(CLBLM_R_X5Y147_SLICE_X7Y147_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X7Y147_AO6),
.Q(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X7Y147_BO6),
.Q(CLBLM_R_X5Y147_SLICE_X7Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y147_SLICE_X7Y147_CO6),
.Q(CLBLM_R_X5Y147_SLICE_X7Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y147_SLICE_X7Y147_DO5),
.O6(CLBLM_R_X5Y147_SLICE_X7Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaa00ccf0ccf0)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_CLUT (
.I0(CLBLM_R_X5Y148_SLICE_X7Y148_AQ),
.I1(CLBLM_R_X5Y147_SLICE_X7Y147_CQ),
.I2(CLBLM_R_X7Y148_SLICE_X8Y148_CQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y127_IOB_X1Y127_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y147_SLICE_X7Y147_CO5),
.O6(CLBLM_R_X5Y147_SLICE_X7Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000ffee3322)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_BLUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X5Y147_SLICE_X6Y147_AQ),
.I5(CLBLM_L_X10Y150_SLICE_X12Y150_CO6),
.O5(CLBLM_R_X5Y147_SLICE_X7Y147_BO5),
.O6(CLBLM_R_X5Y147_SLICE_X7Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeaaeeaaeca0eca0)
  ) CLBLM_R_X5Y147_SLICE_X7Y147_ALUT (
.I0(CLBLM_R_X5Y152_SLICE_X6Y152_CO6),
.I1(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I2(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X5Y148_SLICE_X6Y148_A5Q),
.O5(CLBLM_R_X5Y147_SLICE_X7Y147_AO5),
.O6(CLBLM_R_X5Y147_SLICE_X7Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_L_X8Y148_SLICE_X11Y148_DO5),
.Q(CLBLM_R_X5Y148_SLICE_X6Y148_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y148_SLICE_X6Y148_AO6),
.Q(CLBLM_R_X5Y148_SLICE_X6Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y148_SLICE_X6Y148_BO6),
.Q(CLBLM_R_X5Y148_SLICE_X6Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0333ffff0fffffff)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y150_SLICE_X5Y150_BQ),
.I2(CLBLM_R_X5Y148_SLICE_X6Y148_AQ),
.I3(CLBLM_R_X5Y148_SLICE_X6Y148_BQ),
.I4(CLBLM_R_X5Y149_SLICE_X7Y149_CQ),
.I5(CLBLL_L_X4Y150_SLICE_X5Y150_AQ),
.O5(CLBLM_R_X5Y148_SLICE_X6Y148_DO5),
.O6(CLBLM_R_X5Y148_SLICE_X6Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff153f7fff7fff)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_CLUT (
.I0(CLBLM_R_X7Y148_SLICE_X8Y148_CQ),
.I1(CLBLM_R_X7Y148_SLICE_X8Y148_A5Q),
.I2(CLBLM_L_X10Y149_SLICE_X12Y149_BQ),
.I3(CLBLL_L_X4Y148_SLICE_X5Y148_DQ),
.I4(CLBLM_R_X5Y148_SLICE_X6Y148_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y148_SLICE_X6Y148_CO5),
.O6(CLBLM_R_X5Y148_SLICE_X6Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30cc00cc00fc30)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y149_SLICE_X12Y149_DO5),
.I3(CLBLM_R_X5Y158_SLICE_X6Y158_BQ),
.I4(CLBLM_R_X5Y148_SLICE_X6Y148_CO5),
.I5(CLBLM_R_X5Y148_SLICE_X6Y148_BQ),
.O5(CLBLM_R_X5Y148_SLICE_X6Y148_BO5),
.O6(CLBLM_R_X5Y148_SLICE_X6Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hec20dc10ec20ec20)
  ) CLBLM_R_X5Y148_SLICE_X6Y148_ALUT (
.I0(CLBLM_R_X5Y148_SLICE_X6Y148_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y149_SLICE_X12Y149_DO5),
.I3(CLBLM_L_X10Y149_SLICE_X12Y149_CQ),
.I4(CLBLM_R_X5Y148_SLICE_X6Y148_CO5),
.I5(CLBLM_R_X5Y148_SLICE_X6Y148_BQ),
.O5(CLBLM_R_X5Y148_SLICE_X6Y148_AO5),
.O6(CLBLM_R_X5Y148_SLICE_X6Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X7Y149_DO5),
.Q(CLBLM_R_X5Y148_SLICE_X7Y148_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y148_SLICE_X7Y148_BO5),
.Q(CLBLM_R_X5Y148_SLICE_X7Y148_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y148_SLICE_X7Y148_AO6),
.Q(CLBLM_R_X5Y148_SLICE_X7Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y148_SLICE_X7Y148_BO6),
.Q(CLBLM_R_X5Y148_SLICE_X7Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffdfff)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_DLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(RIOB33_X105Y135_IOB_X1Y135_I),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(RIOB33_X105Y137_IOB_X1Y137_I),
.I4(RIOB33_X105Y129_IOB_X1Y129_I),
.I5(RIOB33_X105Y129_IOB_X1Y130_I),
.O5(CLBLM_R_X5Y148_SLICE_X7Y148_DO5),
.O6(CLBLM_R_X5Y148_SLICE_X7Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ac0000000000)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_CLUT (
.I0(CLBLM_R_X5Y149_SLICE_X7Y149_AQ),
.I1(CLBLM_L_X8Y148_SLICE_X10Y148_AQ),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(RIOB33_X105Y133_IOB_X1Y133_I),
.I4(CLBLM_R_X5Y148_SLICE_X7Y148_DO6),
.I5(RIOB33_X105Y133_IOB_X1Y134_I),
.O5(CLBLM_R_X5Y148_SLICE_X7Y148_CO5),
.O6(CLBLM_R_X5Y148_SLICE_X7Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaf0ccf0ccf0)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_BLUT (
.I0(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.I1(CLBLM_L_X8Y148_SLICE_X10Y148_AQ),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y148_SLICE_X7Y148_BO5),
.O6(CLBLM_R_X5Y148_SLICE_X7Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00fe54fe54fe54)
  ) CLBLM_R_X5Y148_SLICE_X7Y148_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y148_SLICE_X10Y148_BQ),
.I2(CLBLM_R_X5Y148_SLICE_X7Y148_AQ),
.I3(CLBLM_R_X7Y147_SLICE_X9Y147_BQ),
.I4(CLBLM_L_X10Y151_SLICE_X12Y151_CQ),
.I5(CLBLL_L_X4Y151_SLICE_X4Y151_BQ),
.O5(CLBLM_R_X5Y148_SLICE_X7Y148_AO5),
.O6(CLBLM_R_X5Y148_SLICE_X7Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X6Y149_AO5),
.Q(CLBLM_R_X5Y149_SLICE_X6Y149_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X6Y149_BO5),
.Q(CLBLM_R_X5Y149_SLICE_X6Y149_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X6Y149_AO6),
.Q(CLBLM_R_X5Y149_SLICE_X6Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X6Y149_BO6),
.Q(CLBLM_R_X5Y149_SLICE_X6Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_DLUT (
.I0(CLBLM_R_X5Y148_SLICE_X6Y148_BQ),
.I1(CLBLM_R_X7Y148_SLICE_X8Y148_A5Q),
.I2(CLBLM_R_X5Y148_SLICE_X6Y148_AQ),
.I3(CLBLL_L_X4Y148_SLICE_X5Y148_DQ),
.I4(CLBLM_L_X10Y149_SLICE_X12Y149_BQ),
.I5(CLBLM_R_X7Y148_SLICE_X8Y148_CQ),
.O5(CLBLM_R_X5Y149_SLICE_X6Y149_DO5),
.O6(CLBLM_R_X5Y149_SLICE_X6Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f04488888888)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_CLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I2(CLBLM_L_X10Y149_SLICE_X13Y149_A5Q),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y149_SLICE_X8Y149_DO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y149_SLICE_X6Y149_CO5),
.O6(CLBLM_R_X5Y149_SLICE_X6Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0c0bb88bb88)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_BLUT (
.I0(CLBLM_R_X7Y151_SLICE_X9Y151_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X8Y147_SLICE_X11Y147_BQ),
.I3(CLBLM_L_X8Y147_SLICE_X11Y147_CO6),
.I4(CLBLL_L_X4Y153_SLICE_X4Y153_BO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y149_SLICE_X6Y149_BO5),
.O6(CLBLM_R_X5Y149_SLICE_X6Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdddd8888fa50fa50)
  ) CLBLM_R_X5Y149_SLICE_X6Y149_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y150_SLICE_X6Y150_BQ),
.I2(CLBLL_L_X4Y148_SLICE_X4Y148_AQ),
.I3(CLBLM_R_X5Y147_SLICE_X7Y147_BQ),
.I4(CLBLM_R_X5Y148_SLICE_X6Y148_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y149_SLICE_X6Y149_AO5),
.O6(CLBLM_R_X5Y149_SLICE_X6Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X6Y149_CO6),
.Q(CLBLM_R_X5Y149_SLICE_X7Y149_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X7Y149_AO6),
.Q(CLBLM_R_X5Y149_SLICE_X7Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X7Y149_BO6),
.Q(CLBLM_R_X5Y149_SLICE_X7Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y149_SLICE_X7Y149_CO6),
.Q(CLBLM_R_X5Y149_SLICE_X7Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00cc00fafa5050)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y149_SLICE_X15Y149_A5Q),
.I2(CLBLL_L_X4Y150_SLICE_X5Y150_BQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y149_SLICE_X7Y149_DO5),
.O6(CLBLM_R_X5Y149_SLICE_X7Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1e4b1e4a0a0a0a0)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y149_SLICE_X7Y149_CQ),
.I2(CLBLM_L_X8Y155_SLICE_X10Y155_B5Q),
.I3(CLBLL_L_X4Y149_SLICE_X5Y149_BO5),
.I4(1'b1),
.I5(CLBLM_L_X10Y149_SLICE_X12Y149_DO5),
.O5(CLBLM_R_X5Y149_SLICE_X7Y149_CO5),
.O6(CLBLM_R_X5Y149_SLICE_X7Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffee00ee00ee00)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_BLUT (
.I0(CLBLM_L_X8Y151_SLICE_X10Y151_CQ),
.I1(CLBLM_R_X5Y149_SLICE_X7Y149_BQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y152_SLICE_X6Y152_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y149_SLICE_X16Y149_BQ),
.O5(CLBLM_R_X5Y149_SLICE_X7Y149_BO5),
.O6(CLBLM_R_X5Y149_SLICE_X7Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff001f1f1010)
  ) CLBLM_R_X5Y149_SLICE_X7Y149_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLL_L_X4Y153_SLICE_X4Y153_AO6),
.I2(CLBLM_R_X5Y149_SLICE_X6Y149_CO5),
.I3(CLBLM_R_X7Y148_SLICE_X8Y148_BQ),
.I4(CLBLM_R_X5Y149_SLICE_X7Y149_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y149_SLICE_X7Y149_AO5),
.O6(CLBLM_R_X5Y149_SLICE_X7Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y150_SLICE_X6Y150_AO6),
.Q(CLBLM_R_X5Y150_SLICE_X6Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y150_SLICE_X6Y150_BO6),
.Q(CLBLM_R_X5Y150_SLICE_X6Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y150_SLICE_X6Y150_CO6),
.Q(CLBLM_R_X5Y150_SLICE_X6Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y150_SLICE_X6Y150_DO6),
.Q(CLBLM_R_X5Y150_SLICE_X6Y150_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fcfcff005454)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_DLUT (
.I0(CLBLM_L_X10Y150_SLICE_X12Y150_A5Q),
.I1(CLBLM_L_X8Y148_SLICE_X10Y148_BQ),
.I2(CLBLM_R_X5Y150_SLICE_X6Y150_DQ),
.I3(CLBLM_L_X8Y148_SLICE_X11Y148_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y155_SLICE_X16Y155_CO6),
.O5(CLBLM_R_X5Y150_SLICE_X6Y150_DO5),
.O6(CLBLM_R_X5Y150_SLICE_X6Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffccf0f05544)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_CLUT (
.I0(CLBLM_L_X10Y150_SLICE_X12Y150_A5Q),
.I1(CLBLM_R_X5Y150_SLICE_X6Y150_CQ),
.I2(CLBLM_L_X8Y148_SLICE_X10Y148_BQ),
.I3(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y155_SLICE_X16Y155_CO6),
.O5(CLBLM_R_X5Y150_SLICE_X6Y150_CO5),
.O6(CLBLM_R_X5Y150_SLICE_X6Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaffaac0aacc)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_BLUT (
.I0(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.I1(CLBLM_R_X5Y150_SLICE_X6Y150_BQ),
.I2(CLBLM_L_X12Y155_SLICE_X16Y155_CO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y150_SLICE_X12Y150_A5Q),
.I5(CLBLM_L_X8Y149_SLICE_X10Y149_AQ),
.O5(CLBLM_R_X5Y150_SLICE_X6Y150_BO5),
.O6(CLBLM_R_X5Y150_SLICE_X6Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff110011ff220022)
  ) CLBLM_R_X5Y150_SLICE_X6Y150_ALUT (
.I0(CLBLM_R_X5Y150_SLICE_X7Y150_BQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y149_SLICE_X6Y149_A5Q),
.I5(CLBLM_R_X7Y150_SLICE_X9Y150_AO5),
.O5(CLBLM_R_X5Y150_SLICE_X6Y150_AO5),
.O6(CLBLM_R_X5Y150_SLICE_X6Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y150_SLICE_X7Y150_AO5),
.Q(CLBLM_R_X5Y150_SLICE_X7Y150_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y150_SLICE_X7Y150_AO6),
.Q(CLBLM_R_X5Y150_SLICE_X7Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y150_SLICE_X7Y150_BO6),
.Q(CLBLM_R_X5Y150_SLICE_X7Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y150_SLICE_X7Y150_CO6),
.Q(CLBLM_R_X5Y150_SLICE_X7Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc000c00000000000)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y148_SLICE_X6Y148_A5Q),
.I2(CLBLM_L_X8Y151_SLICE_X10Y151_CQ),
.I3(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y150_SLICE_X12Y150_CQ),
.O5(CLBLM_R_X5Y150_SLICE_X7Y150_DO5),
.O6(CLBLM_R_X5Y150_SLICE_X7Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ccccaaaa)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_CLUT (
.I0(CLBLM_R_X5Y151_SLICE_X6Y151_C5Q),
.I1(CLBLM_R_X5Y150_SLICE_X7Y150_CQ),
.I2(1'b1),
.I3(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I4(CLBLL_L_X4Y147_SLICE_X4Y147_BO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y150_SLICE_X7Y150_CO5),
.O6(CLBLM_R_X5Y150_SLICE_X7Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000f303fc0c)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y150_SLICE_X8Y150_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y149_SLICE_X4Y149_BQ),
.I4(CLBLM_R_X7Y150_SLICE_X9Y150_AO6),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y150_SLICE_X7Y150_BO5),
.O6(CLBLM_R_X5Y150_SLICE_X7Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aaf0f0ccf0cc)
  ) CLBLM_R_X5Y150_SLICE_X7Y150_ALUT (
.I0(CLBLM_R_X5Y156_SLICE_X7Y156_AQ),
.I1(CLBLL_L_X4Y150_SLICE_X5Y150_AQ),
.I2(CLBLM_R_X5Y150_SLICE_X7Y150_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y150_SLICE_X7Y150_AO5),
.O6(CLBLM_R_X5Y150_SLICE_X7Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y151_SLICE_X6Y151_CO5),
.Q(CLBLM_R_X5Y151_SLICE_X6Y151_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y151_SLICE_X6Y151_AO6),
.Q(CLBLM_R_X5Y151_SLICE_X6Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y151_SLICE_X6Y151_BO6),
.Q(CLBLM_R_X5Y151_SLICE_X6Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y151_SLICE_X6Y151_CO6),
.Q(CLBLM_R_X5Y151_SLICE_X6Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y151_SLICE_X6Y151_DO6),
.Q(CLBLM_R_X5Y151_SLICE_X6Y151_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc50ccfacc50cc50)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_DLUT (
.I0(CLBLM_R_X5Y149_SLICE_X6Y149_CO5),
.I1(CLBLM_L_X12Y149_SLICE_X17Y149_A5Q),
.I2(CLBLM_R_X5Y151_SLICE_X6Y151_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLL_L_X4Y154_SLICE_X4Y154_BO6),
.O5(CLBLM_R_X5Y151_SLICE_X6Y151_DO5),
.O6(CLBLM_R_X5Y151_SLICE_X6Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5500f0f0cccc)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y148_SLICE_X6Y148_AQ),
.I2(CLBLM_R_X7Y153_SLICE_X8Y153_CQ),
.I3(CLBLM_R_X7Y153_SLICE_X8Y153_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y151_SLICE_X6Y151_CO5),
.O6(CLBLM_R_X5Y151_SLICE_X6Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcfffc000cf00c0)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y151_SLICE_X6Y151_BQ),
.I2(CLBLM_R_X5Y152_SLICE_X6Y152_CO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y150_SLICE_X7Y150_BQ),
.I5(CLBLM_R_X5Y150_SLICE_X6Y150_CQ),
.O5(CLBLM_R_X5Y151_SLICE_X6Y151_BO5),
.O6(CLBLM_R_X5Y151_SLICE_X6Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5554555400540054)
  ) CLBLM_R_X5Y151_SLICE_X6Y151_ALUT (
.I0(CLBLM_R_X5Y152_SLICE_X6Y152_CO6),
.I1(CLBLM_R_X7Y150_SLICE_X8Y150_BQ),
.I2(CLBLM_R_X5Y151_SLICE_X6Y151_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.O5(CLBLM_R_X5Y151_SLICE_X6Y151_AO5),
.O6(CLBLM_R_X5Y151_SLICE_X6Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y151_SLICE_X7Y151_AO6),
.Q(CLBLM_R_X5Y151_SLICE_X7Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y151_SLICE_X7Y151_BO6),
.Q(CLBLM_R_X5Y151_SLICE_X7Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y151_SLICE_X7Y151_CO6),
.Q(CLBLM_R_X5Y151_SLICE_X7Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y151_SLICE_X7Y151_DO6),
.Q(CLBLM_R_X5Y151_SLICE_X7Y151_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbaba1010feba5410)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y149_SLICE_X6Y149_CO5),
.I2(CLBLM_R_X5Y151_SLICE_X7Y151_DQ),
.I3(CLBLL_L_X4Y154_SLICE_X5Y154_BO6),
.I4(CLBLM_R_X5Y150_SLICE_X7Y150_BQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y151_SLICE_X7Y151_DO5),
.O6(CLBLM_R_X5Y151_SLICE_X7Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hae04ae04ae04ae04)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y151_SLICE_X7Y151_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X8Y151_SLICE_X10Y151_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y151_SLICE_X7Y151_CO5),
.O6(CLBLM_R_X5Y151_SLICE_X7Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff005c5cff000c0c)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X5Y151_SLICE_X7Y151_BQ),
.I2(CLBLM_R_X5Y149_SLICE_X6Y149_CO5),
.I3(CLBLM_L_X12Y154_SLICE_X16Y154_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X3Y156_SLICE_X2Y156_DO6),
.O5(CLBLM_R_X5Y151_SLICE_X7Y151_BO5),
.O6(CLBLM_R_X5Y151_SLICE_X7Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddfc1130fcfc3030)
  ) CLBLM_R_X5Y151_SLICE_X7Y151_ALUT (
.I0(CLBLM_R_X3Y152_SLICE_X3Y152_BO5),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y151_SLICE_X7Y151_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLL_L_X4Y151_SLICE_X4Y151_BQ),
.I5(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.O5(CLBLM_R_X5Y151_SLICE_X7Y151_AO5),
.O6(CLBLM_R_X5Y151_SLICE_X7Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X6Y152_AO6),
.Q(CLBLM_R_X5Y152_SLICE_X6Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X6Y152_BO6),
.Q(CLBLM_R_X5Y152_SLICE_X6Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000030aa30)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_DLUT (
.I0(CLBLM_R_X5Y150_SLICE_X6Y150_BQ),
.I1(CLBLL_L_X2Y155_SLICE_X1Y155_CO6),
.I2(CLBLM_R_X5Y151_SLICE_X6Y151_BQ),
.I3(RIOB33_X105Y135_IOB_X1Y136_I),
.I4(CLBLM_R_X3Y156_SLICE_X3Y156_AO5),
.I5(CLBLM_R_X3Y158_SLICE_X2Y158_AO5),
.O5(CLBLM_R_X5Y152_SLICE_X6Y152_DO5),
.O6(CLBLM_R_X5Y152_SLICE_X6Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h44404444ccc0cccc)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_R_X5Y154_SLICE_X6Y154_AQ),
.I4(CLBLM_L_X12Y149_SLICE_X16Y149_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y152_SLICE_X6Y152_CO5),
.O6(CLBLM_R_X5Y152_SLICE_X6Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0afa0af000f000)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_BLUT (
.I0(CLBLM_R_X7Y149_SLICE_X8Y149_CQ),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y152_SLICE_X5Y152_AQ),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y152_SLICE_X6Y152_BO5),
.O6(CLBLM_R_X5Y152_SLICE_X6Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000fa0afa0a)
  ) CLBLM_R_X5Y152_SLICE_X6Y152_ALUT (
.I0(CLBLM_L_X10Y150_SLICE_X13Y150_CQ),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y152_SLICE_X7Y152_BQ),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y152_SLICE_X6Y152_AO5),
.O6(CLBLM_R_X5Y152_SLICE_X6Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X7Y152_AO6),
.Q(CLBLM_R_X5Y152_SLICE_X7Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X7Y152_BO6),
.Q(CLBLM_R_X5Y152_SLICE_X7Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X7Y152_CO6),
.Q(CLBLM_R_X5Y152_SLICE_X7Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y152_SLICE_X7Y152_DO6),
.Q(CLBLM_R_X5Y152_SLICE_X7Y152_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000fcfc0c0c)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y152_SLICE_X12Y152_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X5Y151_SLICE_X7Y151_DQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y152_SLICE_X7Y152_DO5),
.O6(CLBLM_R_X5Y152_SLICE_X7Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0003300cc)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y150_SLICE_X8Y150_CO6),
.I2(CLBLM_R_X5Y152_SLICE_X7Y152_DQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X5Y157_SLICE_X7Y157_DQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y152_SLICE_X7Y152_CO5),
.O6(CLBLM_R_X5Y152_SLICE_X7Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haafcaafcaa0caa0c)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_BLUT (
.I0(CLBLM_R_X7Y149_SLICE_X8Y149_CQ),
.I1(CLBLM_R_X5Y152_SLICE_X7Y152_BQ),
.I2(CLBLM_R_X5Y152_SLICE_X6Y152_CO5),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_L_X10Y152_SLICE_X12Y152_AQ),
.O5(CLBLM_R_X5Y152_SLICE_X7Y152_BO5),
.O6(CLBLM_R_X5Y152_SLICE_X7Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5511541055115410)
  ) CLBLM_R_X5Y152_SLICE_X7Y152_ALUT (
.I0(CLBLM_R_X5Y152_SLICE_X6Y152_CO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X5Y152_SLICE_X7Y152_AQ),
.I3(CLBLM_R_X5Y149_SLICE_X7Y149_AQ),
.I4(CLBLM_L_X8Y151_SLICE_X11Y151_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y152_SLICE_X7Y152_AO5),
.O6(CLBLM_R_X5Y152_SLICE_X7Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y153_SLICE_X6Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y153_SLICE_X6Y153_AO6),
.Q(CLBLM_R_X5Y153_SLICE_X6Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff5d5d0c0c)
  ) CLBLM_R_X5Y153_SLICE_X6Y153_DLUT (
.I0(CLBLM_R_X3Y157_SLICE_X2Y157_AO6),
.I1(CLBLM_R_X5Y147_SLICE_X7Y147_AQ),
.I2(CLBLM_R_X3Y154_SLICE_X3Y154_AO6),
.I3(1'b1),
.I4(RIOB33_X105Y111_IOB_X1Y111_I),
.I5(CLBLM_R_X5Y152_SLICE_X6Y152_DO6),
.O5(CLBLM_R_X5Y153_SLICE_X6Y153_DO5),
.O6(CLBLM_R_X5Y153_SLICE_X6Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccefccefccecccec)
  ) CLBLM_R_X5Y153_SLICE_X6Y153_CLUT (
.I0(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.I1(CLBLM_R_X5Y148_SLICE_X7Y148_CO6),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLM_R_X3Y153_SLICE_X3Y153_AO5),
.I4(1'b1),
.I5(CLBLM_L_X8Y157_SLICE_X10Y157_CQ),
.O5(CLBLM_R_X5Y153_SLICE_X6Y153_CO5),
.O6(CLBLM_R_X5Y153_SLICE_X6Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffbfffdffff)
  ) CLBLM_R_X5Y153_SLICE_X6Y153_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(RIOB33_X105Y133_IOB_X1Y134_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(CLBLL_L_X4Y157_SLICE_X4Y157_CO5),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y153_SLICE_X6Y153_BO5),
.O6(CLBLM_R_X5Y153_SLICE_X6Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000022202220)
  ) CLBLM_R_X5Y153_SLICE_X6Y153_ALUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X5Y153_SLICE_X6Y153_AQ),
.I3(CLBLM_L_X12Y150_SLICE_X16Y150_CQ),
.I4(CLBLL_L_X4Y151_SLICE_X5Y151_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y153_SLICE_X6Y153_AO5),
.O6(CLBLM_R_X5Y153_SLICE_X6Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y153_SLICE_X7Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y153_SLICE_X7Y153_AO6),
.Q(CLBLM_R_X5Y153_SLICE_X7Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffeeffeeff)
  ) CLBLM_R_X5Y153_SLICE_X7Y153_DLUT (
.I0(CLBLM_R_X5Y154_SLICE_X6Y154_AQ),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(1'b1),
.I3(CLBLM_L_X12Y149_SLICE_X16Y149_CQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y152_SLICE_X12Y152_AQ),
.O5(CLBLM_R_X5Y153_SLICE_X7Y153_DO5),
.O6(CLBLM_R_X5Y153_SLICE_X7Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000001)
  ) CLBLM_R_X5Y153_SLICE_X7Y153_CLUT (
.I0(CLBLM_R_X5Y157_SLICE_X7Y157_DQ),
.I1(CLBLM_R_X7Y150_SLICE_X8Y150_BQ),
.I2(CLBLM_R_X7Y153_SLICE_X9Y153_DO6),
.I3(CLBLM_R_X5Y150_SLICE_X7Y150_BQ),
.I4(CLBLM_R_X5Y153_SLICE_X7Y153_DO6),
.I5(CLBLM_R_X5Y152_SLICE_X6Y152_AQ),
.O5(CLBLM_R_X5Y153_SLICE_X7Y153_CO5),
.O6(CLBLM_R_X5Y153_SLICE_X7Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfffffffffffffff)
  ) CLBLM_R_X5Y153_SLICE_X7Y153_BLUT (
.I0(CLBLM_R_X5Y152_SLICE_X7Y152_DQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y150_SLICE_X11Y150_AQ),
.I3(CLBLM_R_X7Y156_SLICE_X9Y156_BQ),
.I4(CLBLM_L_X8Y153_SLICE_X11Y153_DQ),
.I5(CLBLM_R_X5Y152_SLICE_X7Y152_CQ),
.O5(CLBLM_R_X5Y153_SLICE_X7Y153_BO5),
.O6(CLBLM_R_X5Y153_SLICE_X7Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa30ff3030)
  ) CLBLM_R_X5Y153_SLICE_X7Y153_ALUT (
.I0(CLBLM_L_X12Y154_SLICE_X16Y154_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X5Y153_SLICE_X7Y153_AQ),
.I3(CLBLM_R_X5Y153_SLICE_X7Y153_BO6),
.I4(CLBLM_R_X5Y153_SLICE_X7Y153_CO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X5Y153_SLICE_X7Y153_AO5),
.O6(CLBLM_R_X5Y153_SLICE_X7Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y154_SLICE_X6Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y154_SLICE_X6Y154_AO6),
.Q(CLBLM_R_X5Y154_SLICE_X6Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aaaaf0f0fafa)
  ) CLBLM_R_X5Y154_SLICE_X6Y154_DLUT (
.I0(CLBLM_R_X5Y154_SLICE_X7Y154_AQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y151_SLICE_X5Y151_AQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y157_SLICE_X4Y157_BO5),
.I5(CLBLM_R_X5Y153_SLICE_X6Y153_BO6),
.O5(CLBLM_R_X5Y154_SLICE_X6Y154_DO5),
.O6(CLBLM_R_X5Y154_SLICE_X6Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4444ff44f4f4fff4)
  ) CLBLM_R_X5Y154_SLICE_X6Y154_CLUT (
.I0(CLBLM_R_X3Y157_SLICE_X2Y157_AO6),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(CLBLM_R_X7Y154_SLICE_X9Y154_AQ),
.I3(CLBLM_R_X5Y150_SLICE_X6Y150_CQ),
.I4(CLBLL_L_X4Y156_SLICE_X4Y156_CO6),
.I5(CLBLM_R_X5Y153_SLICE_X6Y153_BO6),
.O5(CLBLM_R_X5Y154_SLICE_X6Y154_CO5),
.O6(CLBLM_R_X5Y154_SLICE_X6Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3fbf0faf33bb00aa)
  ) CLBLM_R_X5Y154_SLICE_X6Y154_BLUT (
.I0(CLBLM_R_X11Y155_SLICE_X14Y155_AQ),
.I1(CLBLL_L_X2Y155_SLICE_X1Y155_BO5),
.I2(CLBLM_R_X3Y157_SLICE_X2Y157_AO5),
.I3(CLBLM_R_X3Y154_SLICE_X3Y154_AO5),
.I4(CLBLL_L_X4Y148_SLICE_X5Y148_AQ),
.I5(CLBLM_R_X5Y151_SLICE_X6Y151_DQ),
.O5(CLBLM_R_X5Y154_SLICE_X6Y154_BO5),
.O6(CLBLM_R_X5Y154_SLICE_X6Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00c4c4ff00c0c0)
  ) CLBLM_R_X5Y154_SLICE_X6Y154_ALUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X5Y154_SLICE_X6Y154_AQ),
.I3(CLBLM_R_X5Y151_SLICE_X6Y151_DQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y149_SLICE_X16Y149_CQ),
.O5(CLBLM_R_X5Y154_SLICE_X6Y154_AO5),
.O6(CLBLM_R_X5Y154_SLICE_X6Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y154_SLICE_X7Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y154_SLICE_X7Y154_AO6),
.Q(CLBLM_R_X5Y154_SLICE_X7Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff75307530)
  ) CLBLM_R_X5Y154_SLICE_X7Y154_DLUT (
.I0(CLBLL_L_X2Y155_SLICE_X1Y155_BO5),
.I1(CLBLM_R_X3Y157_SLICE_X2Y157_AO5),
.I2(CLBLM_R_X5Y151_SLICE_X7Y151_AQ),
.I3(CLBLM_R_X5Y148_SLICE_X7Y148_AQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y154_SLICE_X7Y154_BO6),
.O5(CLBLM_R_X5Y154_SLICE_X7Y154_DO5),
.O6(CLBLM_R_X5Y154_SLICE_X7Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fdf0fcf55dd00cc)
  ) CLBLM_R_X5Y154_SLICE_X7Y154_CLUT (
.I0(CLBLL_L_X2Y155_SLICE_X1Y155_BO5),
.I1(CLBLM_R_X5Y155_SLICE_X7Y155_AQ),
.I2(CLBLM_R_X3Y153_SLICE_X3Y153_AO6),
.I3(CLBLM_R_X3Y154_SLICE_X3Y154_AO5),
.I4(CLBLM_R_X7Y149_SLICE_X9Y149_BQ),
.I5(CLBLM_L_X10Y154_SLICE_X12Y154_AQ),
.O5(CLBLM_R_X5Y154_SLICE_X7Y154_CO5),
.O6(CLBLM_R_X5Y154_SLICE_X7Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000003020100)
  ) CLBLM_R_X5Y154_SLICE_X7Y154_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y131_I),
.I1(CLBLL_L_X4Y157_SLICE_X4Y157_CO5),
.I2(RIOB33_X105Y131_IOB_X1Y132_I),
.I3(CLBLM_R_X11Y153_SLICE_X15Y153_BQ),
.I4(CLBLM_L_X8Y153_SLICE_X11Y153_AQ),
.I5(CLBLL_L_X4Y157_SLICE_X4Y157_AO5),
.O5(CLBLM_R_X5Y154_SLICE_X7Y154_BO5),
.O6(CLBLM_R_X5Y154_SLICE_X7Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0ccffccf0cc00)
  ) CLBLM_R_X5Y154_SLICE_X7Y154_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y146_SLICE_X12Y146_C5Q),
.I2(CLBLM_R_X5Y154_SLICE_X7Y154_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y152_SLICE_X6Y152_CO5),
.I5(CLBLM_R_X5Y152_SLICE_X6Y152_AQ),
.O5(CLBLM_R_X5Y154_SLICE_X7Y154_AO5),
.O6(CLBLM_R_X5Y154_SLICE_X7Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y155_SLICE_X6Y155_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y155_SLICE_X6Y155_AO6),
.Q(CLBLM_R_X5Y155_SLICE_X6Y155_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffaafffa)
  ) CLBLM_R_X5Y155_SLICE_X6Y155_DLUT (
.I0(CLBLM_R_X7Y155_SLICE_X9Y155_DO6),
.I1(1'b1),
.I2(CLBLL_L_X4Y156_SLICE_X4Y156_CO5),
.I3(CLBLM_R_X5Y155_SLICE_X6Y155_CO6),
.I4(CLBLM_R_X3Y154_SLICE_X3Y154_DO6),
.I5(CLBLM_R_X5Y156_SLICE_X6Y156_BO6),
.O5(CLBLM_R_X5Y155_SLICE_X6Y155_DO5),
.O6(CLBLM_R_X5Y155_SLICE_X6Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffdfcfffffddcc)
  ) CLBLM_R_X5Y155_SLICE_X6Y155_CLUT (
.I0(CLBLM_R_X3Y157_SLICE_X2Y157_AO6),
.I1(CLBLL_L_X4Y155_SLICE_X5Y155_CO6),
.I2(CLBLL_L_X4Y156_SLICE_X4Y156_CO5),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(CLBLL_L_X4Y156_SLICE_X5Y156_DO6),
.I5(CLBLM_L_X8Y155_SLICE_X10Y155_CQ),
.O5(CLBLM_R_X5Y155_SLICE_X6Y155_CO5),
.O6(CLBLM_R_X5Y155_SLICE_X6Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000040005)
  ) CLBLM_R_X5Y155_SLICE_X6Y155_BLUT (
.I0(CLBLM_R_X7Y155_SLICE_X9Y155_DO6),
.I1(CLBLM_R_X3Y154_SLICE_X3Y154_DO6),
.I2(CLBLM_R_X13Y155_SLICE_X19Y155_AO6),
.I3(CLBLM_R_X5Y156_SLICE_X6Y156_BO6),
.I4(CLBLL_L_X4Y156_SLICE_X4Y156_CO5),
.I5(CLBLM_R_X5Y155_SLICE_X6Y155_CO6),
.O5(CLBLM_R_X5Y155_SLICE_X6Y155_BO5),
.O6(CLBLM_R_X5Y155_SLICE_X6Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaee5044faee5044)
  ) CLBLM_R_X5Y155_SLICE_X6Y155_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y155_SLICE_X11Y155_BQ),
.I2(CLBLM_R_X5Y155_SLICE_X6Y155_AQ),
.I3(CLBLM_R_X7Y153_SLICE_X9Y153_CO6),
.I4(CLBLM_R_X3Y151_SLICE_X3Y151_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y155_SLICE_X6Y155_AO5),
.O6(CLBLM_R_X5Y155_SLICE_X6Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y155_SLICE_X7Y155_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y155_SLICE_X7Y155_AO6),
.Q(CLBLM_R_X5Y155_SLICE_X7Y155_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y155_SLICE_X7Y155_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y155_SLICE_X7Y155_BO6),
.Q(CLBLM_R_X5Y155_SLICE_X7Y155_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff0affce)
  ) CLBLM_R_X5Y155_SLICE_X7Y155_DLUT (
.I0(CLBLM_R_X5Y155_SLICE_X6Y155_AQ),
.I1(CLBLM_R_X5Y151_SLICE_X7Y151_DQ),
.I2(CLBLM_R_X3Y153_SLICE_X3Y153_AO6),
.I3(CLBLM_R_X5Y155_SLICE_X7Y155_CO6),
.I4(CLBLM_R_X3Y157_SLICE_X2Y157_AO5),
.I5(CLBLM_R_X7Y159_SLICE_X9Y159_DO6),
.O5(CLBLM_R_X5Y155_SLICE_X7Y155_DO5),
.O6(CLBLM_R_X5Y155_SLICE_X7Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010000000000)
  ) CLBLM_R_X5Y155_SLICE_X7Y155_CLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLL_L_X4Y157_SLICE_X4Y157_CO5),
.I3(CLBLM_L_X8Y155_SLICE_X11Y155_AQ),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(RIOB33_X105Y133_IOB_X1Y133_I),
.O5(CLBLM_R_X5Y155_SLICE_X7Y155_CO5),
.O6(CLBLM_R_X5Y155_SLICE_X7Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0afacaca0ac)
  ) CLBLM_R_X5Y155_SLICE_X7Y155_BLUT (
.I0(CLBLM_R_X5Y151_SLICE_X7Y151_CQ),
.I1(CLBLM_R_X5Y155_SLICE_X7Y155_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y150_SLICE_X12Y150_A5Q),
.I4(CLBLM_L_X12Y155_SLICE_X16Y155_CO6),
.I5(CLBLM_L_X8Y155_SLICE_X10Y155_B5Q),
.O5(CLBLM_R_X5Y155_SLICE_X7Y155_BO5),
.O6(CLBLM_R_X5Y155_SLICE_X7Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaccccaaaac0c0)
  ) CLBLM_R_X5Y155_SLICE_X7Y155_ALUT (
.I0(CLBLL_L_X4Y151_SLICE_X4Y151_DQ),
.I1(CLBLM_R_X7Y153_SLICE_X9Y153_CO6),
.I2(CLBLM_R_X5Y155_SLICE_X7Y155_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y156_SLICE_X10Y156_CQ),
.O5(CLBLM_R_X5Y155_SLICE_X7Y155_AO5),
.O6(CLBLM_R_X5Y155_SLICE_X7Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00c000c0a0e0a0e0)
  ) CLBLM_R_X5Y156_SLICE_X6Y156_DLUT (
.I0(CLBLM_L_X8Y155_SLICE_X10Y155_CQ),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(CLBLM_R_X3Y158_SLICE_X2Y158_AO6),
.I3(CLBLL_L_X2Y155_SLICE_X1Y155_CO6),
.I4(1'b1),
.I5(CLBLL_L_X2Y155_SLICE_X1Y155_CO5),
.O5(CLBLM_R_X5Y156_SLICE_X6Y156_DO5),
.O6(CLBLM_R_X5Y156_SLICE_X6Y156_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000c000c0a0e0a0e)
  ) CLBLM_R_X5Y156_SLICE_X6Y156_CLUT (
.I0(CLBLM_R_X7Y148_SLICE_X9Y148_AQ),
.I1(CLBLM_R_X5Y151_SLICE_X6Y151_AQ),
.I2(CLBLL_L_X4Y157_SLICE_X4Y157_CO5),
.I3(CLBLL_L_X2Y155_SLICE_X1Y155_CO6),
.I4(1'b1),
.I5(CLBLL_L_X2Y155_SLICE_X1Y155_CO5),
.O5(CLBLM_R_X5Y156_SLICE_X6Y156_CO5),
.O6(CLBLM_R_X5Y156_SLICE_X6Y156_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h44f444f4ffff44f4)
  ) CLBLM_R_X5Y156_SLICE_X6Y156_BLUT (
.I0(CLBLL_L_X4Y156_SLICE_X4Y156_CO6),
.I1(CLBLM_R_X5Y155_SLICE_X7Y155_BQ),
.I2(CLBLM_R_X5Y151_SLICE_X6Y151_AQ),
.I3(CLBLL_L_X4Y157_SLICE_X4Y157_BO6),
.I4(CLBLM_R_X7Y148_SLICE_X9Y148_AQ),
.I5(CLBLM_R_X3Y154_SLICE_X3Y154_AO6),
.O5(CLBLM_R_X5Y156_SLICE_X6Y156_BO5),
.O6(CLBLM_R_X5Y156_SLICE_X6Y156_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffafe)
  ) CLBLM_R_X5Y156_SLICE_X6Y156_ALUT (
.I0(CLBLM_R_X5Y156_SLICE_X6Y156_DO6),
.I1(CLBLM_R_X5Y155_SLICE_X7Y155_BQ),
.I2(CLBLL_L_X4Y156_SLICE_X5Y156_DO6),
.I3(CLBLL_L_X4Y156_SLICE_X4Y156_CO6),
.I4(CLBLL_L_X4Y155_SLICE_X5Y155_CO6),
.I5(CLBLM_R_X5Y156_SLICE_X6Y156_CO6),
.O5(CLBLM_R_X5Y156_SLICE_X6Y156_AO5),
.O6(CLBLM_R_X5Y156_SLICE_X6Y156_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y156_SLICE_X7Y156_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y156_SLICE_X7Y156_AO6),
.Q(CLBLM_R_X5Y156_SLICE_X7Y156_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffff0fffa)
  ) CLBLM_R_X5Y156_SLICE_X7Y156_DLUT (
.I0(CLBLM_R_X7Y156_SLICE_X9Y156_AQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y157_SLICE_X6Y157_BO6),
.I3(CLBLM_R_X5Y156_SLICE_X7Y156_CO6),
.I4(CLBLM_R_X3Y154_SLICE_X3Y154_AO6),
.I5(CLBLM_R_X5Y156_SLICE_X7Y156_BO6),
.O5(CLBLM_R_X5Y156_SLICE_X7Y156_DO5),
.O6(CLBLM_R_X5Y156_SLICE_X7Y156_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h50ff000050500000)
  ) CLBLM_R_X5Y156_SLICE_X7Y156_CLUT (
.I0(CLBLL_L_X2Y155_SLICE_X1Y155_CO6),
.I1(1'b1),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(CLBLM_R_X3Y156_SLICE_X3Y156_AO5),
.I4(CLBLM_R_X3Y158_SLICE_X2Y158_AO6),
.I5(CLBLM_L_X8Y154_SLICE_X10Y154_DQ),
.O5(CLBLM_R_X5Y156_SLICE_X7Y156_CO5),
.O6(CLBLM_R_X5Y156_SLICE_X7Y156_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000ca0000)
  ) CLBLM_R_X5Y156_SLICE_X7Y156_BLUT (
.I0(CLBLM_R_X7Y157_SLICE_X9Y157_BQ),
.I1(CLBLM_R_X5Y152_SLICE_X7Y152_BQ),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(CLBLL_L_X4Y157_SLICE_X4Y157_CO5),
.I4(RIOB33_X105Y131_IOB_X1Y132_I),
.I5(CLBLL_L_X4Y157_SLICE_X4Y157_AO5),
.O5(CLBLM_R_X5Y156_SLICE_X7Y156_BO5),
.O6(CLBLM_R_X5Y156_SLICE_X7Y156_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0aaccccf0aa)
  ) CLBLM_R_X5Y156_SLICE_X7Y156_ALUT (
.I0(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I1(CLBLM_L_X12Y158_SLICE_X16Y158_A5Q),
.I2(CLBLM_R_X5Y156_SLICE_X7Y156_AQ),
.I3(CLBLL_L_X4Y147_SLICE_X4Y147_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y156_SLICE_X7Y156_AO5),
.O6(CLBLM_R_X5Y156_SLICE_X7Y156_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y157_SLICE_X6Y157_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y157_SLICE_X6Y157_AO6),
.Q(CLBLM_R_X5Y157_SLICE_X6Y157_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcecececeffceffce)
  ) CLBLM_R_X5Y157_SLICE_X6Y157_DLUT (
.I0(CLBLL_L_X4Y156_SLICE_X4Y156_AQ),
.I1(CLBLM_R_X5Y158_SLICE_X7Y158_AO6),
.I2(CLBLL_L_X4Y156_SLICE_X4Y156_CO5),
.I3(CLBLM_R_X7Y158_SLICE_X8Y158_AQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y157_SLICE_X4Y157_BO5),
.O5(CLBLM_R_X5Y157_SLICE_X6Y157_DO5),
.O6(CLBLM_R_X5Y157_SLICE_X6Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000000e2e2)
  ) CLBLM_R_X5Y157_SLICE_X6Y157_CLUT (
.I0(CLBLM_R_X5Y152_SLICE_X7Y152_AQ),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(CLBLM_R_X7Y157_SLICE_X9Y157_CQ),
.I3(1'b1),
.I4(CLBLL_L_X4Y157_SLICE_X5Y157_AO5),
.I5(CLBLL_L_X4Y157_SLICE_X4Y157_CO5),
.O5(CLBLM_R_X5Y157_SLICE_X6Y157_CO5),
.O6(CLBLM_R_X5Y157_SLICE_X6Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000041014000)
  ) CLBLM_R_X5Y157_SLICE_X6Y157_BLUT (
.I0(CLBLL_L_X4Y157_SLICE_X5Y157_AO5),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y135_IOB_X1Y136_I),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_AQ),
.I4(CLBLM_R_X7Y158_SLICE_X9Y158_AQ),
.I5(CLBLM_R_X3Y158_SLICE_X2Y158_AO5),
.O5(CLBLM_R_X5Y157_SLICE_X6Y157_BO5),
.O6(CLBLM_R_X5Y157_SLICE_X6Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0ccccaaaa)
  ) CLBLM_R_X5Y157_SLICE_X6Y157_ALUT (
.I0(CLBLM_L_X12Y158_SLICE_X16Y158_A5Q),
.I1(CLBLM_R_X7Y157_SLICE_X8Y157_AQ),
.I2(CLBLM_R_X5Y157_SLICE_X6Y157_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y153_SLICE_X9Y153_CO6),
.O5(CLBLM_R_X5Y157_SLICE_X6Y157_AO5),
.O6(CLBLM_R_X5Y157_SLICE_X6Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y157_SLICE_X7Y157_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y157_SLICE_X7Y157_AO6),
.Q(CLBLM_R_X5Y157_SLICE_X7Y157_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y157_SLICE_X7Y157_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y157_SLICE_X7Y157_BO6),
.Q(CLBLM_R_X5Y157_SLICE_X7Y157_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y157_SLICE_X7Y157_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y157_SLICE_X7Y157_CO6),
.Q(CLBLM_R_X5Y157_SLICE_X7Y157_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y157_SLICE_X7Y157_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y157_SLICE_X7Y157_DO6),
.Q(CLBLM_R_X5Y157_SLICE_X7Y157_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00af05fa50)
  ) CLBLM_R_X5Y157_SLICE_X7Y157_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X5Y149_SLICE_X7Y149_DO6),
.I3(CLBLM_R_X5Y157_SLICE_X7Y157_BQ),
.I4(CLBLM_L_X8Y153_SLICE_X11Y153_DQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X5Y157_SLICE_X7Y157_DO5),
.O6(CLBLM_R_X5Y157_SLICE_X7Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffee440000ee44)
  ) CLBLM_R_X5Y157_SLICE_X7Y157_CLUT (
.I0(CLBLM_R_X5Y152_SLICE_X6Y152_CO5),
.I1(CLBLM_R_X5Y157_SLICE_X7Y157_CQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y156_SLICE_X9Y156_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X5Y154_SLICE_X7Y154_AQ),
.O5(CLBLM_R_X5Y157_SLICE_X7Y157_CO5),
.O6(CLBLM_R_X5Y157_SLICE_X7Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaee5044faee5044)
  ) CLBLM_R_X5Y157_SLICE_X7Y157_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X5Y157_SLICE_X7Y157_BQ),
.I2(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.I3(CLBLM_R_X5Y152_SLICE_X6Y152_CO5),
.I4(CLBLM_L_X8Y157_SLICE_X10Y157_AQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y157_SLICE_X7Y157_BO5),
.O6(CLBLM_R_X5Y157_SLICE_X7Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafff0aaaa0000)
  ) CLBLM_R_X5Y157_SLICE_X7Y157_ALUT (
.I0(CLBLM_R_X5Y157_SLICE_X7Y157_CQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y157_SLICE_X7Y157_AQ),
.I3(CLBLM_L_X10Y153_SLICE_X13Y153_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y153_SLICE_X9Y153_CO6),
.O5(CLBLM_R_X5Y157_SLICE_X7Y157_AO5),
.O6(CLBLM_R_X5Y157_SLICE_X7Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y158_SLICE_X6Y158_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y158_SLICE_X6Y158_AO6),
.Q(CLBLM_R_X5Y158_SLICE_X6Y158_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y158_SLICE_X6Y158_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X5Y158_SLICE_X6Y158_BO6),
.Q(CLBLM_R_X5Y158_SLICE_X6Y158_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y158_SLICE_X6Y158_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y158_SLICE_X6Y158_DO5),
.O6(CLBLM_R_X5Y158_SLICE_X6Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0010001022320010)
  ) CLBLM_R_X5Y158_SLICE_X6Y158_CLUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(CLBLM_R_X3Y158_SLICE_X2Y158_AO5),
.I2(CLBLM_R_X5Y158_SLICE_X6Y158_AQ),
.I3(CLBLL_L_X2Y155_SLICE_X1Y155_CO6),
.I4(CLBLM_R_X7Y153_SLICE_X8Y153_CQ),
.I5(CLBLM_R_X3Y156_SLICE_X3Y156_AO5),
.O5(CLBLM_R_X5Y158_SLICE_X6Y158_CO5),
.O6(CLBLM_R_X5Y158_SLICE_X6Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff0ccf000f0cc)
  ) CLBLM_R_X5Y158_SLICE_X6Y158_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y158_SLICE_X6Y158_BQ),
.I2(CLBLM_R_X5Y158_SLICE_X6Y158_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y152_SLICE_X6Y152_CO5),
.I5(CLBLM_L_X10Y150_SLICE_X12Y150_CQ),
.O5(CLBLM_R_X5Y158_SLICE_X6Y158_BO5),
.O6(CLBLM_R_X5Y158_SLICE_X6Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccf0ccaaccf0)
  ) CLBLM_R_X5Y158_SLICE_X6Y158_ALUT (
.I0(CLBLL_L_X4Y153_SLICE_X5Y153_AQ),
.I1(CLBLM_L_X8Y153_SLICE_X11Y153_AQ),
.I2(CLBLM_R_X5Y158_SLICE_X6Y158_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y152_SLICE_X6Y152_CO5),
.I5(1'b1),
.O5(CLBLM_R_X5Y158_SLICE_X6Y158_AO5),
.O6(CLBLM_R_X5Y158_SLICE_X6Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y158_SLICE_X7Y158_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y158_SLICE_X7Y158_DO5),
.O6(CLBLM_R_X5Y158_SLICE_X7Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y158_SLICE_X7Y158_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y158_SLICE_X7Y158_CO5),
.O6(CLBLM_R_X5Y158_SLICE_X7Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y158_SLICE_X7Y158_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y158_SLICE_X7Y158_BO5),
.O6(CLBLM_R_X5Y158_SLICE_X7Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000330022223322)
  ) CLBLM_R_X5Y158_SLICE_X7Y158_ALUT (
.I0(CLBLM_L_X8Y158_SLICE_X11Y158_BQ),
.I1(CLBLL_L_X4Y157_SLICE_X4Y157_CO5),
.I2(1'b1),
.I3(CLBLM_R_X5Y158_SLICE_X6Y158_BQ),
.I4(CLBLL_L_X2Y155_SLICE_X1Y155_CO5),
.I5(CLBLL_L_X2Y155_SLICE_X1Y155_CO6),
.O5(CLBLM_R_X5Y158_SLICE_X7Y158_AO5),
.O6(CLBLM_R_X5Y158_SLICE_X7Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y144_SLICE_X8Y144_AO6),
.Q(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y144_SLICE_X8Y144_DO5),
.O6(CLBLM_R_X7Y144_SLICE_X8Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y144_SLICE_X8Y144_CO5),
.O6(CLBLM_R_X7Y144_SLICE_X8Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa000000000000)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_BLUT (
.I0(CLBLM_R_X7Y145_SLICE_X8Y145_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X5Y146_SLICE_X6Y146_AQ),
.I5(CLBLM_R_X5Y146_SLICE_X6Y146_A5Q),
.O5(CLBLM_R_X7Y144_SLICE_X8Y144_BO5),
.O6(CLBLM_R_X7Y144_SLICE_X8Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888bb888888888)
  ) CLBLM_R_X7Y144_SLICE_X8Y144_ALUT (
.I0(CLBLM_R_X7Y157_SLICE_X8Y157_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.I3(CLBLM_R_X7Y144_SLICE_X8Y144_BO6),
.I4(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y144_SLICE_X8Y144_AO5),
.O6(CLBLM_R_X7Y144_SLICE_X8Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y144_SLICE_X9Y144_DO5),
.O6(CLBLM_R_X7Y144_SLICE_X9Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y144_SLICE_X9Y144_CO5),
.O6(CLBLM_R_X7Y144_SLICE_X9Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y144_SLICE_X9Y144_BO5),
.O6(CLBLM_R_X7Y144_SLICE_X9Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y144_SLICE_X9Y144_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y144_SLICE_X9Y144_AO5),
.O6(CLBLM_R_X7Y144_SLICE_X9Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y145_SLICE_X8Y145_AO6),
.Q(CLBLM_R_X7Y145_SLICE_X8Y145_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y145_SLICE_X8Y145_DO5),
.O6(CLBLM_R_X7Y145_SLICE_X8Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y145_SLICE_X8Y145_CO5),
.O6(CLBLM_R_X7Y145_SLICE_X8Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y145_SLICE_X8Y145_BO5),
.O6(CLBLM_R_X7Y145_SLICE_X8Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff12ff0000120000)
  ) CLBLM_R_X7Y145_SLICE_X8Y145_ALUT (
.I0(CLBLM_R_X5Y146_SLICE_X6Y146_A5Q),
.I1(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I2(CLBLM_R_X7Y145_SLICE_X8Y145_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X10Y145_SLICE_X12Y145_AQ),
.O5(CLBLM_R_X7Y145_SLICE_X8Y145_AO5),
.O6(CLBLM_R_X7Y145_SLICE_X8Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y145_SLICE_X9Y145_DO5),
.O6(CLBLM_R_X7Y145_SLICE_X9Y145_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y145_SLICE_X9Y145_CO5),
.O6(CLBLM_R_X7Y145_SLICE_X9Y145_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y145_SLICE_X9Y145_BO5),
.O6(CLBLM_R_X7Y145_SLICE_X9Y145_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y145_SLICE_X9Y145_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y145_SLICE_X9Y145_AO5),
.O6(CLBLM_R_X7Y145_SLICE_X9Y145_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y146_SLICE_X8Y146_AO6),
.Q(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff05ffffff05)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_DLUT (
.I0(CLBLM_R_X7Y148_SLICE_X9Y148_CO5),
.I1(1'b1),
.I2(CLBLM_R_X7Y146_SLICE_X9Y146_BO6),
.I3(CLBLM_R_X7Y147_SLICE_X8Y147_CO6),
.I4(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y146_SLICE_X8Y146_DO5),
.O6(CLBLM_R_X7Y146_SLICE_X8Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffcd)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_CLUT (
.I0(CLBLM_R_X7Y148_SLICE_X9Y148_CO5),
.I1(CLBLM_R_X7Y147_SLICE_X8Y147_DO6),
.I2(CLBLM_R_X7Y146_SLICE_X9Y146_BO6),
.I3(CLBLM_R_X5Y147_SLICE_X7Y147_C5Q),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_BO5),
.I5(CLBLL_L_X4Y146_SLICE_X5Y146_AQ),
.O5(CLBLM_R_X7Y146_SLICE_X8Y146_CO5),
.O6(CLBLM_R_X7Y146_SLICE_X8Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffeffffaaaaffff)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_BLUT (
.I0(CLBLM_R_X5Y150_SLICE_X7Y150_A5Q),
.I1(CLBLM_R_X5Y147_SLICE_X7Y147_C5Q),
.I2(CLBLM_R_X7Y147_SLICE_X8Y147_DO6),
.I3(CLBLL_L_X4Y146_SLICE_X5Y146_AQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y146_SLICE_X8Y146_BO5),
.O6(CLBLM_R_X7Y146_SLICE_X8Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaafeba55005410)
  ) CLBLM_R_X7Y146_SLICE_X8Y146_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I3(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I4(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I5(CLBLM_R_X5Y146_SLICE_X6Y146_A5Q),
.O5(CLBLM_R_X7Y146_SLICE_X8Y146_AO5),
.O6(CLBLM_R_X7Y146_SLICE_X8Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y146_SLICE_X9Y146_AO6),
.Q(CLBLM_R_X7Y146_SLICE_X9Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffff0)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I3(CLBLM_R_X7Y146_SLICE_X9Y146_CO6),
.I4(CLBLM_R_X5Y150_SLICE_X7Y150_A5Q),
.I5(CLBLM_R_X7Y147_SLICE_X9Y147_A5Q),
.O5(CLBLM_R_X7Y146_SLICE_X9Y146_DO5),
.O6(CLBLM_R_X7Y146_SLICE_X9Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0fffffff5ffff)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_CLUT (
.I0(CLBLM_R_X7Y148_SLICE_X9Y148_CO5),
.I1(1'b1),
.I2(CLBLM_L_X8Y153_SLICE_X11Y153_C5Q),
.I3(CLBLM_R_X7Y147_SLICE_X8Y147_BO5),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y146_SLICE_X9Y146_BO6),
.O5(CLBLM_R_X7Y146_SLICE_X9Y146_CO5),
.O6(CLBLM_R_X7Y146_SLICE_X9Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_BLUT (
.I0(CLBLM_R_X3Y156_SLICE_X2Y156_DO6),
.I1(CLBLM_R_X3Y155_SLICE_X2Y155_BO6),
.I2(CLBLL_L_X4Y154_SLICE_X5Y154_CO6),
.I3(CLBLL_L_X4Y153_SLICE_X4Y153_BO6),
.I4(CLBLL_L_X4Y154_SLICE_X5Y154_BO6),
.I5(CLBLM_R_X5Y155_SLICE_X6Y155_DO6),
.O5(CLBLM_R_X7Y146_SLICE_X9Y146_BO5),
.O6(CLBLM_R_X7Y146_SLICE_X9Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa33aa30aa33aa30)
  ) CLBLM_R_X7Y146_SLICE_X9Y146_ALUT (
.I0(CLBLM_R_X5Y150_SLICE_X7Y150_A5Q),
.I1(CLBLM_R_X7Y146_SLICE_X8Y146_DO6),
.I2(CLBLM_R_X7Y146_SLICE_X9Y146_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y146_SLICE_X12Y146_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y146_SLICE_X9Y146_AO5),
.O6(CLBLM_R_X7Y146_SLICE_X9Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X8Y147_AO6),
.Q(CLBLM_R_X7Y147_SLICE_X8Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_DLUT (
.I0(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.I1(CLBLM_R_X7Y147_SLICE_X9Y147_A5Q),
.I2(CLBLM_R_X5Y149_SLICE_X6Y149_AQ),
.I3(CLBLM_L_X8Y153_SLICE_X11Y153_C5Q),
.I4(CLBLM_R_X5Y148_SLICE_X7Y148_A5Q),
.I5(CLBLM_R_X5Y151_SLICE_X6Y151_C5Q),
.O5(CLBLM_R_X7Y147_SLICE_X8Y147_DO5),
.O6(CLBLM_R_X7Y147_SLICE_X8Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffeffff)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_CLUT (
.I0(CLBLM_R_X7Y147_SLICE_X9Y147_A5Q),
.I1(CLBLM_R_X5Y149_SLICE_X6Y149_AQ),
.I2(CLBLM_L_X8Y153_SLICE_X11Y153_C5Q),
.I3(CLBLM_R_X5Y150_SLICE_X7Y150_A5Q),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X7Y147_SLICE_X8Y147_BO6),
.O5(CLBLM_R_X7Y147_SLICE_X8Y147_CO5),
.O6(CLBLM_R_X7Y147_SLICE_X8Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffcfffffffe)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_BLUT (
.I0(CLBLM_R_X5Y149_SLICE_X6Y149_AQ),
.I1(CLBLM_R_X5Y148_SLICE_X7Y148_A5Q),
.I2(CLBLM_R_X5Y147_SLICE_X7Y147_C5Q),
.I3(CLBLM_R_X5Y151_SLICE_X6Y151_C5Q),
.I4(CLBLL_L_X4Y146_SLICE_X5Y146_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y147_SLICE_X8Y147_BO5),
.O6(CLBLM_R_X7Y147_SLICE_X8Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff000f0ffaa00aa)
  ) CLBLM_R_X7Y147_SLICE_X8Y147_ALUT (
.I0(CLBLM_R_X5Y149_SLICE_X6Y149_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y147_SLICE_X8Y147_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y145_SLICE_X8Y145_AQ),
.I5(CLBLL_L_X4Y147_SLICE_X4Y147_BO6),
.O5(CLBLM_R_X7Y147_SLICE_X8Y147_AO5),
.O6(CLBLM_R_X7Y147_SLICE_X8Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X9Y147_AO5),
.Q(CLBLM_R_X7Y147_SLICE_X9Y147_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X9Y147_AO6),
.Q(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X9Y147_BO6),
.Q(CLBLM_R_X7Y147_SLICE_X9Y147_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y147_SLICE_X9Y147_CO6),
.Q(CLBLM_R_X7Y147_SLICE_X9Y147_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00002000ffffdf5f)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_DLUT (
.I0(CLBLM_L_X8Y147_SLICE_X10Y147_BQ),
.I1(CLBLM_R_X7Y147_SLICE_X9Y147_CQ),
.I2(CLBLM_L_X8Y147_SLICE_X10Y147_AQ),
.I3(CLBLM_R_X7Y147_SLICE_X9Y147_BQ),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y147_SLICE_X9Y147_DO5),
.O6(CLBLM_R_X7Y147_SLICE_X9Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00f000c0)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_CLUT (
.I0(CLBLM_R_X7Y151_SLICE_X9Y151_AQ),
.I1(CLBLM_R_X7Y147_SLICE_X9Y147_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y154_SLICE_X13Y154_CQ),
.I4(CLBLM_R_X7Y147_SLICE_X9Y147_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y147_SLICE_X9Y147_CO5),
.O6(CLBLM_R_X7Y147_SLICE_X9Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f8f20802)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y147_SLICE_X9Y147_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y147_SLICE_X9Y147_DO5),
.I4(CLBLM_R_X7Y147_SLICE_X8Y147_AQ),
.I5(CLBLM_L_X10Y154_SLICE_X13Y154_CQ),
.O5(CLBLM_R_X7Y147_SLICE_X9Y147_BO5),
.O6(CLBLM_R_X7Y147_SLICE_X9Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdd88dd88f5f5a0a0)
  ) CLBLM_R_X7Y147_SLICE_X9Y147_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X3Y151_SLICE_X2Y151_AQ),
.I2(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I3(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I4(CLBLM_L_X10Y149_SLICE_X12Y149_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y147_SLICE_X9Y147_AO5),
.O6(CLBLM_R_X7Y147_SLICE_X9Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X8Y148_DO6),
.Q(CLBLM_R_X7Y148_SLICE_X8Y148_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X8Y148_AO6),
.Q(CLBLM_R_X7Y148_SLICE_X8Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X8Y148_BO6),
.Q(CLBLM_R_X7Y148_SLICE_X8Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X8Y148_CO6),
.Q(CLBLM_R_X7Y148_SLICE_X8Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f077ddcc00cc00)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_DLUT (
.I0(CLBLM_L_X10Y149_SLICE_X12Y149_DO5),
.I1(CLBLM_L_X10Y149_SLICE_X12Y149_BQ),
.I2(CLBLM_L_X12Y151_SLICE_X16Y151_AQ),
.I3(CLBLM_R_X7Y148_SLICE_X8Y148_A5Q),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y148_SLICE_X8Y148_DO5),
.O6(CLBLM_R_X7Y148_SLICE_X8Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf2f80208f8f80808)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_CLUT (
.I0(CLBLM_L_X10Y149_SLICE_X12Y149_DO5),
.I1(CLBLM_R_X7Y148_SLICE_X8Y148_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y148_SLICE_X5Y148_DQ),
.I4(CLBLM_R_X7Y151_SLICE_X9Y151_CQ),
.I5(CLBLM_R_X7Y148_SLICE_X8Y148_DO5),
.O5(CLBLM_R_X7Y148_SLICE_X8Y148_CO5),
.O6(CLBLM_R_X7Y148_SLICE_X8Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf2fa020af2f80208)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_BLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_R_X7Y148_SLICE_X8Y148_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y159_SLICE_X8Y159_BO6),
.I4(CLBLM_R_X7Y146_SLICE_X9Y146_AQ),
.I5(CLBLM_R_X7Y158_SLICE_X8Y158_CO5),
.O5(CLBLM_R_X7Y148_SLICE_X8Y148_BO5),
.O6(CLBLM_R_X7Y148_SLICE_X8Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff440044ff500050)
  ) CLBLM_R_X7Y148_SLICE_X8Y148_ALUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_R_X7Y148_SLICE_X8Y148_BQ),
.I2(CLBLM_R_X7Y148_SLICE_X8Y148_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y144_SLICE_X6Y144_AQ),
.I5(CLBLM_L_X10Y159_SLICE_X12Y159_AO6),
.O5(CLBLM_R_X7Y148_SLICE_X8Y148_AO5),
.O6(CLBLM_R_X7Y148_SLICE_X8Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X9Y148_AO6),
.Q(CLBLM_R_X7Y148_SLICE_X9Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y148_SLICE_X9Y148_BO6),
.Q(CLBLM_R_X7Y148_SLICE_X9Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff1155ffff33ff)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_DLUT (
.I0(CLBLL_L_X4Y154_SLICE_X5Y154_CO6),
.I1(CLBLM_R_X5Y155_SLICE_X6Y155_DO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y155_SLICE_X2Y155_BO6),
.I4(CLBLM_L_X10Y150_SLICE_X13Y150_BQ),
.I5(CLBLL_L_X4Y153_SLICE_X4Y153_BO6),
.O5(CLBLM_R_X7Y148_SLICE_X9Y148_DO5),
.O6(CLBLM_R_X7Y148_SLICE_X9Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000dc50ff55ff55)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_CLUT (
.I0(CLBLL_L_X4Y153_SLICE_X4Y153_AO6),
.I1(CLBLM_R_X3Y156_SLICE_X2Y156_DO6),
.I2(CLBLL_L_X4Y154_SLICE_X5Y154_BO6),
.I3(CLBLL_L_X4Y154_SLICE_X4Y154_BO6),
.I4(CLBLM_R_X7Y148_SLICE_X9Y148_DO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y148_SLICE_X9Y148_CO5),
.O6(CLBLM_R_X7Y148_SLICE_X9Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffee5544faea5040)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y148_SLICE_X9Y148_BQ),
.I2(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I3(CLBLM_L_X8Y146_SLICE_X10Y146_AQ),
.I4(CLBLM_R_X5Y147_SLICE_X7Y147_C5Q),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X7Y148_SLICE_X9Y148_BO5),
.O6(CLBLM_R_X7Y148_SLICE_X9Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heeeaccc0eeeaccc0)
  ) CLBLM_R_X7Y148_SLICE_X9Y148_ALUT (
.I0(CLBLM_L_X8Y148_SLICE_X10Y148_CQ),
.I1(CLBLM_R_X5Y152_SLICE_X6Y152_CO6),
.I2(CLBLM_R_X7Y148_SLICE_X9Y148_AQ),
.I3(CLBLM_R_X7Y151_SLICE_X8Y151_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y148_SLICE_X9Y148_AO5),
.O6(CLBLM_R_X7Y148_SLICE_X9Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y149_SLICE_X8Y149_AO6),
.Q(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y149_SLICE_X8Y149_BO6),
.Q(CLBLM_R_X7Y149_SLICE_X8Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y149_SLICE_X8Y149_CO6),
.Q(CLBLM_R_X7Y149_SLICE_X8Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h223332330000ffaa)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_DLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I1(CLBLM_R_X5Y149_SLICE_X7Y149_A5Q),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.I4(CLBLL_L_X4Y154_SLICE_X5Y154_BO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y149_SLICE_X8Y149_DO5),
.O6(CLBLM_R_X7Y149_SLICE_X8Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc0000ff00)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y149_SLICE_X7Y149_A5Q),
.I2(1'b1),
.I3(CLBLM_R_X5Y151_SLICE_X6Y151_CQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y149_SLICE_X8Y149_CO5),
.O6(CLBLM_R_X7Y149_SLICE_X8Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55fe54aa00ae04)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y149_SLICE_X8Y149_BQ),
.I2(RIOB33_X105Y117_IOB_X1Y118_I),
.I3(CLBLM_R_X5Y150_SLICE_X7Y150_CQ),
.I4(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I5(CLBLM_L_X8Y149_SLICE_X11Y149_CQ),
.O5(CLBLM_R_X7Y149_SLICE_X8Y149_BO5),
.O6(CLBLM_R_X7Y149_SLICE_X8Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffaffeaaafaaaea)
  ) CLBLM_R_X7Y149_SLICE_X8Y149_ALUT (
.I0(CLBLM_R_X7Y150_SLICE_X9Y150_CO6),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I5(CLBLL_L_X4Y149_SLICE_X5Y149_A5Q),
.O5(CLBLM_R_X7Y149_SLICE_X8Y149_AO5),
.O6(CLBLM_R_X7Y149_SLICE_X8Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_C5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y149_SLICE_X9Y149_CO5),
.Q(CLBLM_R_X7Y149_SLICE_X9Y149_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y149_SLICE_X9Y149_AO6),
.Q(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y149_SLICE_X9Y149_BO6),
.Q(CLBLM_R_X7Y149_SLICE_X9Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X7Y149_SLICE_X9Y149_CO6),
.Q(CLBLM_R_X7Y149_SLICE_X9Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00005f5f0000ffcc)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_DLUT (
.I0(CLBLM_R_X3Y156_SLICE_X2Y156_DO6),
.I1(CLBLM_L_X8Y148_SLICE_X10Y148_CQ),
.I2(CLBLM_L_X8Y155_SLICE_X10Y155_B5Q),
.I3(CLBLM_R_X5Y149_SLICE_X7Y149_A5Q),
.I4(CLBLM_L_X10Y150_SLICE_X13Y150_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y149_SLICE_X9Y149_DO5),
.O6(CLBLM_R_X7Y149_SLICE_X9Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f000ffcccc5500)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_CLUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_C5Q),
.I1(CLBLM_R_X11Y149_SLICE_X15Y149_A5Q),
.I2(CLBLM_R_X7Y156_SLICE_X9Y156_BQ),
.I3(RIOB33_X105Y119_IOB_X1Y119_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y149_SLICE_X9Y149_CO5),
.O6(CLBLM_R_X7Y149_SLICE_X9Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafffaeee05550444)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y149_SLICE_X9Y149_BQ),
.I2(CLBLL_L_X4Y151_SLICE_X4Y151_BQ),
.I3(CLBLM_L_X10Y151_SLICE_X12Y151_CQ),
.I4(CLBLM_L_X8Y149_SLICE_X10Y149_AQ),
.I5(CLBLM_R_X7Y149_SLICE_X9Y149_C5Q),
.O5(CLBLM_R_X7Y149_SLICE_X9Y149_BO5),
.O6(CLBLM_R_X7Y149_SLICE_X9Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccd0001cccc0000)
  ) CLBLM_R_X7Y149_SLICE_X9Y149_ALUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X5Y152_SLICE_X7Y152_AQ),
.I5(RIOB33_X105Y119_IOB_X1Y119_I),
.O5(CLBLM_R_X7Y149_SLICE_X9Y149_AO5),
.O6(CLBLM_R_X7Y149_SLICE_X9Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y150_SLICE_X8Y150_AO6),
.Q(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y150_SLICE_X8Y150_BO6),
.Q(CLBLM_R_X7Y150_SLICE_X8Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000030000)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y150_SLICE_X5Y150_DQ),
.I2(CLBLM_R_X7Y152_SLICE_X9Y152_DO6),
.I3(CLBLM_R_X7Y152_SLICE_X8Y152_A5Q),
.I4(CLBLM_R_X5Y150_SLICE_X7Y150_DO6),
.I5(CLBLM_R_X7Y151_SLICE_X9Y151_DO6),
.O5(CLBLM_R_X7Y150_SLICE_X8Y150_DO5),
.O6(CLBLM_R_X7Y150_SLICE_X8Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff00000eeee0000)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_CLUT (
.I0(CLBLM_L_X8Y150_SLICE_X11Y150_BQ),
.I1(CLBLM_R_X5Y152_SLICE_X6Y152_BQ),
.I2(CLBLL_L_X4Y150_SLICE_X4Y150_BQ),
.I3(CLBLM_L_X10Y149_SLICE_X12Y149_C5Q),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y150_SLICE_X8Y150_CO5),
.O6(CLBLM_R_X7Y150_SLICE_X8Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc05cc50cc05cc50)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y150_SLICE_X13Y150_BQ),
.I2(CLBLM_R_X7Y156_SLICE_X9Y156_BQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y150_SLICE_X8Y150_CO5),
.I5(1'b1),
.O5(CLBLM_R_X7Y150_SLICE_X8Y150_BO5),
.O6(CLBLM_R_X7Y150_SLICE_X8Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccfaccaaccfa)
  ) CLBLM_R_X7Y150_SLICE_X8Y150_ALUT (
.I0(CLBLM_R_X7Y150_SLICE_X8Y150_DO6),
.I1(CLBLM_R_X7Y155_SLICE_X9Y155_AQ),
.I2(CLBLM_R_X7Y150_SLICE_X8Y150_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y150_SLICE_X8Y150_AO5),
.O6(CLBLM_R_X7Y150_SLICE_X8Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffbfffffffff)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_DLUT (
.I0(CLBLM_R_X5Y147_SLICE_X7Y147_C5Q),
.I1(CLBLM_R_X5Y146_SLICE_X6Y146_A5Q),
.I2(RIOB33_X105Y119_IOB_X1Y119_I),
.I3(CLBLM_R_X7Y152_SLICE_X9Y152_BQ),
.I4(CLBLM_L_X10Y156_SLICE_X13Y156_AO6),
.I5(CLBLM_R_X13Y150_SLICE_X18Y150_DO5),
.O5(CLBLM_R_X7Y150_SLICE_X9Y150_DO5),
.O6(CLBLM_R_X7Y150_SLICE_X9Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cccc0800)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_CLUT (
.I0(CLBLM_R_X7Y152_SLICE_X9Y152_CO5),
.I1(CLBLM_R_X7Y154_SLICE_X8Y154_AO5),
.I2(CLBLL_L_X4Y153_SLICE_X4Y153_AO6),
.I3(CLBLM_R_X7Y150_SLICE_X9Y150_AO5),
.I4(CLBLM_L_X10Y152_SLICE_X12Y152_CO5),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y150_SLICE_X9Y150_CO5),
.O6(CLBLM_R_X7Y150_SLICE_X9Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5544555554445555)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_BLUT (
.I0(CLBLM_L_X10Y152_SLICE_X12Y152_CO5),
.I1(CLBLM_R_X3Y156_SLICE_X2Y156_DO6),
.I2(CLBLM_L_X8Y151_SLICE_X10Y151_AQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(CLBLM_R_X7Y152_SLICE_X9Y152_CO5),
.I5(CLBLM_R_X11Y149_SLICE_X15Y149_A5Q),
.O5(CLBLM_R_X7Y150_SLICE_X9Y150_BO5),
.O6(CLBLM_R_X7Y150_SLICE_X9Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaff00c0c0ffff)
  ) CLBLM_R_X7Y150_SLICE_X9Y150_ALUT (
.I0(CLBLM_R_X11Y151_SLICE_X15Y151_AQ),
.I1(CLBLM_R_X7Y151_SLICE_X9Y151_AQ),
.I2(CLBLM_R_X7Y151_SLICE_X8Y151_DQ),
.I3(CLBLM_L_X10Y151_SLICE_X13Y151_AQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y150_SLICE_X9Y150_AO5),
.O6(CLBLM_R_X7Y150_SLICE_X9Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X8Y151_AO6),
.Q(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X8Y151_BO6),
.Q(CLBLM_R_X7Y151_SLICE_X8Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X8Y151_CO6),
.Q(CLBLM_R_X7Y151_SLICE_X8Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X8Y151_DO6),
.Q(CLBLM_R_X7Y151_SLICE_X8Y151_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaac0c0c0c0)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_DLUT (
.I0(CLBLM_R_X7Y157_SLICE_X8Y157_BQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X7Y151_SLICE_X9Y151_C5Q),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y151_SLICE_X8Y151_DO5),
.O6(CLBLM_R_X7Y151_SLICE_X8Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00c000c0)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_CLUT (
.I0(CLBLM_R_X7Y150_SLICE_X8Y150_BQ),
.I1(CLBLM_R_X7Y151_SLICE_X8Y151_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y151_SLICE_X9Y151_CQ),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y151_SLICE_X8Y151_CO5),
.O6(CLBLM_R_X7Y151_SLICE_X8Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000cccc0ff0)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y149_SLICE_X8Y149_BQ),
.I2(CLBLM_R_X7Y151_SLICE_X8Y151_AQ),
.I3(CLBLM_L_X8Y153_SLICE_X10Y153_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y151_SLICE_X8Y151_BO5),
.O6(CLBLM_R_X7Y151_SLICE_X8Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff11ff2200110022)
  ) CLBLM_R_X7Y151_SLICE_X8Y151_ALUT (
.I0(CLBLM_L_X10Y151_SLICE_X13Y151_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X8Y151_SLICE_X11Y151_AQ),
.I5(CLBLM_R_X7Y148_SLICE_X8Y148_CQ),
.O5(CLBLM_R_X7Y151_SLICE_X8Y151_AO5),
.O6(CLBLM_R_X7Y151_SLICE_X8Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X9Y151_CO5),
.Q(CLBLM_R_X7Y151_SLICE_X9Y151_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X9Y151_AO6),
.Q(CLBLM_R_X7Y151_SLICE_X9Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X9Y151_BO6),
.Q(CLBLM_R_X7Y151_SLICE_X9Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y151_SLICE_X9Y151_CO6),
.Q(CLBLM_R_X7Y151_SLICE_X9Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff3fffffff)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y150_SLICE_X4Y150_CQ),
.I2(CLBLM_R_X7Y151_SLICE_X9Y151_BQ),
.I3(CLBLM_R_X7Y154_SLICE_X9Y154_CQ),
.I4(CLBLM_R_X7Y152_SLICE_X9Y152_BQ),
.I5(CLBLM_R_X7Y151_SLICE_X8Y151_BQ),
.O5(CLBLM_R_X7Y151_SLICE_X9Y151_DO5),
.O6(CLBLM_R_X7Y151_SLICE_X9Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0aaaacccc00f0)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_CLUT (
.I0(CLBLM_R_X7Y155_SLICE_X9Y155_AQ),
.I1(CLBLM_R_X5Y151_SLICE_X6Y151_BQ),
.I2(CLBLM_R_X11Y151_SLICE_X15Y151_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y151_SLICE_X9Y151_CO5),
.O6(CLBLM_R_X7Y151_SLICE_X9Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc0000ddee1122)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_BLUT (
.I0(CLBLM_L_X8Y151_SLICE_X10Y151_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_L_X8Y151_SLICE_X11Y151_CO6),
.I4(CLBLM_L_X10Y152_SLICE_X12Y152_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y151_SLICE_X9Y151_BO5),
.O6(CLBLM_R_X7Y151_SLICE_X9Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccfedc33003210)
  ) CLBLM_R_X7Y151_SLICE_X9Y151_ALUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y151_SLICE_X9Y151_AQ),
.I3(CLBLM_L_X8Y153_SLICE_X10Y153_BO6),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_L_X8Y152_SLICE_X10Y152_CQ),
.O5(CLBLM_R_X7Y151_SLICE_X9Y151_AO5),
.O6(CLBLM_R_X7Y151_SLICE_X9Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y152_SLICE_X8Y152_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y152_SLICE_X8Y152_BO6),
.Q(CLBLM_R_X7Y152_SLICE_X8Y152_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y152_SLICE_X8Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y152_SLICE_X8Y152_AO6),
.Q(CLBLM_R_X7Y152_SLICE_X8Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffeffff)
  ) CLBLM_R_X7Y152_SLICE_X8Y152_DLUT (
.I0(CLBLM_R_X5Y150_SLICE_X7Y150_AQ),
.I1(CLBLM_R_X7Y157_SLICE_X9Y157_DQ),
.I2(CLBLM_L_X10Y150_SLICE_X13Y150_BQ),
.I3(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X5Y151_SLICE_X7Y151_CQ),
.O5(CLBLM_R_X7Y152_SLICE_X8Y152_DO5),
.O6(CLBLM_R_X7Y152_SLICE_X8Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffefffffffcf)
  ) CLBLM_R_X7Y152_SLICE_X8Y152_CLUT (
.I0(CLBLM_R_X7Y148_SLICE_X8Y148_AQ),
.I1(CLBLM_R_X7Y150_SLICE_X9Y150_DO6),
.I2(CLBLM_L_X8Y158_SLICE_X10Y158_AQ),
.I3(CLBLM_L_X8Y148_SLICE_X10Y148_DO6),
.I4(CLBLM_R_X7Y152_SLICE_X8Y152_DO6),
.I5(CLBLM_R_X7Y148_SLICE_X8Y148_BQ),
.O5(CLBLM_R_X7Y152_SLICE_X8Y152_CO5),
.O6(CLBLM_R_X7Y152_SLICE_X8Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0aca0ac0000ff00)
  ) CLBLM_R_X7Y152_SLICE_X8Y152_BLUT (
.I0(CLBLM_L_X8Y157_SLICE_X10Y157_DQ),
.I1(CLBLM_L_X8Y157_SLICE_X11Y157_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X7Y147_SLICE_X9Y147_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y152_SLICE_X8Y152_BO5),
.O6(CLBLM_R_X7Y152_SLICE_X8Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccff5accccff5a)
  ) CLBLM_R_X7Y152_SLICE_X8Y152_ALUT (
.I0(CLBLM_R_X7Y155_SLICE_X8Y155_DO6),
.I1(CLBLM_R_X7Y151_SLICE_X8Y151_BQ),
.I2(CLBLM_R_X7Y152_SLICE_X8Y152_AQ),
.I3(CLBLM_R_X7Y158_SLICE_X8Y158_CO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y152_SLICE_X8Y152_AO5),
.O6(CLBLM_R_X7Y152_SLICE_X8Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y152_SLICE_X9Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y152_SLICE_X9Y152_AO6),
.Q(CLBLM_R_X7Y152_SLICE_X9Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y152_SLICE_X9Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y152_SLICE_X9Y152_BO6),
.Q(CLBLM_R_X7Y152_SLICE_X9Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffbfffffffff)
  ) CLBLM_R_X7Y152_SLICE_X9Y152_DLUT (
.I0(CLBLM_R_X5Y154_SLICE_X6Y154_AQ),
.I1(CLBLM_R_X7Y153_SLICE_X9Y153_CO5),
.I2(CLBLM_L_X10Y157_SLICE_X12Y157_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X8Y151_SLICE_X11Y151_AQ),
.I5(CLBLM_L_X8Y157_SLICE_X11Y157_BQ),
.O5(CLBLM_R_X7Y152_SLICE_X9Y152_DO5),
.O6(CLBLM_R_X7Y152_SLICE_X9Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaaeae50505050)
  ) CLBLM_R_X7Y152_SLICE_X9Y152_CLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I1(CLBLM_R_X3Y155_SLICE_X2Y155_BO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X7Y150_SLICE_X8Y150_CO6),
.I4(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y152_SLICE_X9Y152_CO5),
.O6(CLBLM_R_X7Y152_SLICE_X9Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f10101f2f20202)
  ) CLBLM_R_X7Y152_SLICE_X9Y152_BLUT (
.I0(CLBLM_L_X8Y152_SLICE_X10Y152_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X13Y154_SLICE_X19Y154_AQ),
.I5(CLBLM_R_X7Y154_SLICE_X9Y154_CQ),
.O5(CLBLM_R_X7Y152_SLICE_X9Y152_BO5),
.O6(CLBLM_R_X7Y152_SLICE_X9Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffa8a8a8a8a8a8)
  ) CLBLM_R_X7Y152_SLICE_X9Y152_ALUT (
.I0(CLBLM_R_X5Y152_SLICE_X6Y152_CO6),
.I1(CLBLM_R_X7Y152_SLICE_X9Y152_BQ),
.I2(CLBLM_R_X7Y152_SLICE_X9Y152_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y152_SLICE_X16Y152_BQ),
.O5(CLBLM_R_X7Y152_SLICE_X9Y152_AO5),
.O6(CLBLM_R_X7Y152_SLICE_X9Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y153_SLICE_X8Y153_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y153_SLICE_X8Y153_AO5),
.Q(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y153_SLICE_X8Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y153_SLICE_X8Y153_AO6),
.Q(CLBLM_R_X7Y153_SLICE_X8Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y153_SLICE_X8Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y153_SLICE_X8Y153_BO6),
.Q(CLBLM_R_X7Y153_SLICE_X8Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y153_SLICE_X8Y153_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y153_SLICE_X8Y153_CO6),
.Q(CLBLM_R_X7Y153_SLICE_X8Y153_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffeffffffffffff)
  ) CLBLM_R_X7Y153_SLICE_X8Y153_DLUT (
.I0(CLBLM_R_X3Y151_SLICE_X2Y151_CO5),
.I1(CLBLM_R_X7Y152_SLICE_X8Y152_CO6),
.I2(CLBLM_R_X13Y156_SLICE_X18Y156_CO6),
.I3(CLBLM_R_X7Y155_SLICE_X8Y155_BO6),
.I4(CLBLM_L_X8Y155_SLICE_X11Y155_DO6),
.I5(CLBLM_R_X7Y153_SLICE_X9Y153_BQ),
.O5(CLBLM_R_X7Y153_SLICE_X8Y153_DO5),
.O6(CLBLM_R_X7Y153_SLICE_X8Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0aaaaccaa)
  ) CLBLM_R_X7Y153_SLICE_X8Y153_CLUT (
.I0(CLBLM_L_X10Y148_SLICE_X13Y148_AQ),
.I1(CLBLM_R_X7Y153_SLICE_X8Y153_CQ),
.I2(CLBLM_R_X7Y155_SLICE_X9Y155_A5Q),
.I3(CLBLM_L_X10Y150_SLICE_X12Y150_A5Q),
.I4(CLBLM_L_X12Y155_SLICE_X16Y155_CO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y153_SLICE_X8Y153_CO5),
.O6(CLBLM_R_X7Y153_SLICE_X8Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0afa0afa0)
  ) CLBLM_R_X7Y153_SLICE_X8Y153_BLUT (
.I0(CLBLM_R_X7Y156_SLICE_X8Y156_CQ),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y151_SLICE_X13Y151_BQ),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X7Y153_SLICE_X8Y153_BO5),
.O6(CLBLM_R_X7Y153_SLICE_X8Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa0afa0afcfc0c0c)
  ) CLBLM_R_X7Y153_SLICE_X8Y153_ALUT (
.I0(CLBLM_L_X8Y157_SLICE_X10Y157_AQ),
.I1(CLBLL_L_X4Y148_SLICE_X5Y148_DQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y158_SLICE_X10Y158_AQ),
.I4(CLBLM_L_X12Y150_SLICE_X16Y150_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y153_SLICE_X8Y153_AO5),
.O6(CLBLM_R_X7Y153_SLICE_X8Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y153_SLICE_X9Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y153_SLICE_X9Y153_AO6),
.Q(CLBLM_R_X7Y153_SLICE_X9Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y153_SLICE_X9Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y153_SLICE_X9Y153_BO6),
.Q(CLBLM_R_X7Y153_SLICE_X9Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5fff5fffffffffff)
  ) CLBLM_R_X7Y153_SLICE_X9Y153_DLUT (
.I0(CLBLL_L_X4Y153_SLICE_X5Y153_AQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y150_SLICE_X6Y150_AQ),
.I3(CLBLM_L_X10Y150_SLICE_X13Y150_CQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y153_SLICE_X12Y153_BQ),
.O5(CLBLM_R_X7Y153_SLICE_X9Y153_DO5),
.O6(CLBLM_R_X7Y153_SLICE_X9Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc8c8c50505050)
  ) CLBLM_R_X7Y153_SLICE_X9Y153_CLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X12Y149_SLICE_X16Y149_CQ),
.I3(1'b1),
.I4(CLBLM_R_X13Y150_SLICE_X18Y150_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y153_SLICE_X9Y153_CO5),
.O6(CLBLM_R_X7Y153_SLICE_X9Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000fffc0f0c)
  ) CLBLM_R_X7Y153_SLICE_X9Y153_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y153_SLICE_X9Y153_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y150_SLICE_X7Y150_A5Q),
.I4(CLBLM_L_X10Y158_SLICE_X13Y158_AQ),
.I5(CLBLL_L_X4Y147_SLICE_X4Y147_BO6),
.O5(CLBLM_R_X7Y153_SLICE_X9Y153_BO5),
.O6(CLBLM_R_X7Y153_SLICE_X9Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffa0f00000a0f0)
  ) CLBLM_R_X7Y153_SLICE_X9Y153_ALUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I1(1'b1),
.I2(CLBLM_R_X7Y153_SLICE_X9Y153_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y156_SLICE_X4Y156_AQ),
.O5(CLBLM_R_X7Y153_SLICE_X9Y153_AO5),
.O6(CLBLM_R_X7Y153_SLICE_X9Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y154_SLICE_X8Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y154_SLICE_X8Y154_AO6),
.Q(CLBLM_R_X7Y154_SLICE_X8Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y154_SLICE_X8Y154_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y154_SLICE_X8Y154_BO6),
.Q(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y154_SLICE_X8Y154_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y154_SLICE_X8Y154_CO6),
.Q(CLBLM_R_X7Y154_SLICE_X8Y154_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000055555544)
  ) CLBLM_R_X7Y154_SLICE_X8Y154_DLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.I4(CLBLL_L_X4Y153_SLICE_X4Y153_AO6),
.I5(CLBLM_R_X7Y154_SLICE_X8Y154_AQ),
.O5(CLBLM_R_X7Y154_SLICE_X8Y154_DO5),
.O6(CLBLM_R_X7Y154_SLICE_X8Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000ff0ff101)
  ) CLBLM_R_X7Y154_SLICE_X8Y154_CLUT (
.I0(CLBLM_R_X7Y148_SLICE_X8Y148_AQ),
.I1(CLBLM_R_X7Y148_SLICE_X8Y148_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y151_SLICE_X4Y151_CQ),
.I4(CLBLM_L_X8Y154_SLICE_X10Y154_A5Q),
.I5(CLBLM_L_X8Y158_SLICE_X10Y158_AQ),
.O5(CLBLM_R_X7Y154_SLICE_X8Y154_CO5),
.O6(CLBLM_R_X7Y154_SLICE_X8Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ff54ff54)
  ) CLBLM_R_X7Y154_SLICE_X8Y154_BLUT (
.I0(CLBLM_R_X7Y155_SLICE_X8Y155_CO6),
.I1(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.I2(CLBLM_L_X8Y157_SLICE_X11Y157_AQ),
.I3(CLBLM_R_X7Y158_SLICE_X8Y158_CO5),
.I4(CLBLM_R_X5Y154_SLICE_X6Y154_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y154_SLICE_X8Y154_BO5),
.O6(CLBLM_R_X7Y154_SLICE_X8Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f2000200550055)
  ) CLBLM_R_X7Y154_SLICE_X8Y154_ALUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I1(CLBLM_R_X7Y154_SLICE_X8Y154_DO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLL_L_X4Y150_SLICE_X4Y150_CQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y154_SLICE_X8Y154_AO5),
.O6(CLBLM_R_X7Y154_SLICE_X8Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y154_SLICE_X9Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y154_SLICE_X9Y154_AO6),
.Q(CLBLM_R_X7Y154_SLICE_X9Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y154_SLICE_X9Y154_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y154_SLICE_X9Y154_BO6),
.Q(CLBLM_R_X7Y154_SLICE_X9Y154_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y154_SLICE_X9Y154_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y154_SLICE_X9Y154_CO6),
.Q(CLBLM_R_X7Y154_SLICE_X9Y154_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f1ef0f0f0f0)
  ) CLBLM_R_X7Y154_SLICE_X9Y154_DLUT (
.I0(CLBLM_R_X3Y155_SLICE_X3Y155_AO6),
.I1(CLBLM_R_X13Y155_SLICE_X19Y155_AO6),
.I2(CLBLM_R_X7Y148_SLICE_X9Y148_BQ),
.I3(CLBLM_R_X7Y155_SLICE_X9Y155_DO6),
.I4(CLBLM_R_X5Y156_SLICE_X6Y156_AO6),
.I5(CLBLM_R_X13Y154_SLICE_X19Y154_AQ),
.O5(CLBLM_R_X7Y154_SLICE_X9Y154_DO5),
.O6(CLBLM_R_X7Y154_SLICE_X9Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haabeaabe00140014)
  ) CLBLM_R_X7Y154_SLICE_X9Y154_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y150_SLICE_X4Y150_CQ),
.I2(CLBLM_L_X8Y153_SLICE_X10Y153_CO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(CLBLM_L_X10Y154_SLICE_X12Y154_AQ),
.O5(CLBLM_R_X7Y154_SLICE_X9Y154_CO5),
.O6(CLBLM_R_X7Y154_SLICE_X9Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0fcfc0f000c0c)
  ) CLBLM_R_X7Y154_SLICE_X9Y154_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y154_SLICE_X9Y154_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y152_SLICE_X7Y152_CQ),
.I4(CLBLM_R_X5Y152_SLICE_X6Y152_CO5),
.I5(CLBLM_L_X8Y154_SLICE_X10Y154_B5Q),
.O5(CLBLM_R_X7Y154_SLICE_X9Y154_BO5),
.O6(CLBLM_R_X7Y154_SLICE_X9Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ffa0af000fa0a)
  ) CLBLM_R_X7Y154_SLICE_X9Y154_ALUT (
.I0(CLBLM_R_X7Y154_SLICE_X9Y154_AQ),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y146_SLICE_X15Y146_AQ),
.I4(CLBLM_R_X5Y152_SLICE_X6Y152_CO5),
.I5(CLBLL_L_X4Y150_SLICE_X4Y150_CQ),
.O5(CLBLM_R_X7Y154_SLICE_X9Y154_AO5),
.O6(CLBLM_R_X7Y154_SLICE_X9Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y155_SLICE_X8Y155_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y155_SLICE_X8Y155_AO5),
.Q(CLBLM_R_X7Y155_SLICE_X8Y155_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y155_SLICE_X8Y155_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y155_SLICE_X8Y155_AO6),
.Q(CLBLM_R_X7Y155_SLICE_X8Y155_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000f000f0)
  ) CLBLM_R_X7Y155_SLICE_X8Y155_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X7Y158_SLICE_X8Y158_BQ),
.I3(CLBLM_R_X7Y156_SLICE_X8Y156_CQ),
.I4(1'b1),
.I5(CLBLM_R_X7Y156_SLICE_X8Y156_BQ),
.O5(CLBLM_R_X7Y155_SLICE_X8Y155_DO5),
.O6(CLBLM_R_X7Y155_SLICE_X8Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000040)
  ) CLBLM_R_X7Y155_SLICE_X8Y155_CLUT (
.I0(CLBLM_R_X7Y152_SLICE_X8Y152_AQ),
.I1(CLBLM_R_X7Y155_SLICE_X8Y155_AQ),
.I2(CLBLM_R_X7Y158_SLICE_X8Y158_BQ),
.I3(CLBLM_R_X7Y156_SLICE_X8Y156_CQ),
.I4(CLBLM_L_X8Y154_SLICE_X10Y154_A5Q),
.I5(CLBLM_R_X7Y156_SLICE_X8Y156_BQ),
.O5(CLBLM_R_X7Y155_SLICE_X8Y155_CO5),
.O6(CLBLM_R_X7Y155_SLICE_X8Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0e0f00001100)
  ) CLBLM_R_X7Y155_SLICE_X8Y155_BLUT (
.I0(CLBLM_R_X7Y156_SLICE_X8Y156_CQ),
.I1(CLBLM_R_X7Y156_SLICE_X8Y156_BQ),
.I2(CLBLM_R_X7Y158_SLICE_X8Y158_CO5),
.I3(CLBLM_R_X7Y158_SLICE_X8Y158_BQ),
.I4(CLBLM_R_X7Y152_SLICE_X8Y152_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y155_SLICE_X8Y155_BO5),
.O6(CLBLM_R_X7Y155_SLICE_X8Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaaafaaac0c0cfcf)
  ) CLBLM_R_X7Y155_SLICE_X8Y155_ALUT (
.I0(CLBLM_R_X7Y158_SLICE_X8Y158_DO6),
.I1(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y154_SLICE_X11Y154_A5Q),
.I4(CLBLL_L_X4Y153_SLICE_X4Y153_AO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y155_SLICE_X8Y155_AO5),
.O6(CLBLM_R_X7Y155_SLICE_X8Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y155_SLICE_X9Y155_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y155_SLICE_X9Y155_CO5),
.Q(CLBLM_R_X7Y155_SLICE_X9Y155_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y155_SLICE_X9Y155_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y155_SLICE_X9Y155_AO6),
.Q(CLBLM_R_X7Y155_SLICE_X9Y155_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y155_SLICE_X9Y155_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y155_SLICE_X9Y155_BO6),
.Q(CLBLM_R_X7Y155_SLICE_X9Y155_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0aceffff0ace0ace)
  ) CLBLM_R_X7Y155_SLICE_X9Y155_DLUT (
.I0(CLBLM_L_X8Y155_SLICE_X10Y155_AQ),
.I1(CLBLM_L_X8Y156_SLICE_X10Y156_AQ),
.I2(CLBLM_R_X3Y153_SLICE_X3Y153_AO6),
.I3(CLBLM_R_X3Y157_SLICE_X2Y157_AO5),
.I4(CLBLL_L_X2Y155_SLICE_X1Y155_BO5),
.I5(CLBLM_L_X8Y156_SLICE_X10Y156_BQ),
.O5(CLBLM_R_X7Y155_SLICE_X9Y155_DO5),
.O6(CLBLM_R_X7Y155_SLICE_X9Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f0f0b3a0b3a0)
  ) CLBLM_R_X7Y155_SLICE_X9Y155_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLL_L_X4Y149_SLICE_X4Y149_CO6),
.I2(CLBLM_L_X8Y156_SLICE_X11Y156_AQ),
.I3(CLBLM_R_X7Y155_SLICE_X9Y155_A5Q),
.I4(CLBLM_R_X7Y155_SLICE_X8Y155_CO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y155_SLICE_X9Y155_CO5),
.O6(CLBLM_R_X7Y155_SLICE_X9Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f0fdf805000d08)
  ) CLBLM_R_X7Y155_SLICE_X9Y155_BLUT (
.I0(CLBLM_R_X7Y155_SLICE_X8Y155_CO6),
.I1(CLBLM_R_X7Y155_SLICE_X9Y155_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.I4(CLBLM_R_X7Y158_SLICE_X8Y158_CO5),
.I5(CLBLM_R_X5Y149_SLICE_X7Y149_CQ),
.O5(CLBLM_R_X7Y155_SLICE_X9Y155_BO5),
.O6(CLBLM_R_X7Y155_SLICE_X9Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafafafafacafaf)
  ) CLBLM_R_X7Y155_SLICE_X9Y155_ALUT (
.I0(CLBLM_L_X10Y154_SLICE_X12Y154_A5Q),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLL_L_X4Y158_SLICE_X4Y158_AO6),
.I4(RIOB33_X105Y135_IOB_X1Y136_I),
.I5(RIOB33_X105Y135_IOB_X1Y135_I),
.O5(CLBLM_R_X7Y155_SLICE_X9Y155_AO5),
.O6(CLBLM_R_X7Y155_SLICE_X9Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y156_SLICE_X8Y156_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y156_SLICE_X8Y156_AO6),
.Q(CLBLM_R_X7Y156_SLICE_X8Y156_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y156_SLICE_X8Y156_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y156_SLICE_X8Y156_BO6),
.Q(CLBLM_R_X7Y156_SLICE_X8Y156_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y156_SLICE_X8Y156_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y156_SLICE_X8Y156_CO6),
.Q(CLBLM_R_X7Y156_SLICE_X8Y156_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y156_SLICE_X8Y156_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y156_SLICE_X8Y156_DO6),
.Q(CLBLM_R_X7Y156_SLICE_X8Y156_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaff0055aafa0050)
  ) CLBLM_R_X7Y156_SLICE_X8Y156_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X7Y156_SLICE_X8Y156_DQ),
.I3(CLBLL_L_X4Y147_SLICE_X4Y147_BO6),
.I4(CLBLM_L_X8Y159_SLICE_X10Y159_AQ),
.I5(CLBLM_R_X7Y147_SLICE_X9Y147_A5Q),
.O5(CLBLM_R_X7Y156_SLICE_X8Y156_DO5),
.O6(CLBLM_R_X7Y156_SLICE_X8Y156_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb1a0b1a0e4a0e4a0)
  ) CLBLM_R_X7Y156_SLICE_X8Y156_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y156_SLICE_X8Y156_CQ),
.I2(CLBLM_R_X7Y157_SLICE_X8Y157_DQ),
.I3(CLBLM_R_X7Y155_SLICE_X8Y155_BO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y158_SLICE_X8Y158_BQ),
.O5(CLBLM_R_X7Y156_SLICE_X8Y156_CO5),
.O6(CLBLM_R_X7Y156_SLICE_X8Y156_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf9fc090cf0f00000)
  ) CLBLM_R_X7Y156_SLICE_X8Y156_BLUT (
.I0(CLBLM_R_X7Y156_SLICE_X8Y156_CQ),
.I1(CLBLM_R_X7Y156_SLICE_X8Y156_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y158_SLICE_X8Y158_BQ),
.I4(CLBLM_R_X7Y156_SLICE_X9Y156_AQ),
.I5(CLBLM_R_X7Y155_SLICE_X8Y155_BO6),
.O5(CLBLM_R_X7Y156_SLICE_X8Y156_BO5),
.O6(CLBLM_R_X7Y156_SLICE_X8Y156_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf5ccffcca0cc00)
  ) CLBLM_R_X7Y156_SLICE_X8Y156_ALUT (
.I0(CLBLM_L_X10Y151_SLICE_X12Y151_CQ),
.I1(CLBLM_L_X8Y157_SLICE_X11Y157_CQ),
.I2(CLBLM_R_X7Y156_SLICE_X8Y156_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y151_SLICE_X4Y151_BQ),
.I5(CLBLM_L_X10Y148_SLICE_X13Y148_AQ),
.O5(CLBLM_R_X7Y156_SLICE_X8Y156_AO5),
.O6(CLBLM_R_X7Y156_SLICE_X8Y156_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y156_SLICE_X9Y156_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y156_SLICE_X9Y156_AO6),
.Q(CLBLM_R_X7Y156_SLICE_X9Y156_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y156_SLICE_X9Y156_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y156_SLICE_X9Y156_BO6),
.Q(CLBLM_R_X7Y156_SLICE_X9Y156_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y156_SLICE_X9Y156_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y156_SLICE_X9Y156_CO6),
.Q(CLBLM_R_X7Y156_SLICE_X9Y156_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4af000005af00000)
  ) CLBLM_R_X7Y156_SLICE_X9Y156_DLUT (
.I0(CLBLM_R_X7Y155_SLICE_X8Y155_AQ),
.I1(CLBLM_L_X10Y159_SLICE_X12Y159_AO6),
.I2(CLBLM_L_X8Y154_SLICE_X10Y154_A5Q),
.I3(CLBLM_R_X7Y155_SLICE_X8Y155_BO5),
.I4(CLBLL_L_X4Y156_SLICE_X4Y156_AO5),
.I5(CLBLM_L_X8Y158_SLICE_X10Y158_AQ),
.O5(CLBLM_R_X7Y156_SLICE_X9Y156_DO5),
.O6(CLBLM_R_X7Y156_SLICE_X9Y156_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44ee44fa50fa50)
  ) CLBLM_R_X7Y156_SLICE_X9Y156_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y156_SLICE_X9Y156_CQ),
.I2(CLBLM_R_X5Y147_SLICE_X7Y147_C5Q),
.I3(CLBLM_R_X11Y157_SLICE_X14Y157_AQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y147_SLICE_X4Y147_BO6),
.O5(CLBLM_R_X7Y156_SLICE_X9Y156_CO5),
.O6(CLBLM_R_X7Y156_SLICE_X9Y156_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000303ff000303)
  ) CLBLM_R_X7Y156_SLICE_X9Y156_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X8Y152_SLICE_X11Y152_AO6),
.I3(CLBLM_L_X8Y156_SLICE_X10Y156_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y156_SLICE_X9Y156_BO5),
.O6(CLBLM_R_X7Y156_SLICE_X9Y156_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00d8d8ff00d8d8)
  ) CLBLM_R_X7Y156_SLICE_X9Y156_ALUT (
.I0(CLBLM_R_X5Y152_SLICE_X6Y152_CO5),
.I1(CLBLM_L_X10Y157_SLICE_X12Y157_AQ),
.I2(CLBLM_R_X7Y156_SLICE_X9Y156_AQ),
.I3(CLBLM_L_X12Y155_SLICE_X17Y155_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y156_SLICE_X9Y156_AO5),
.O6(CLBLM_R_X7Y156_SLICE_X9Y156_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y157_SLICE_X8Y157_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y157_SLICE_X8Y157_AO6),
.Q(CLBLM_R_X7Y157_SLICE_X8Y157_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y157_SLICE_X8Y157_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y157_SLICE_X8Y157_BO6),
.Q(CLBLM_R_X7Y157_SLICE_X8Y157_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y157_SLICE_X8Y157_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y157_SLICE_X8Y157_CO6),
.Q(CLBLM_R_X7Y157_SLICE_X8Y157_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y157_SLICE_X8Y157_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y157_SLICE_X8Y157_DO6),
.Q(CLBLM_R_X7Y157_SLICE_X8Y157_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfc3030eeee2222)
  ) CLBLM_R_X7Y157_SLICE_X8Y157_DLUT (
.I0(CLBLM_L_X8Y157_SLICE_X11Y157_BQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y157_SLICE_X8Y157_DQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y157_SLICE_X7Y157_DQ),
.I5(CLBLM_R_X5Y152_SLICE_X6Y152_CO5),
.O5(CLBLM_R_X7Y157_SLICE_X8Y157_DO5),
.O6(CLBLM_R_X7Y157_SLICE_X8Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888b8b88888b8b8)
  ) CLBLM_R_X7Y157_SLICE_X8Y157_CLUT (
.I0(CLBLM_R_X11Y155_SLICE_X14Y155_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y157_SLICE_X8Y157_BQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y159_SLICE_X8Y159_BO5),
.I5(1'b1),
.O5(CLBLM_R_X7Y157_SLICE_X8Y157_CO5),
.O6(CLBLM_R_X7Y157_SLICE_X8Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc5050cccc5050)
  ) CLBLM_R_X7Y157_SLICE_X8Y157_BLUT (
.I0(CLBLM_R_X7Y159_SLICE_X8Y159_BO5),
.I1(CLBLM_L_X10Y145_SLICE_X12Y145_CQ),
.I2(CLBLM_R_X7Y157_SLICE_X8Y157_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y157_SLICE_X8Y157_BO5),
.O6(CLBLM_R_X7Y157_SLICE_X8Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffa0f0afffa0f0a)
  ) CLBLM_R_X7Y157_SLICE_X8Y157_ALUT (
.I0(CLBLM_R_X7Y159_SLICE_X8Y159_BO5),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y158_SLICE_X8Y158_BQ),
.I4(CLBLM_L_X8Y156_SLICE_X11Y156_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X7Y157_SLICE_X8Y157_AO5),
.O6(CLBLM_R_X7Y157_SLICE_X8Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y157_SLICE_X9Y157_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y157_SLICE_X9Y157_AO6),
.Q(CLBLM_R_X7Y157_SLICE_X9Y157_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y157_SLICE_X9Y157_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y157_SLICE_X9Y157_BO6),
.Q(CLBLM_R_X7Y157_SLICE_X9Y157_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y157_SLICE_X9Y157_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y157_SLICE_X9Y157_CO6),
.Q(CLBLM_R_X7Y157_SLICE_X9Y157_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y157_SLICE_X9Y157_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y157_SLICE_X9Y157_DO6),
.Q(CLBLM_R_X7Y157_SLICE_X9Y157_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff50ff5000500050)
  ) CLBLM_R_X7Y157_SLICE_X9Y157_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(1'b1),
.I2(CLBLM_R_X7Y157_SLICE_X9Y157_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(CLBLM_R_X7Y158_SLICE_X8Y158_BQ),
.O5(CLBLM_R_X7Y157_SLICE_X9Y157_DO5),
.O6(CLBLM_R_X7Y157_SLICE_X9Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa50ee44ee44)
  ) CLBLM_R_X7Y157_SLICE_X9Y157_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y157_SLICE_X9Y157_CQ),
.I2(CLBLM_R_X7Y152_SLICE_X8Y152_A5Q),
.I3(CLBLM_L_X10Y153_SLICE_X12Y153_BQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y152_SLICE_X6Y152_CO5),
.O5(CLBLM_R_X7Y157_SLICE_X9Y157_CO5),
.O6(CLBLM_R_X7Y157_SLICE_X9Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fe000ef0fe000e)
  ) CLBLM_R_X7Y157_SLICE_X9Y157_BLUT (
.I0(CLBLM_R_X5Y157_SLICE_X7Y157_DQ),
.I1(CLBLM_R_X7Y157_SLICE_X9Y157_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X5Y152_SLICE_X6Y152_CO5),
.I4(CLBLM_L_X12Y156_SLICE_X16Y156_BQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y157_SLICE_X9Y157_BO5),
.O6(CLBLM_R_X7Y157_SLICE_X9Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff500050ffcc00cc)
  ) CLBLM_R_X7Y157_SLICE_X9Y157_ALUT (
.I0(CLBLM_R_X7Y158_SLICE_X8Y158_CO5),
.I1(CLBLM_R_X7Y155_SLICE_X9Y155_BQ),
.I2(CLBLM_R_X7Y157_SLICE_X9Y157_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLL_L_X4Y155_SLICE_X4Y155_BQ),
.I5(CLBLM_R_X7Y155_SLICE_X8Y155_CO6),
.O5(CLBLM_R_X7Y157_SLICE_X9Y157_AO5),
.O6(CLBLM_R_X7Y157_SLICE_X9Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y158_SLICE_X8Y158_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y158_SLICE_X8Y158_AO6),
.Q(CLBLM_R_X7Y158_SLICE_X8Y158_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y158_SLICE_X8Y158_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y158_SLICE_X8Y158_BO6),
.Q(CLBLM_R_X7Y158_SLICE_X8Y158_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000000dfda)
  ) CLBLM_R_X7Y158_SLICE_X8Y158_DLUT (
.I0(CLBLM_L_X8Y157_SLICE_X11Y157_AQ),
.I1(CLBLM_R_X7Y155_SLICE_X8Y155_CO6),
.I2(CLBLM_R_X7Y155_SLICE_X8Y155_AQ),
.I3(CLBLM_R_X7Y158_SLICE_X8Y158_CO6),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X7Y158_SLICE_X8Y158_DO5),
.O6(CLBLM_R_X7Y158_SLICE_X8Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0100000000000101)
  ) CLBLM_R_X7Y158_SLICE_X8Y158_CLUT (
.I0(CLBLM_R_X7Y148_SLICE_X8Y148_BQ),
.I1(CLBLM_R_X7Y148_SLICE_X8Y148_AQ),
.I2(CLBLM_L_X8Y154_SLICE_X10Y154_A5Q),
.I3(CLBLM_R_X7Y155_SLICE_X8Y155_BO5),
.I4(CLBLM_L_X8Y158_SLICE_X10Y158_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y158_SLICE_X8Y158_CO5),
.O6(CLBLM_R_X7Y158_SLICE_X8Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5c5c0c0c5c5c0c0)
  ) CLBLM_R_X7Y158_SLICE_X8Y158_BLUT (
.I0(CLBLM_R_X7Y159_SLICE_X8Y159_BO5),
.I1(CLBLL_L_X4Y155_SLICE_X5Y155_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_R_X7Y159_SLICE_X8Y159_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y158_SLICE_X8Y158_BO5),
.O6(CLBLM_R_X7Y158_SLICE_X8Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccfff0cccc00f0)
  ) CLBLM_R_X7Y158_SLICE_X8Y158_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y156_SLICE_X8Y156_AQ),
.I2(CLBLM_R_X7Y158_SLICE_X8Y158_AQ),
.I3(CLBLM_R_X5Y152_SLICE_X6Y152_CO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X8Y153_SLICE_X11Y153_DQ),
.O5(CLBLM_R_X7Y158_SLICE_X8Y158_AO5),
.O6(CLBLM_R_X7Y158_SLICE_X8Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y158_SLICE_X9Y158_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y158_SLICE_X9Y158_AO6),
.Q(CLBLM_R_X7Y158_SLICE_X9Y158_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff4fffffff4fff4)
  ) CLBLM_R_X7Y158_SLICE_X9Y158_DLUT (
.I0(CLBLM_R_X3Y157_SLICE_X2Y157_AO5),
.I1(CLBLM_R_X5Y151_SLICE_X7Y151_BQ),
.I2(CLBLM_R_X7Y158_SLICE_X9Y158_BO6),
.I3(CLBLM_R_X7Y158_SLICE_X9Y158_CO6),
.I4(CLBLL_L_X2Y155_SLICE_X1Y155_BO5),
.I5(CLBLM_R_X7Y156_SLICE_X8Y156_AQ),
.O5(CLBLM_R_X7Y158_SLICE_X9Y158_DO5),
.O6(CLBLM_R_X7Y158_SLICE_X9Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000080000)
  ) CLBLM_R_X7Y158_SLICE_X9Y158_CLUT (
.I0(CLBLM_L_X10Y158_SLICE_X12Y158_AQ),
.I1(RIOB33_X105Y131_IOB_X1Y132_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y133_IOB_X1Y134_I),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(CLBLL_L_X4Y157_SLICE_X4Y157_CO5),
.O5(CLBLM_R_X7Y158_SLICE_X9Y158_CO5),
.O6(CLBLM_R_X7Y158_SLICE_X9Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000008)
  ) CLBLM_R_X7Y158_SLICE_X9Y158_BLUT (
.I0(RIOB33_X105Y131_IOB_X1Y132_I),
.I1(CLBLM_R_X13Y150_SLICE_X18Y150_AQ),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(CLBLL_L_X4Y157_SLICE_X4Y157_CO5),
.I4(RIOB33_X105Y131_IOB_X1Y131_I),
.I5(RIOB33_X105Y133_IOB_X1Y134_I),
.O5(CLBLM_R_X7Y158_SLICE_X9Y158_BO5),
.O6(CLBLM_R_X7Y158_SLICE_X9Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaafcfcaaaa3030)
  ) CLBLM_R_X7Y158_SLICE_X9Y158_ALUT (
.I0(CLBLM_L_X8Y154_SLICE_X10Y154_A5Q),
.I1(CLBLM_R_X5Y152_SLICE_X6Y152_CO5),
.I2(CLBLM_R_X7Y158_SLICE_X9Y158_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y154_SLICE_X9Y154_CQ),
.O5(CLBLM_R_X7Y158_SLICE_X9Y158_AO5),
.O6(CLBLM_R_X7Y158_SLICE_X9Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X7Y159_SLICE_X8Y159_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X7Y159_SLICE_X8Y159_AO6),
.Q(CLBLM_R_X7Y159_SLICE_X8Y159_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y159_SLICE_X8Y159_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y159_SLICE_X8Y159_DO5),
.O6(CLBLM_R_X7Y159_SLICE_X8Y159_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y159_SLICE_X8Y159_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y159_SLICE_X8Y159_CO5),
.O6(CLBLM_R_X7Y159_SLICE_X8Y159_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc030303022222233)
  ) CLBLM_R_X7Y159_SLICE_X8Y159_BLUT (
.I0(CLBLM_L_X8Y154_SLICE_X10Y154_A5Q),
.I1(CLBLM_L_X8Y158_SLICE_X10Y158_AQ),
.I2(CLBLM_L_X10Y159_SLICE_X12Y159_AO6),
.I3(CLBLM_R_X7Y148_SLICE_X8Y148_BQ),
.I4(CLBLM_R_X7Y148_SLICE_X8Y148_AQ),
.I5(1'b1),
.O5(CLBLM_R_X7Y159_SLICE_X8Y159_BO5),
.O6(CLBLM_R_X7Y159_SLICE_X8Y159_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5c5c5c5c0c0c0c0)
  ) CLBLM_R_X7Y159_SLICE_X8Y159_ALUT (
.I0(CLBLM_R_X7Y159_SLICE_X8Y159_BO5),
.I1(CLBLM_R_X11Y158_SLICE_X15Y158_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X7Y157_SLICE_X8Y157_CQ),
.O5(CLBLM_R_X7Y159_SLICE_X8Y159_AO5),
.O6(CLBLM_R_X7Y159_SLICE_X8Y159_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000001000000)
  ) CLBLM_R_X7Y159_SLICE_X9Y159_DLUT (
.I0(RIOB33_X105Y133_IOB_X1Y134_I),
.I1(RIOB33_X105Y131_IOB_X1Y131_I),
.I2(RIOB33_X105Y133_IOB_X1Y133_I),
.I3(RIOB33_X105Y131_IOB_X1Y132_I),
.I4(CLBLM_R_X11Y159_SLICE_X14Y159_CQ),
.I5(CLBLL_L_X4Y157_SLICE_X4Y157_CO5),
.O5(CLBLM_R_X7Y159_SLICE_X9Y159_DO5),
.O6(CLBLM_R_X7Y159_SLICE_X9Y159_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00ff30c50af5fa0)
  ) CLBLM_R_X7Y159_SLICE_X9Y159_CLUT (
.I0(CLBLM_R_X7Y148_SLICE_X8Y148_AQ),
.I1(CLBLM_R_X7Y148_SLICE_X8Y148_BQ),
.I2(CLBLM_L_X8Y150_SLICE_X11Y150_CQ),
.I3(CLBLM_R_X3Y152_SLICE_X3Y152_BO5),
.I4(CLBLM_L_X8Y154_SLICE_X10Y154_A5Q),
.I5(CLBLM_L_X8Y158_SLICE_X10Y158_AQ),
.O5(CLBLM_R_X7Y159_SLICE_X9Y159_CO5),
.O6(CLBLM_R_X7Y159_SLICE_X9Y159_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffef554400000000)
  ) CLBLM_R_X7Y159_SLICE_X9Y159_BLUT (
.I0(CLBLM_L_X8Y154_SLICE_X10Y154_A5Q),
.I1(CLBLM_R_X7Y148_SLICE_X8Y148_AQ),
.I2(CLBLM_R_X7Y155_SLICE_X8Y155_AQ),
.I3(CLBLM_R_X7Y148_SLICE_X8Y148_BQ),
.I4(CLBLM_L_X8Y158_SLICE_X10Y158_AQ),
.I5(CLBLM_R_X7Y157_SLICE_X8Y157_CQ),
.O5(CLBLM_R_X7Y159_SLICE_X9Y159_BO5),
.O6(CLBLM_R_X7Y159_SLICE_X9Y159_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f3f0f050735050)
  ) CLBLM_R_X7Y159_SLICE_X9Y159_ALUT (
.I0(CLBLM_R_X7Y159_SLICE_X9Y159_BO6),
.I1(CLBLM_R_X7Y148_SLICE_X8Y148_AQ),
.I2(CLBLM_L_X8Y159_SLICE_X10Y159_AQ),
.I3(CLBLM_L_X8Y158_SLICE_X10Y158_AQ),
.I4(CLBLM_R_X7Y148_SLICE_X8Y148_BQ),
.I5(CLBLM_R_X7Y159_SLICE_X9Y159_CO6),
.O5(CLBLM_R_X7Y159_SLICE_X9Y159_AO5),
.O6(CLBLM_R_X7Y159_SLICE_X9Y159_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y144_SLICE_X14Y144_DO5),
.O6(CLBLM_R_X11Y144_SLICE_X14Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y144_SLICE_X14Y144_CO5),
.O6(CLBLM_R_X11Y144_SLICE_X14Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y144_SLICE_X14Y144_BO5),
.O6(CLBLM_R_X11Y144_SLICE_X14Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y144_SLICE_X14Y144_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y144_SLICE_X14Y144_AO5),
.O6(CLBLM_R_X11Y144_SLICE_X14Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y144_SLICE_X15Y144_AO5),
.Q(CLBLM_R_X11Y144_SLICE_X15Y144_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y144_SLICE_X15Y144_AO6),
.Q(CLBLM_R_X11Y144_SLICE_X15Y144_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y144_SLICE_X15Y144_DO5),
.O6(CLBLM_R_X11Y144_SLICE_X15Y144_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y144_SLICE_X15Y144_CO5),
.O6(CLBLM_R_X11Y144_SLICE_X15Y144_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y144_SLICE_X15Y144_BO5),
.O6(CLBLM_R_X11Y144_SLICE_X15Y144_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5a0a0dddd8888)
  ) CLBLM_R_X11Y144_SLICE_X15Y144_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y157_SLICE_X17Y157_BQ),
.I2(CLBLM_R_X5Y146_SLICE_X6Y146_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y125_IOB_X1Y126_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y144_SLICE_X15Y144_AO5),
.O6(CLBLM_R_X11Y144_SLICE_X15Y144_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y146_SLICE_X14Y146_AO6),
.Q(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y146_SLICE_X14Y146_BO6),
.Q(CLBLM_R_X11Y146_SLICE_X14Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y146_SLICE_X14Y146_CO6),
.Q(CLBLM_R_X11Y146_SLICE_X14Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y146_SLICE_X14Y146_DO6),
.Q(CLBLM_R_X11Y146_SLICE_X14Y146_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00ffcccc00f0)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y147_SLICE_X13Y147_BQ),
.I2(CLBLM_R_X11Y146_SLICE_X14Y146_DQ),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y146_SLICE_X15Y146_BQ),
.O5(CLBLM_R_X11Y146_SLICE_X14Y146_DO5),
.O6(CLBLM_R_X11Y146_SLICE_X14Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff8f008fffcf00cf)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_CLUT (
.I0(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.I1(CLBLM_R_X11Y146_SLICE_X14Y146_CQ),
.I2(CLBLM_R_X13Y147_SLICE_X18Y147_CO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y159_SLICE_X14Y159_CQ),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_R_X11Y146_SLICE_X14Y146_CO5),
.O6(CLBLM_R_X11Y146_SLICE_X14Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8fcf8fc080c080c)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_BLUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I1(CLBLM_R_X11Y146_SLICE_X14Y146_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(1'b1),
.I5(CLBLM_L_X10Y150_SLICE_X13Y150_B5Q),
.O5(CLBLM_R_X11Y146_SLICE_X14Y146_BO5),
.O6(CLBLM_R_X11Y146_SLICE_X14Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffccf0ccaacca0)
  ) CLBLM_R_X11Y146_SLICE_X14Y146_ALUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I1(CLBLM_R_X11Y148_SLICE_X14Y148_AQ),
.I2(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y150_SLICE_X13Y150_B5Q),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X11Y146_SLICE_X14Y146_AO5),
.O6(CLBLM_R_X11Y146_SLICE_X14Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y146_SLICE_X15Y146_AO6),
.Q(CLBLM_R_X11Y146_SLICE_X15Y146_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y146_SLICE_X15Y146_BO6),
.Q(CLBLM_R_X11Y146_SLICE_X15Y146_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y146_SLICE_X15Y146_CO6),
.Q(CLBLM_R_X11Y146_SLICE_X15Y146_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfe01ff005f5fffff)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_DLUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_CQ),
.I1(CLBLM_L_X10Y145_SLICE_X13Y145_BQ),
.I2(CLBLM_L_X10Y146_SLICE_X12Y146_C5Q),
.I3(CLBLM_L_X10Y147_SLICE_X12Y147_CQ),
.I4(CLBLM_L_X10Y146_SLICE_X12Y146_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y146_SLICE_X15Y146_DO5),
.O6(CLBLM_R_X11Y146_SLICE_X15Y146_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0afa0afa0aca0ac)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_CLUT (
.I0(CLBLM_R_X11Y154_SLICE_X15Y154_BQ),
.I1(CLBLM_R_X11Y146_SLICE_X15Y146_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.I4(1'b1),
.I5(CLBLM_L_X8Y146_SLICE_X11Y146_AQ),
.O5(CLBLM_R_X11Y146_SLICE_X15Y146_CO5),
.O6(CLBLM_R_X11Y146_SLICE_X15Y146_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaee00550044)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y146_SLICE_X15Y146_BQ),
.I2(1'b1),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_DO6),
.I4(CLBLM_L_X8Y146_SLICE_X11Y146_CQ),
.I5(CLBLM_R_X11Y153_SLICE_X15Y153_BQ),
.O5(CLBLM_R_X11Y146_SLICE_X15Y146_BO5),
.O6(CLBLM_R_X11Y146_SLICE_X15Y146_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haafe0054aafe0054)
  ) CLBLM_R_X11Y146_SLICE_X15Y146_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y147_SLICE_X12Y147_AQ),
.I2(CLBLM_R_X11Y146_SLICE_X15Y146_AQ),
.I3(CLBLM_R_X7Y146_SLICE_X9Y146_DO6),
.I4(CLBLM_L_X12Y147_SLICE_X16Y147_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y146_SLICE_X15Y146_AO5),
.O6(CLBLM_R_X11Y146_SLICE_X15Y146_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2010201002010201)
  ) CLBLM_R_X11Y147_SLICE_X14Y147_DLUT (
.I0(CLBLM_R_X11Y146_SLICE_X15Y146_AQ),
.I1(CLBLM_L_X10Y146_SLICE_X13Y146_DO6),
.I2(CLBLM_R_X11Y152_SLICE_X14Y152_B5Q),
.I3(CLBLM_L_X12Y157_SLICE_X17Y157_A5Q),
.I4(1'b1),
.I5(CLBLM_L_X10Y147_SLICE_X12Y147_AQ),
.O5(CLBLM_R_X11Y147_SLICE_X14Y147_DO5),
.O6(CLBLM_R_X11Y147_SLICE_X14Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0201000020100000)
  ) CLBLM_R_X11Y147_SLICE_X14Y147_CLUT (
.I0(CLBLM_L_X12Y149_SLICE_X16Y149_B5Q),
.I1(CLBLM_R_X11Y147_SLICE_X15Y147_CO6),
.I2(CLBLM_R_X13Y153_SLICE_X18Y153_CQ),
.I3(CLBLM_L_X8Y147_SLICE_X11Y147_AQ),
.I4(CLBLM_R_X11Y147_SLICE_X14Y147_DO6),
.I5(CLBLM_L_X10Y147_SLICE_X13Y147_DO6),
.O5(CLBLM_R_X11Y147_SLICE_X14Y147_CO5),
.O6(CLBLM_R_X11Y147_SLICE_X14Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h010200030d0e0c0f)
  ) CLBLM_R_X11Y147_SLICE_X14Y147_BLUT (
.I0(CLBLM_R_X13Y147_SLICE_X18Y147_AO5),
.I1(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.I2(CLBLM_L_X10Y147_SLICE_X12Y147_BQ),
.I3(CLBLM_R_X11Y150_SLICE_X14Y150_AQ),
.I4(CLBLM_R_X11Y147_SLICE_X14Y147_AO6),
.I5(CLBLM_L_X10Y149_SLICE_X12Y149_CQ),
.O5(CLBLM_R_X11Y147_SLICE_X14Y147_BO5),
.O6(CLBLM_R_X11Y147_SLICE_X14Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h550055000f0f1e0f)
  ) CLBLM_R_X11Y147_SLICE_X14Y147_ALUT (
.I0(CLBLM_L_X10Y146_SLICE_X12Y146_C5Q),
.I1(CLBLM_L_X10Y146_SLICE_X12Y146_CQ),
.I2(CLBLM_L_X12Y149_SLICE_X17Y149_A5Q),
.I3(CLBLM_L_X10Y145_SLICE_X13Y145_BQ),
.I4(CLBLM_L_X10Y145_SLICE_X13Y145_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y147_SLICE_X14Y147_AO5),
.O6(CLBLM_R_X11Y147_SLICE_X14Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h77bbddee77bbddee)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_DLUT (
.I0(CLBLM_L_X8Y146_SLICE_X11Y146_AQ),
.I1(CLBLM_L_X8Y148_SLICE_X11Y148_B5Q),
.I2(1'b1),
.I3(CLBLM_L_X12Y154_SLICE_X16Y154_A5Q),
.I4(CLBLM_L_X10Y146_SLICE_X12Y146_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y147_SLICE_X15Y147_DO5),
.O6(CLBLM_R_X11Y147_SLICE_X15Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5affffffff5a)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_CLUT (
.I0(CLBLM_R_X11Y146_SLICE_X15Y146_CQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y150_SLICE_X13Y150_C5Q),
.I3(CLBLM_L_X10Y147_SLICE_X13Y147_BQ),
.I4(CLBLM_R_X11Y147_SLICE_X15Y147_DO6),
.I5(CLBLM_L_X8Y155_SLICE_X10Y155_BQ),
.O5(CLBLM_R_X11Y147_SLICE_X15Y147_CO5),
.O6(CLBLM_R_X11Y147_SLICE_X15Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1111303011110303)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_BLUT (
.I0(CLBLM_L_X10Y150_SLICE_X13Y150_C5Q),
.I1(CLBLM_L_X10Y147_SLICE_X13Y147_AQ),
.I2(CLBLM_R_X11Y153_SLICE_X15Y153_DQ),
.I3(1'b1),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.I5(CLBLM_L_X12Y147_SLICE_X16Y147_BO6),
.O5(CLBLM_R_X11Y147_SLICE_X15Y147_BO5),
.O6(CLBLM_R_X11Y147_SLICE_X15Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa5555aa3c553c)
  ) CLBLM_R_X11Y147_SLICE_X15Y147_ALUT (
.I0(CLBLM_R_X11Y152_SLICE_X14Y152_B5Q),
.I1(CLBLM_R_X11Y146_SLICE_X15Y146_DO6),
.I2(CLBLM_R_X11Y147_SLICE_X14Y147_AO5),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_BO6),
.I4(CLBLM_L_X8Y155_SLICE_X10Y155_BQ),
.I5(CLBLM_R_X3Y154_SLICE_X2Y154_AO6),
.O5(CLBLM_R_X11Y147_SLICE_X15Y147_AO5),
.O6(CLBLM_R_X11Y147_SLICE_X15Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y148_SLICE_X14Y148_AO6),
.Q(CLBLM_R_X11Y148_SLICE_X14Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y148_SLICE_X14Y148_BO6),
.Q(CLBLM_R_X11Y148_SLICE_X14Y148_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y148_SLICE_X14Y148_CO6),
.Q(CLBLM_R_X11Y148_SLICE_X14Y148_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1111111100330033)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_DLUT (
.I0(CLBLM_R_X11Y152_SLICE_X14Y152_B5Q),
.I1(CLBLM_R_X11Y148_SLICE_X14Y148_CQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y146_SLICE_X15Y146_DO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.O5(CLBLM_R_X11Y148_SLICE_X14Y148_DO5),
.O6(CLBLM_R_X11Y148_SLICE_X14Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff000000cfcf)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_CLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.I2(RIOB33_X105Y141_IOB_X1Y142_I),
.I3(CLBLM_L_X10Y151_SLICE_X12Y151_DQ),
.I4(CLBLM_R_X11Y148_SLICE_X14Y148_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y148_SLICE_X14Y148_CO5),
.O6(CLBLM_R_X11Y148_SLICE_X14Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00aaccaacc)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_BLUT (
.I0(CLBLM_L_X10Y150_SLICE_X13Y150_C5Q),
.I1(CLBLM_R_X11Y148_SLICE_X14Y148_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y148_SLICE_X14Y148_BO5),
.O6(CLBLM_R_X11Y148_SLICE_X14Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfecccc00320000)
  ) CLBLM_R_X11Y148_SLICE_X14Y148_ALUT (
.I0(CLBLM_R_X11Y148_SLICE_X14Y148_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y148_SLICE_X14Y148_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I5(CLBLM_L_X8Y150_SLICE_X11Y150_AQ),
.O5(CLBLM_R_X11Y148_SLICE_X14Y148_AO5),
.O6(CLBLM_R_X11Y148_SLICE_X14Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y148_SLICE_X15Y148_AO6),
.Q(CLBLM_R_X11Y148_SLICE_X15Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000f0005000700)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_DLUT (
.I0(CLBLM_R_X11Y150_SLICE_X14Y150_AQ),
.I1(CLBLM_R_X7Y148_SLICE_X9Y148_CO5),
.I2(CLBLM_R_X11Y157_SLICE_X14Y157_DO6),
.I3(CLBLM_L_X12Y152_SLICE_X16Y152_DO6),
.I4(CLBLM_R_X7Y146_SLICE_X9Y146_BO6),
.I5(CLBLM_R_X7Y146_SLICE_X8Y146_BO6),
.O5(CLBLM_R_X11Y148_SLICE_X15Y148_DO5),
.O6(CLBLM_R_X11Y148_SLICE_X15Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffccfffffffeff)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_CLUT (
.I0(CLBLM_R_X7Y148_SLICE_X9Y148_CO5),
.I1(CLBLM_L_X12Y156_SLICE_X16Y156_CO6),
.I2(CLBLM_R_X7Y146_SLICE_X9Y146_BO6),
.I3(CLBLM_L_X8Y148_SLICE_X11Y148_B5Q),
.I4(CLBLM_R_X11Y156_SLICE_X15Y156_CO6),
.I5(CLBLM_R_X7Y146_SLICE_X8Y146_BO6),
.O5(CLBLM_R_X11Y148_SLICE_X15Y148_CO5),
.O6(CLBLM_R_X11Y148_SLICE_X15Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00010a0b05040f0e)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_BLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.I1(CLBLM_L_X12Y148_SLICE_X16Y148_AO6),
.I2(CLBLM_R_X11Y148_SLICE_X15Y148_AQ),
.I3(CLBLM_L_X10Y146_SLICE_X12Y146_CQ),
.I4(CLBLM_L_X12Y149_SLICE_X16Y149_B5Q),
.I5(CLBLM_L_X10Y145_SLICE_X12Y145_CQ),
.O5(CLBLM_R_X11Y148_SLICE_X15Y148_BO5),
.O6(CLBLM_R_X11Y148_SLICE_X15Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcceeccff00220033)
  ) CLBLM_R_X11Y148_SLICE_X15Y148_ALUT (
.I0(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(1'b1),
.I3(CLBLM_R_X11Y148_SLICE_X15Y148_BO6),
.I4(RIOB33_X105Y141_IOB_X1Y142_I),
.I5(CLBLM_R_X13Y151_SLICE_X18Y151_DQ),
.O5(CLBLM_R_X11Y148_SLICE_X15Y148_AO5),
.O6(CLBLM_R_X11Y148_SLICE_X15Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y149_SLICE_X14Y149_AO6),
.Q(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y149_SLICE_X14Y149_BO6),
.Q(CLBLM_R_X11Y149_SLICE_X14Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y149_SLICE_X14Y149_CO6),
.Q(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y149_SLICE_X14Y149_DO6),
.Q(CLBLM_R_X11Y149_SLICE_X14Y149_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff003c0000003c)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_DLUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y148_SLICE_X13Y148_DO6),
.I2(CLBLM_R_X11Y149_SLICE_X14Y149_DQ),
.I3(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X13Y152_SLICE_X19Y152_AQ),
.O5(CLBLM_R_X11Y149_SLICE_X14Y149_DO5),
.O6(CLBLM_R_X11Y149_SLICE_X14Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa003c00cc)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_CLUT (
.I0(CLBLM_L_X12Y150_SLICE_X17Y150_AQ),
.I1(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.I2(CLBLM_R_X11Y149_SLICE_X14Y149_DQ),
.I3(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I4(CLBLM_L_X10Y148_SLICE_X13Y148_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y149_SLICE_X14Y149_CO5),
.O6(CLBLM_R_X11Y149_SLICE_X14Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaf0f0f0cc)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_BLUT (
.I0(CLBLM_R_X7Y157_SLICE_X9Y157_BQ),
.I1(CLBLM_R_X11Y149_SLICE_X14Y149_BQ),
.I2(CLBLM_R_X11Y148_SLICE_X14Y148_AQ),
.I3(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y149_SLICE_X14Y149_BO5),
.O6(CLBLM_R_X11Y149_SLICE_X14Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc000c0ffaa00aa)
  ) CLBLM_R_X11Y149_SLICE_X14Y149_ALUT (
.I0(CLBLM_R_X13Y151_SLICE_X18Y151_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y147_SLICE_X12Y147_BQ),
.I5(CLBLM_R_X11Y149_SLICE_X15Y149_DO6),
.O5(CLBLM_R_X11Y149_SLICE_X14Y149_AO5),
.O6(CLBLM_R_X11Y149_SLICE_X14Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y149_SLICE_X15Y149_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y149_SLICE_X15Y149_AO5),
.Q(CLBLM_R_X11Y149_SLICE_X15Y149_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y149_SLICE_X15Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X11Y149_SLICE_X15Y149_AO6),
.Q(CLBLM_R_X11Y149_SLICE_X15Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0011001100000000)
  ) CLBLM_R_X11Y149_SLICE_X15Y149_DLUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I1(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I2(1'b1),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y149_SLICE_X5Y149_AQ),
.O5(CLBLM_R_X11Y149_SLICE_X15Y149_DO5),
.O6(CLBLM_R_X11Y149_SLICE_X15Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9669966969966996)
  ) CLBLM_R_X11Y149_SLICE_X15Y149_CLUT (
.I0(CLBLM_L_X10Y151_SLICE_X12Y151_AQ),
.I1(CLBLM_R_X11Y150_SLICE_X15Y150_CO6),
.I2(CLBLM_R_X7Y148_SLICE_X9Y148_BQ),
.I3(CLBLM_L_X12Y151_SLICE_X16Y151_AQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y149_SLICE_X14Y149_BQ),
.O5(CLBLM_R_X11Y149_SLICE_X15Y149_CO5),
.O6(CLBLM_R_X11Y149_SLICE_X15Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0054540054000054)
  ) CLBLM_R_X11Y149_SLICE_X15Y149_BLUT (
.I0(CLBLM_L_X10Y149_SLICE_X13Y149_A5Q),
.I1(CLBLM_R_X13Y155_SLICE_X19Y155_AO6),
.I2(CLBLM_R_X5Y155_SLICE_X6Y155_DO6),
.I3(CLBLM_R_X13Y153_SLICE_X18Y153_AQ),
.I4(CLBLM_L_X10Y153_SLICE_X13Y153_AQ),
.I5(CLBLM_R_X11Y149_SLICE_X15Y149_CO6),
.O5(CLBLM_R_X11Y149_SLICE_X15Y149_BO5),
.O6(CLBLM_R_X11Y149_SLICE_X15Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbbb8888c0e2c0e2)
  ) CLBLM_R_X11Y149_SLICE_X15Y149_ALUT (
.I0(CLBLM_R_X13Y149_SLICE_X18Y149_CQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y149_SLICE_X14Y149_CQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y149_SLICE_X15Y149_AO5),
.O6(CLBLM_R_X11Y149_SLICE_X15Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y150_SLICE_X14Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y150_SLICE_X14Y150_AO6),
.Q(CLBLM_R_X11Y150_SLICE_X14Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffeeffee)
  ) CLBLM_R_X11Y150_SLICE_X14Y150_DLUT (
.I0(CLBLM_L_X8Y150_SLICE_X10Y150_A5Q),
.I1(CLBLM_R_X7Y151_SLICE_X8Y151_DQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y151_SLICE_X15Y151_AQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y151_SLICE_X6Y151_CQ),
.O5(CLBLM_R_X11Y150_SLICE_X14Y150_DO5),
.O6(CLBLM_R_X11Y150_SLICE_X14Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hefffefffefffefff)
  ) CLBLM_R_X11Y150_SLICE_X14Y150_CLUT (
.I0(CLBLM_R_X11Y146_SLICE_X15Y146_BQ),
.I1(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I2(CLBLM_R_X11Y146_SLICE_X14Y146_DQ),
.I3(CLBLL_L_X4Y148_SLICE_X5Y148_DQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y150_SLICE_X14Y150_CO5),
.O6(CLBLM_R_X11Y150_SLICE_X14Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffefffe)
  ) CLBLM_R_X11Y150_SLICE_X14Y150_BLUT (
.I0(CLBLM_R_X11Y150_SLICE_X14Y150_DO6),
.I1(CLBLM_R_X11Y149_SLICE_X15Y149_A5Q),
.I2(CLBLM_R_X5Y152_SLICE_X6Y152_BQ),
.I3(CLBLM_L_X10Y150_SLICE_X13Y150_AQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y152_SLICE_X12Y152_BQ),
.O5(CLBLM_R_X11Y150_SLICE_X14Y150_BO5),
.O6(CLBLM_R_X11Y150_SLICE_X14Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000fffa5550)
  ) CLBLM_R_X11Y150_SLICE_X14Y150_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X11Y150_SLICE_X14Y150_AQ),
.I3(CLBLM_L_X12Y149_SLICE_X17Y149_A5Q),
.I4(CLBLM_L_X10Y150_SLICE_X12Y150_BQ),
.I5(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.O5(CLBLM_R_X11Y150_SLICE_X14Y150_AO5),
.O6(CLBLM_R_X11Y150_SLICE_X14Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5faf5faff5faf5fa)
  ) CLBLM_R_X11Y150_SLICE_X15Y150_DLUT (
.I0(CLBLM_L_X8Y147_SLICE_X11Y147_BQ),
.I1(1'b1),
.I2(CLBLM_R_X11Y149_SLICE_X14Y149_AQ),
.I3(CLBLM_R_X13Y152_SLICE_X19Y152_AQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y155_SLICE_X14Y155_BQ),
.O5(CLBLM_R_X11Y150_SLICE_X15Y150_DO5),
.O6(CLBLM_R_X11Y150_SLICE_X15Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969696996969696)
  ) CLBLM_R_X11Y150_SLICE_X15Y150_CLUT (
.I0(CLBLM_R_X13Y150_SLICE_X19Y150_AQ),
.I1(CLBLM_R_X11Y155_SLICE_X14Y155_BQ),
.I2(CLBLM_R_X7Y149_SLICE_X8Y149_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_L_X8Y147_SLICE_X11Y147_BQ),
.O5(CLBLM_R_X11Y150_SLICE_X15Y150_CO5),
.O6(CLBLM_R_X11Y150_SLICE_X15Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000004)
  ) CLBLM_R_X11Y150_SLICE_X15Y150_BLUT (
.I0(CLBLM_R_X11Y150_SLICE_X14Y150_CO6),
.I1(CLBLM_L_X10Y149_SLICE_X12Y149_DO5),
.I2(CLBLM_R_X13Y148_SLICE_X18Y148_AQ),
.I3(CLBLM_R_X13Y149_SLICE_X19Y149_AQ),
.I4(CLBLM_R_X13Y150_SLICE_X18Y150_CQ),
.I5(CLBLL_L_X4Y157_SLICE_X4Y157_BO6),
.O5(CLBLM_R_X11Y150_SLICE_X15Y150_BO5),
.O6(CLBLM_R_X11Y150_SLICE_X15Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcec3020f0a0f0a0)
  ) CLBLM_R_X11Y150_SLICE_X15Y150_ALUT (
.I0(CLBLM_R_X11Y149_SLICE_X15Y149_A5Q),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(RIOB33_X105Y121_IOB_X1Y121_I),
.I3(CLBLM_L_X12Y150_SLICE_X16Y150_AQ),
.I4(CLBLM_R_X11Y150_SLICE_X14Y150_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y150_SLICE_X15Y150_AO5),
.O6(CLBLM_R_X11Y150_SLICE_X15Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y151_SLICE_X14Y151_AO6),
.Q(CLBLM_R_X11Y151_SLICE_X14Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y151_SLICE_X14Y151_BO6),
.Q(CLBLM_R_X11Y151_SLICE_X14Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h77bb77bbddeeddee)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_DLUT (
.I0(CLBLM_R_X7Y149_SLICE_X8Y149_BQ),
.I1(CLBLM_R_X11Y151_SLICE_X14Y151_AQ),
.I2(1'b1),
.I3(CLBLM_L_X12Y153_SLICE_X17Y153_BQ),
.I4(1'b1),
.I5(CLBLM_L_X10Y151_SLICE_X12Y151_AQ),
.O5(CLBLM_R_X11Y151_SLICE_X14Y151_DO5),
.O6(CLBLM_R_X11Y151_SLICE_X14Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_CLUT (
.I0(CLBLM_R_X7Y151_SLICE_X9Y151_C5Q),
.I1(CLBLM_L_X12Y152_SLICE_X17Y152_AQ),
.I2(CLBLM_L_X10Y151_SLICE_X13Y151_BQ),
.I3(CLBLM_L_X10Y151_SLICE_X13Y151_CQ),
.I4(CLBLM_L_X12Y151_SLICE_X17Y151_AQ),
.I5(CLBLM_L_X10Y149_SLICE_X12Y149_C5Q),
.O5(CLBLM_R_X11Y151_SLICE_X14Y151_CO5),
.O6(CLBLM_R_X11Y151_SLICE_X14Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f033003300)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X10Y153_SLICE_X13Y153_AQ),
.I3(CLBLM_L_X10Y149_SLICE_X12Y149_C5Q),
.I4(1'b1),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y151_SLICE_X14Y151_BO5),
.O6(CLBLM_R_X11Y151_SLICE_X14Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaac0ffaaaac000)
  ) CLBLM_R_X11Y151_SLICE_X14Y151_ALUT (
.I0(CLBLM_R_X5Y151_SLICE_X7Y151_AQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_R_X11Y151_SLICE_X14Y151_AQ),
.I3(CLBLM_R_X11Y149_SLICE_X15Y149_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X13Y152_SLICE_X19Y152_AQ),
.O5(CLBLM_R_X11Y151_SLICE_X14Y151_AO5),
.O6(CLBLM_R_X11Y151_SLICE_X14Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y151_SLICE_X15Y151_AO5),
.Q(CLBLM_R_X11Y151_SLICE_X15Y151_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y151_SLICE_X15Y151_AO6),
.Q(CLBLM_R_X11Y151_SLICE_X15Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y151_SLICE_X15Y151_BO6),
.Q(CLBLM_R_X11Y151_SLICE_X15Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_DLUT (
.I0(CLBLM_R_X7Y153_SLICE_X8Y153_BQ),
.I1(CLBLM_R_X11Y151_SLICE_X14Y151_CO6),
.I2(CLBLM_L_X10Y154_SLICE_X13Y154_BQ),
.I3(CLBLM_R_X13Y149_SLICE_X18Y149_CQ),
.I4(CLBLM_L_X12Y151_SLICE_X17Y151_BQ),
.I5(CLBLM_R_X11Y151_SLICE_X14Y151_BQ),
.O5(CLBLM_R_X11Y151_SLICE_X15Y151_DO5),
.O6(CLBLM_R_X11Y151_SLICE_X15Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffe)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_CLUT (
.I0(CLBLM_L_X12Y152_SLICE_X16Y152_BQ),
.I1(CLBLM_R_X11Y150_SLICE_X14Y150_BO6),
.I2(CLBLM_L_X10Y158_SLICE_X13Y158_BQ),
.I3(CLBLM_R_X7Y149_SLICE_X8Y149_CQ),
.I4(CLBLM_L_X12Y151_SLICE_X17Y151_A5Q),
.I5(CLBLM_R_X11Y151_SLICE_X15Y151_DO6),
.O5(CLBLM_R_X11Y151_SLICE_X15Y151_CO5),
.O6(CLBLM_R_X11Y151_SLICE_X15Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ee00f0f0eeee)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_BLUT (
.I0(CLBLM_R_X11Y152_SLICE_X15Y152_DQ),
.I1(CLBLM_R_X11Y151_SLICE_X15Y151_BQ),
.I2(CLBLM_R_X13Y149_SLICE_X19Y149_CQ),
.I3(CLBLM_L_X12Y155_SLICE_X16Y155_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y150_SLICE_X12Y150_A5Q),
.O5(CLBLM_R_X11Y151_SLICE_X15Y151_BO5),
.O6(CLBLM_R_X11Y151_SLICE_X15Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcac0cac0afafa0a0)
  ) CLBLM_R_X11Y151_SLICE_X15Y151_ALUT (
.I0(CLBLM_L_X12Y151_SLICE_X17Y151_A5Q),
.I1(CLBLM_L_X10Y147_SLICE_X12Y147_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X8Y154_SLICE_X10Y154_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y151_SLICE_X15Y151_AO5),
.O6(CLBLM_R_X11Y151_SLICE_X15Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_B5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y152_SLICE_X14Y152_BO5),
.Q(CLBLM_R_X11Y152_SLICE_X14Y152_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y152_SLICE_X14Y152_AO6),
.Q(CLBLM_R_X11Y152_SLICE_X14Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y152_SLICE_X14Y152_BO6),
.Q(CLBLM_R_X11Y152_SLICE_X14Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y152_SLICE_X14Y152_CO6),
.Q(CLBLM_R_X11Y152_SLICE_X14Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaa0aaa0dddd8888)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_DLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_L_X10Y158_SLICE_X13Y158_BQ),
.I2(CLBLM_L_X8Y154_SLICE_X11Y154_CQ),
.I3(CLBLM_L_X10Y151_SLICE_X13Y151_BQ),
.I4(CLBLM_L_X12Y150_SLICE_X17Y150_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y152_SLICE_X14Y152_DO5),
.O6(CLBLM_R_X11Y152_SLICE_X14Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0ffc0cfa0af808)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_CLUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X11Y152_SLICE_X14Y152_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X8Y152_SLICE_X10Y152_BQ),
.I4(CLBLM_L_X10Y152_SLICE_X12Y152_CO6),
.I5(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.O5(CLBLM_R_X11Y152_SLICE_X14Y152_CO5),
.O6(CLBLM_R_X11Y152_SLICE_X14Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0aaf0aaffcc00cc)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_BLUT (
.I0(CLBLM_L_X12Y152_SLICE_X17Y152_A5Q),
.I1(CLBLM_L_X12Y152_SLICE_X16Y152_B5Q),
.I2(CLBLM_R_X11Y156_SLICE_X15Y156_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X5Y151_SLICE_X6Y151_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y152_SLICE_X14Y152_BO5),
.O6(CLBLM_R_X11Y152_SLICE_X14Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaa00aaffa000a0)
  ) CLBLM_R_X11Y152_SLICE_X14Y152_ALUT (
.I0(CLBLM_R_X7Y153_SLICE_X9Y153_CO6),
.I1(1'b1),
.I2(CLBLM_R_X11Y152_SLICE_X14Y152_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y150_SLICE_X13Y150_AQ),
.I5(CLBLM_L_X8Y153_SLICE_X11Y153_CQ),
.O5(CLBLM_R_X11Y152_SLICE_X14Y152_AO5),
.O6(CLBLM_R_X11Y152_SLICE_X14Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y152_SLICE_X15Y152_AO6),
.Q(CLBLM_R_X11Y152_SLICE_X15Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y152_SLICE_X15Y152_BO6),
.Q(CLBLM_R_X11Y152_SLICE_X15Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y152_SLICE_X15Y152_CO6),
.Q(CLBLM_R_X11Y152_SLICE_X15Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y152_SLICE_X15Y152_DO6),
.Q(CLBLM_R_X11Y152_SLICE_X15Y152_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff7800000078)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_DLUT (
.I0(CLBLM_L_X10Y152_SLICE_X13Y152_CO6),
.I1(CLBLM_L_X10Y148_SLICE_X13Y148_AQ),
.I2(CLBLM_R_X11Y152_SLICE_X15Y152_DQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y146_SLICE_X14Y146_AQ),
.I5(CLBLM_R_X7Y151_SLICE_X8Y151_DQ),
.O5(CLBLM_R_X11Y152_SLICE_X15Y152_DO5),
.O6(CLBLM_R_X11Y152_SLICE_X15Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffc000c0ffaa00aa)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_CLUT (
.I0(CLBLM_L_X12Y153_SLICE_X17Y153_BQ),
.I1(CLBLM_R_X11Y152_SLICE_X15Y152_CQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y154_SLICE_X14Y154_DQ),
.I5(CLBLM_R_X11Y149_SLICE_X15Y149_DO6),
.O5(CLBLM_R_X11Y152_SLICE_X15Y152_CO5),
.O6(CLBLM_R_X11Y152_SLICE_X15Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00d5d58080)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_BLUT (
.I0(CLBLM_R_X11Y149_SLICE_X15Y149_DO6),
.I1(CLBLM_R_X11Y152_SLICE_X15Y152_BQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X8Y152_SLICE_X10Y152_AQ),
.I4(CLBLM_R_X13Y153_SLICE_X18Y153_BQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y152_SLICE_X15Y152_BO5),
.O6(CLBLM_R_X11Y152_SLICE_X15Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0000ccc0)
  ) CLBLM_R_X11Y152_SLICE_X15Y152_ALUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_AQ),
.I1(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I2(CLBLM_R_X11Y152_SLICE_X15Y152_AQ),
.I3(CLBLM_R_X11Y153_SLICE_X14Y153_BO6),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y152_SLICE_X15Y152_AO5),
.O6(CLBLM_R_X11Y152_SLICE_X15Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y153_SLICE_X14Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y153_SLICE_X14Y153_AO6),
.Q(CLBLM_R_X11Y153_SLICE_X14Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffbfffb)
  ) CLBLM_R_X11Y153_SLICE_X14Y153_DLUT (
.I0(CLBLM_L_X10Y152_SLICE_X13Y152_AQ),
.I1(CLBLM_L_X10Y150_SLICE_X13Y150_BQ),
.I2(CLBLM_L_X12Y152_SLICE_X17Y152_BO5),
.I3(CLBLM_R_X11Y153_SLICE_X14Y153_CO6),
.I4(1'b1),
.I5(CLBLM_R_X5Y147_SLICE_X7Y147_BQ),
.O5(CLBLM_R_X11Y153_SLICE_X14Y153_DO5),
.O6(CLBLM_R_X11Y153_SLICE_X14Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffff7)
  ) CLBLM_R_X11Y153_SLICE_X14Y153_CLUT (
.I0(CLBLM_R_X13Y149_SLICE_X19Y149_AQ),
.I1(CLBLM_L_X8Y153_SLICE_X11Y153_BQ),
.I2(CLBLM_L_X12Y154_SLICE_X17Y154_A5Q),
.I3(CLBLL_L_X4Y151_SLICE_X4Y151_AQ),
.I4(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.I5(CLBLM_L_X8Y158_SLICE_X10Y158_BQ),
.O5(CLBLM_R_X11Y153_SLICE_X14Y153_CO5),
.O6(CLBLM_R_X11Y153_SLICE_X14Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaacc88a0a0cc80)
  ) CLBLM_R_X11Y153_SLICE_X14Y153_BLUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_L_X10Y149_SLICE_X13Y149_AQ),
.I2(CLBLM_L_X8Y154_SLICE_X11Y154_CQ),
.I3(CLBLM_R_X13Y152_SLICE_X18Y152_BO5),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_AQ),
.I5(CLBLM_L_X10Y151_SLICE_X13Y151_BQ),
.O5(CLBLM_R_X11Y153_SLICE_X14Y153_BO5),
.O6(CLBLM_R_X11Y153_SLICE_X14Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffc3330eeec2220)
  ) CLBLM_R_X11Y153_SLICE_X14Y153_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X11Y153_SLICE_X14Y153_AQ),
.I3(CLBLM_R_X11Y153_SLICE_X14Y153_BO6),
.I4(CLBLM_L_X10Y148_SLICE_X13Y148_AQ),
.I5(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.O5(CLBLM_R_X11Y153_SLICE_X14Y153_AO5),
.O6(CLBLM_R_X11Y153_SLICE_X14Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y153_SLICE_X15Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y153_SLICE_X15Y153_AO6),
.Q(CLBLM_R_X11Y153_SLICE_X15Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y153_SLICE_X15Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y153_SLICE_X15Y153_BO6),
.Q(CLBLM_R_X11Y153_SLICE_X15Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y153_SLICE_X15Y153_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y153_SLICE_X15Y153_CO6),
.Q(CLBLM_R_X11Y153_SLICE_X15Y153_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y153_SLICE_X15Y153_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y153_SLICE_X15Y153_DO6),
.Q(CLBLM_R_X11Y153_SLICE_X15Y153_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000fffa5550)
  ) CLBLM_R_X11Y153_SLICE_X15Y153_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(1'b1),
.I2(CLBLM_R_X11Y153_SLICE_X15Y153_DQ),
.I3(CLBLM_R_X13Y153_SLICE_X19Y153_CQ),
.I4(CLBLM_L_X8Y154_SLICE_X10Y154_DQ),
.I5(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.O5(CLBLM_R_X11Y153_SLICE_X15Y153_DO5),
.O6(CLBLM_R_X11Y153_SLICE_X15Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hefaf4505eaaa4000)
  ) CLBLM_R_X11Y153_SLICE_X15Y153_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y153_SLICE_X15Y153_CQ),
.I2(CLBLM_R_X11Y149_SLICE_X15Y149_DO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y152_SLICE_X13Y152_AQ),
.I5(CLBLM_R_X13Y153_SLICE_X19Y153_AQ),
.O5(CLBLM_R_X11Y153_SLICE_X15Y153_CO5),
.O6(CLBLM_R_X11Y153_SLICE_X15Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ccccf0f0aaaa)
  ) CLBLM_R_X11Y153_SLICE_X15Y153_BLUT (
.I0(CLBLM_L_X8Y155_SLICE_X11Y155_CQ),
.I1(CLBLM_R_X11Y153_SLICE_X15Y153_BQ),
.I2(CLBLM_R_X11Y153_SLICE_X15Y153_CQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y153_SLICE_X9Y153_CO6),
.O5(CLBLM_R_X11Y153_SLICE_X15Y153_BO5),
.O6(CLBLM_R_X11Y153_SLICE_X15Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffe0ff00ffe0)
  ) CLBLM_R_X11Y153_SLICE_X15Y153_ALUT (
.I0(RIOB33_X105Y117_IOB_X1Y118_I),
.I1(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I2(CLBLM_R_X11Y153_SLICE_X15Y153_AQ),
.I3(CLBLM_L_X10Y152_SLICE_X12Y152_DO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y153_SLICE_X15Y153_DQ),
.O5(CLBLM_R_X11Y153_SLICE_X15Y153_AO5),
.O6(CLBLM_R_X11Y153_SLICE_X15Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y154_SLICE_X14Y154_D5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y154_SLICE_X14Y154_DO5),
.Q(CLBLM_R_X11Y154_SLICE_X14Y154_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y154_SLICE_X14Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y154_SLICE_X14Y154_AO6),
.Q(CLBLM_R_X11Y154_SLICE_X14Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y154_SLICE_X14Y154_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y154_SLICE_X14Y154_CO6),
.Q(CLBLM_R_X11Y154_SLICE_X14Y154_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y154_SLICE_X14Y154_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y154_SLICE_X14Y154_DO6),
.Q(CLBLM_R_X11Y154_SLICE_X14Y154_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff55aa00d8d8d8d8)
  ) CLBLM_R_X11Y154_SLICE_X14Y154_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y154_SLICE_X14Y154_CQ),
.I2(CLBLM_L_X8Y159_SLICE_X10Y159_AQ),
.I3(CLBLM_R_X11Y148_SLICE_X14Y148_CQ),
.I4(CLBLM_L_X12Y157_SLICE_X17Y157_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y154_SLICE_X14Y154_DO5),
.O6(CLBLM_R_X11Y154_SLICE_X14Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h888d88d8888d88d8)
  ) CLBLM_R_X11Y154_SLICE_X14Y154_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y152_SLICE_X16Y152_AQ),
.I2(CLBLM_R_X13Y151_SLICE_X18Y151_CQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y154_SLICE_X14Y154_BO5),
.I5(1'b1),
.O5(CLBLM_R_X11Y154_SLICE_X14Y154_CO5),
.O6(CLBLM_R_X11Y154_SLICE_X14Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafaca0a0ffcc0000)
  ) CLBLM_R_X11Y154_SLICE_X14Y154_BLUT (
.I0(CLBLM_R_X13Y153_SLICE_X19Y153_CQ),
.I1(CLBLM_L_X10Y149_SLICE_X12Y149_C5Q),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y154_SLICE_X13Y154_DQ),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y154_SLICE_X14Y154_BO5),
.O6(CLBLM_R_X11Y154_SLICE_X14Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888ddd88888)
  ) CLBLM_R_X11Y154_SLICE_X14Y154_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y160_SLICE_X14Y160_AQ),
.I2(CLBLM_R_X11Y154_SLICE_X14Y154_AQ),
.I3(CLBLM_R_X7Y150_SLICE_X9Y150_BO6),
.I4(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X11Y154_SLICE_X14Y154_AO5),
.O6(CLBLM_R_X11Y154_SLICE_X14Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y154_SLICE_X15Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y154_SLICE_X15Y154_AO6),
.Q(CLBLM_R_X11Y154_SLICE_X15Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y154_SLICE_X15Y154_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y154_SLICE_X15Y154_BO6),
.Q(CLBLM_R_X11Y154_SLICE_X15Y154_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffd)
  ) CLBLM_R_X11Y154_SLICE_X15Y154_DLUT (
.I0(CLBLM_R_X11Y146_SLICE_X15Y146_AQ),
.I1(CLBLL_L_X4Y155_SLICE_X4Y155_CO6),
.I2(CLBLM_R_X11Y156_SLICE_X15Y156_DO6),
.I3(CLBLM_R_X11Y155_SLICE_X15Y155_CO6),
.I4(CLBLM_R_X13Y152_SLICE_X18Y152_BO5),
.I5(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.O5(CLBLM_R_X11Y154_SLICE_X15Y154_DO5),
.O6(CLBLM_R_X11Y154_SLICE_X15Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4e4a0cccccc00)
  ) CLBLM_R_X11Y154_SLICE_X15Y154_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_R_X11Y154_SLICE_X14Y154_D5Q),
.I3(CLBLM_L_X10Y155_SLICE_X13Y155_BQ),
.I4(CLBLM_R_X11Y151_SLICE_X15Y151_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y154_SLICE_X15Y154_CO5),
.O6(CLBLM_R_X11Y154_SLICE_X15Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f6f0f000060000)
  ) CLBLM_R_X11Y154_SLICE_X15Y154_BLUT (
.I0(CLBLM_L_X12Y154_SLICE_X16Y154_DO6),
.I1(CLBLM_R_X11Y154_SLICE_X15Y154_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y153_SLICE_X8Y153_AQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X8Y150_SLICE_X10Y150_BQ),
.O5(CLBLM_R_X11Y154_SLICE_X15Y154_BO5),
.O6(CLBLM_R_X11Y154_SLICE_X15Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccaaaacccca0a0)
  ) CLBLM_R_X11Y154_SLICE_X15Y154_ALUT (
.I0(CLBLM_R_X7Y153_SLICE_X9Y153_CO6),
.I1(CLBLM_R_X11Y155_SLICE_X15Y155_AQ),
.I2(CLBLM_R_X11Y154_SLICE_X15Y154_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X13Y151_SLICE_X18Y151_CQ),
.O5(CLBLM_R_X11Y154_SLICE_X15Y154_AO5),
.O6(CLBLM_R_X11Y154_SLICE_X15Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y155_SLICE_X14Y155_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y155_SLICE_X14Y155_AO6),
.Q(CLBLM_R_X11Y155_SLICE_X14Y155_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y155_SLICE_X14Y155_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y155_SLICE_X14Y155_BO6),
.Q(CLBLM_R_X11Y155_SLICE_X14Y155_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y155_SLICE_X14Y155_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y155_SLICE_X14Y155_CO6),
.Q(CLBLM_R_X11Y155_SLICE_X14Y155_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y155_SLICE_X14Y155_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y155_SLICE_X14Y155_DO6),
.Q(CLBLM_R_X11Y155_SLICE_X14Y155_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haafeaaaa00540000)
  ) CLBLM_R_X11Y155_SLICE_X14Y155_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y152_SLICE_X12Y152_CO6),
.I2(CLBLM_R_X11Y155_SLICE_X14Y155_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I5(CLBLM_L_X8Y155_SLICE_X11Y155_AQ),
.O5(CLBLM_R_X11Y155_SLICE_X14Y155_DO5),
.O6(CLBLM_R_X11Y155_SLICE_X14Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffaaf0aaffaaf0)
  ) CLBLM_R_X11Y155_SLICE_X14Y155_CLUT (
.I0(CLBLM_R_X7Y153_SLICE_X8Y153_AQ),
.I1(1'b1),
.I2(CLBLM_L_X10Y159_SLICE_X12Y159_CO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y156_SLICE_X14Y156_DO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y155_SLICE_X14Y155_CO5),
.O6(CLBLM_R_X11Y155_SLICE_X14Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafafa0a0afaca0ac)
  ) CLBLM_R_X11Y155_SLICE_X14Y155_BLUT (
.I0(CLBLM_L_X10Y154_SLICE_X13Y154_DQ),
.I1(CLBLM_R_X11Y155_SLICE_X14Y155_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I4(CLBLM_L_X12Y155_SLICE_X17Y155_BQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X11Y155_SLICE_X14Y155_BO5),
.O6(CLBLM_R_X11Y155_SLICE_X14Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00a8a8ff00a8a8)
  ) CLBLM_R_X11Y155_SLICE_X14Y155_ALUT (
.I0(CLBLM_R_X7Y153_SLICE_X9Y153_CO6),
.I1(CLBLM_R_X11Y154_SLICE_X14Y154_CQ),
.I2(CLBLM_R_X11Y155_SLICE_X14Y155_AQ),
.I3(CLBLM_R_X11Y152_SLICE_X15Y152_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y155_SLICE_X14Y155_AO5),
.O6(CLBLM_R_X11Y155_SLICE_X14Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y155_SLICE_X15Y155_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y155_SLICE_X15Y155_AO6),
.Q(CLBLM_R_X11Y155_SLICE_X15Y155_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefefefffefefefc)
  ) CLBLM_R_X11Y155_SLICE_X15Y155_DLUT (
.I0(CLBLM_L_X12Y155_SLICE_X17Y155_BQ),
.I1(CLBLM_L_X12Y153_SLICE_X16Y153_DO6),
.I2(CLBLM_L_X8Y157_SLICE_X11Y157_DO6),
.I3(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X11Y155_SLICE_X14Y155_BQ),
.O5(CLBLM_R_X11Y155_SLICE_X15Y155_DO5),
.O6(CLBLM_R_X11Y155_SLICE_X15Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffdfffffff)
  ) CLBLM_R_X11Y155_SLICE_X15Y155_CLUT (
.I0(CLBLM_R_X11Y157_SLICE_X15Y157_AQ),
.I1(CLBLM_R_X3Y157_SLICE_X2Y157_AO5),
.I2(CLBLM_L_X12Y155_SLICE_X16Y155_BO5),
.I3(CLBLM_L_X12Y155_SLICE_X16Y155_DO6),
.I4(CLBLM_R_X5Y149_SLICE_X7Y149_AQ),
.I5(CLBLM_R_X11Y155_SLICE_X15Y155_DO6),
.O5(CLBLM_R_X11Y155_SLICE_X15Y155_CO5),
.O6(CLBLM_R_X11Y155_SLICE_X15Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffffbf)
  ) CLBLM_R_X11Y155_SLICE_X15Y155_BLUT (
.I0(CLBLM_R_X11Y156_SLICE_X14Y156_DO6),
.I1(CLBLM_R_X7Y149_SLICE_X8Y149_DO5),
.I2(CLBLM_L_X8Y155_SLICE_X10Y155_DO6),
.I3(CLBLM_L_X12Y156_SLICE_X16Y156_DO6),
.I4(CLBLM_R_X13Y156_SLICE_X18Y156_BO6),
.I5(CLBLM_L_X10Y159_SLICE_X12Y159_CO6),
.O5(CLBLM_R_X11Y155_SLICE_X15Y155_BO5),
.O6(CLBLM_R_X11Y155_SLICE_X15Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccafafccccfafa)
  ) CLBLM_R_X11Y155_SLICE_X15Y155_ALUT (
.I0(CLBLM_R_X11Y158_SLICE_X15Y158_BO6),
.I1(CLBLM_R_X5Y150_SLICE_X6Y150_DQ),
.I2(CLBLM_R_X11Y155_SLICE_X15Y155_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y155_SLICE_X16Y155_BO6),
.O5(CLBLM_R_X11Y155_SLICE_X15Y155_AO5),
.O6(CLBLM_R_X11Y155_SLICE_X15Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y156_SLICE_X14Y156_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y156_SLICE_X14Y156_AO6),
.Q(CLBLM_R_X11Y156_SLICE_X14Y156_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y156_SLICE_X14Y156_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y156_SLICE_X14Y156_BO6),
.Q(CLBLM_R_X11Y156_SLICE_X14Y156_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc300c300c300c300)
  ) CLBLM_R_X11Y156_SLICE_X14Y156_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y155_SLICE_X14Y155_CQ),
.I2(CLBLM_L_X10Y157_SLICE_X12Y157_DO6),
.I3(CLBLM_L_X10Y159_SLICE_X12Y159_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y156_SLICE_X14Y156_DO5),
.O6(CLBLM_R_X11Y156_SLICE_X14Y156_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000dffeffff)
  ) CLBLM_R_X11Y156_SLICE_X14Y156_CLUT (
.I0(CLBLM_R_X11Y156_SLICE_X15Y156_AQ),
.I1(CLBLM_L_X8Y156_SLICE_X11Y156_DO6),
.I2(CLBLM_L_X10Y157_SLICE_X13Y157_AO5),
.I3(CLBLM_L_X12Y157_SLICE_X16Y157_CQ),
.I4(CLBLM_R_X7Y157_SLICE_X9Y157_AQ),
.I5(CLBLM_L_X8Y157_SLICE_X11Y157_DO6),
.O5(CLBLM_R_X11Y156_SLICE_X14Y156_CO5),
.O6(CLBLM_R_X11Y156_SLICE_X14Y156_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfc0d0cfdfc0d0c)
  ) CLBLM_R_X11Y156_SLICE_X14Y156_BLUT (
.I0(CLBLM_L_X10Y157_SLICE_X13Y157_CO6),
.I1(CLBLM_L_X10Y159_SLICE_X12Y159_CO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y159_SLICE_X12Y159_DO6),
.I4(CLBLM_R_X11Y152_SLICE_X15Y152_DQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y156_SLICE_X14Y156_BO5),
.O6(CLBLM_R_X11Y156_SLICE_X14Y156_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff007575ff002020)
  ) CLBLM_R_X11Y156_SLICE_X14Y156_ALUT (
.I0(CLBLM_R_X11Y159_SLICE_X15Y159_DO5),
.I1(CLBLM_R_X11Y158_SLICE_X15Y158_BO6),
.I2(CLBLM_R_X11Y156_SLICE_X14Y156_AQ),
.I3(CLBLM_R_X3Y150_SLICE_X3Y150_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y157_SLICE_X16Y157_BQ),
.O5(CLBLM_R_X11Y156_SLICE_X14Y156_AO5),
.O6(CLBLM_R_X11Y156_SLICE_X14Y156_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y156_SLICE_X15Y156_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y156_SLICE_X15Y156_AO6),
.Q(CLBLM_R_X11Y156_SLICE_X15Y156_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y156_SLICE_X15Y156_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y156_SLICE_X15Y156_BO6),
.Q(CLBLM_R_X11Y156_SLICE_X15Y156_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00eeffff00ee)
  ) CLBLM_R_X11Y156_SLICE_X15Y156_DLUT (
.I0(CLBLM_L_X10Y158_SLICE_X13Y158_AQ),
.I1(CLBLM_R_X11Y157_SLICE_X14Y157_CQ),
.I2(1'b1),
.I3(CLBLM_R_X11Y159_SLICE_X15Y159_DO5),
.I4(CLBLM_R_X11Y158_SLICE_X15Y158_BO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y156_SLICE_X15Y156_DO5),
.O6(CLBLM_R_X11Y156_SLICE_X15Y156_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfdf5f5f7f7f5f5f)
  ) CLBLM_R_X11Y156_SLICE_X15Y156_CLUT (
.I0(CLBLM_R_X11Y158_SLICE_X15Y158_DO6),
.I1(CLBLM_R_X11Y156_SLICE_X14Y156_CO6),
.I2(CLBLM_R_X11Y150_SLICE_X15Y150_BO6),
.I3(1'b1),
.I4(CLBLM_L_X10Y159_SLICE_X12Y159_DO6),
.I5(CLBLM_L_X10Y157_SLICE_X12Y157_BQ),
.O5(CLBLM_R_X11Y156_SLICE_X15Y156_CO5),
.O6(CLBLM_R_X11Y156_SLICE_X15Y156_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cff0ffc0cfc0c)
  ) CLBLM_R_X11Y156_SLICE_X15Y156_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y156_SLICE_X15Y156_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y159_SLICE_X15Y159_BQ),
.I4(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.I5(RIOB33_X105Y141_IOB_X1Y142_I),
.O5(CLBLM_R_X11Y156_SLICE_X15Y156_BO5),
.O6(CLBLM_R_X11Y156_SLICE_X15Y156_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffff820000ff82)
  ) CLBLM_R_X11Y156_SLICE_X15Y156_ALUT (
.I0(CLBLM_L_X10Y159_SLICE_X12Y159_DO6),
.I1(CLBLM_R_X11Y157_SLICE_X15Y157_CO6),
.I2(CLBLM_R_X11Y156_SLICE_X15Y156_AQ),
.I3(CLBLM_L_X10Y159_SLICE_X12Y159_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLL_L_X4Y149_SLICE_X5Y149_AQ),
.O5(CLBLM_R_X11Y156_SLICE_X15Y156_AO5),
.O6(CLBLM_R_X11Y156_SLICE_X15Y156_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y157_SLICE_X14Y157_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y157_SLICE_X14Y157_AO6),
.Q(CLBLM_R_X11Y157_SLICE_X14Y157_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y157_SLICE_X14Y157_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y157_SLICE_X14Y157_BO6),
.Q(CLBLM_R_X11Y157_SLICE_X14Y157_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y157_SLICE_X14Y157_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y157_SLICE_X14Y157_CO6),
.Q(CLBLM_R_X11Y157_SLICE_X14Y157_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffcfe)
  ) CLBLM_R_X11Y157_SLICE_X14Y157_DLUT (
.I0(CLBLM_L_X10Y159_SLICE_X12Y159_DO6),
.I1(CLBLM_L_X10Y155_SLICE_X13Y155_CO6),
.I2(CLBLM_R_X3Y153_SLICE_X3Y153_BO6),
.I3(CLBLM_L_X10Y159_SLICE_X13Y159_CO6),
.I4(CLBLM_L_X12Y157_SLICE_X17Y157_DO6),
.I5(CLBLM_L_X10Y159_SLICE_X12Y159_CO6),
.O5(CLBLM_R_X11Y157_SLICE_X14Y157_DO5),
.O6(CLBLM_R_X11Y157_SLICE_X14Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00f0aaaaccf0)
  ) CLBLM_R_X11Y157_SLICE_X14Y157_CLUT (
.I0(CLBLM_R_X7Y157_SLICE_X9Y157_AQ),
.I1(CLBLM_R_X11Y157_SLICE_X14Y157_CQ),
.I2(CLBLM_R_X11Y157_SLICE_X14Y157_BQ),
.I3(CLBLM_R_X11Y159_SLICE_X15Y159_DO5),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y158_SLICE_X15Y158_BO6),
.O5(CLBLM_R_X11Y157_SLICE_X14Y157_CO5),
.O6(CLBLM_R_X11Y157_SLICE_X14Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc5cfc0cac5c5c0c0)
  ) CLBLM_R_X11Y157_SLICE_X14Y157_BLUT (
.I0(CLBLM_R_X11Y159_SLICE_X15Y159_DO5),
.I1(CLBLL_L_X4Y152_SLICE_X5Y152_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y158_SLICE_X15Y158_BO6),
.I4(CLBLM_R_X11Y158_SLICE_X14Y158_BQ),
.I5(CLBLM_R_X11Y157_SLICE_X14Y157_BQ),
.O5(CLBLM_R_X11Y157_SLICE_X14Y157_BO5),
.O6(CLBLM_R_X11Y157_SLICE_X14Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ff000ff0f90009)
  ) CLBLM_R_X11Y157_SLICE_X14Y157_ALUT (
.I0(CLBLM_L_X12Y157_SLICE_X17Y157_DO6),
.I1(CLBLM_R_X11Y157_SLICE_X14Y157_AQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y159_SLICE_X15Y159_CO5),
.I4(CLBLM_L_X8Y157_SLICE_X11Y157_BQ),
.I5(CLBLM_R_X11Y158_SLICE_X14Y158_DO5),
.O5(CLBLM_R_X11Y157_SLICE_X14Y157_AO5),
.O6(CLBLM_R_X11Y157_SLICE_X14Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y157_SLICE_X15Y157_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y157_SLICE_X15Y157_AO6),
.Q(CLBLM_R_X11Y157_SLICE_X15Y157_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y157_SLICE_X15Y157_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y157_SLICE_X15Y157_BO6),
.Q(CLBLM_R_X11Y157_SLICE_X15Y157_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2200222288aa8888)
  ) CLBLM_R_X11Y157_SLICE_X15Y157_DLUT (
.I0(CLBLM_L_X10Y159_SLICE_X12Y159_DO6),
.I1(CLBLM_L_X8Y157_SLICE_X11Y157_DO6),
.I2(1'b1),
.I3(CLBLM_L_X8Y156_SLICE_X11Y156_DO6),
.I4(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.I5(CLBLM_L_X12Y157_SLICE_X16Y157_CQ),
.O5(CLBLM_R_X11Y157_SLICE_X15Y157_DO5),
.O6(CLBLM_R_X11Y157_SLICE_X15Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00be00be00ff00ff)
  ) CLBLM_R_X11Y157_SLICE_X15Y157_CLUT (
.I0(CLBLM_L_X8Y156_SLICE_X11Y156_DO6),
.I1(CLBLM_L_X12Y157_SLICE_X16Y157_CQ),
.I2(CLBLM_L_X10Y157_SLICE_X13Y157_AO5),
.I3(CLBLM_L_X8Y157_SLICE_X11Y157_DO6),
.I4(1'b1),
.I5(CLBLM_R_X7Y155_SLICE_X9Y155_BQ),
.O5(CLBLM_R_X11Y157_SLICE_X15Y157_CO5),
.O6(CLBLM_R_X11Y157_SLICE_X15Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaf3f3aaaaf0f0)
  ) CLBLM_R_X11Y157_SLICE_X15Y157_BLUT (
.I0(CLBLM_L_X8Y149_SLICE_X11Y149_CQ),
.I1(CLBLM_R_X11Y159_SLICE_X15Y159_CO5),
.I2(CLBLM_L_X12Y156_SLICE_X16Y156_DO6),
.I3(1'b1),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y158_SLICE_X14Y158_DO5),
.O5(CLBLM_R_X11Y157_SLICE_X15Y157_BO5),
.O6(CLBLM_R_X11Y157_SLICE_X15Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff000303ff003232)
  ) CLBLM_R_X11Y157_SLICE_X15Y157_ALUT (
.I0(CLBLM_R_X11Y158_SLICE_X15Y158_BO5),
.I1(RIOB33_X105Y121_IOB_X1Y121_I),
.I2(CLBLM_R_X11Y157_SLICE_X15Y157_AQ),
.I3(CLBLM_L_X10Y155_SLICE_X13Y155_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y157_SLICE_X16Y157_DO6),
.O5(CLBLM_R_X11Y157_SLICE_X15Y157_AO5),
.O6(CLBLM_R_X11Y157_SLICE_X15Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y158_SLICE_X14Y158_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y158_SLICE_X14Y158_AO6),
.Q(CLBLM_R_X11Y158_SLICE_X14Y158_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y158_SLICE_X14Y158_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y158_SLICE_X14Y158_BO6),
.Q(CLBLM_R_X11Y158_SLICE_X14Y158_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y158_SLICE_X14Y158_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y158_SLICE_X14Y158_CO6),
.Q(CLBLM_R_X11Y158_SLICE_X14Y158_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h40404043bfb000bc)
  ) CLBLM_R_X11Y158_SLICE_X14Y158_DLUT (
.I0(CLBLM_R_X11Y157_SLICE_X15Y157_AQ),
.I1(CLBLM_R_X11Y159_SLICE_X14Y159_BQ),
.I2(CLBLM_L_X12Y158_SLICE_X16Y158_AQ),
.I3(CLBLM_R_X11Y159_SLICE_X15Y159_AQ),
.I4(CLBLM_L_X12Y158_SLICE_X17Y158_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y158_SLICE_X14Y158_DO5),
.O6(CLBLM_R_X11Y158_SLICE_X14Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heaeaeaea44444440)
  ) CLBLM_R_X11Y158_SLICE_X14Y158_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y154_SLICE_X12Y154_CQ),
.I2(CLBLM_L_X12Y158_SLICE_X16Y158_AQ),
.I3(CLBLM_R_X11Y159_SLICE_X15Y159_AQ),
.I4(CLBLM_L_X12Y158_SLICE_X17Y158_AQ),
.I5(CLBLM_R_X11Y159_SLICE_X14Y159_BQ),
.O5(CLBLM_R_X11Y158_SLICE_X14Y158_CO5),
.O6(CLBLM_R_X11Y158_SLICE_X14Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff72ff5000720050)
  ) CLBLM_R_X11Y158_SLICE_X14Y158_BLUT (
.I0(CLBLM_R_X11Y159_SLICE_X15Y159_DO5),
.I1(CLBLM_R_X11Y158_SLICE_X15Y158_BO6),
.I2(CLBLM_R_X11Y156_SLICE_X14Y156_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y158_SLICE_X14Y158_BQ),
.I5(CLBLM_R_X7Y154_SLICE_X9Y154_CQ),
.O5(CLBLM_R_X11Y158_SLICE_X14Y158_BO5),
.O6(CLBLM_R_X11Y158_SLICE_X14Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000cfcccfcc)
  ) CLBLM_R_X11Y158_SLICE_X14Y158_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y156_SLICE_X18Y156_BO6),
.I2(CLBLM_R_X11Y159_SLICE_X15Y159_CO5),
.I3(CLBLM_R_X11Y158_SLICE_X14Y158_DO5),
.I4(CLBLM_R_X7Y158_SLICE_X8Y158_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X11Y158_SLICE_X14Y158_AO5),
.O6(CLBLM_R_X11Y158_SLICE_X14Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y158_SLICE_X15Y158_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y158_SLICE_X15Y158_AO6),
.Q(CLBLM_R_X11Y158_SLICE_X15Y158_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5554ffff5555ffff)
  ) CLBLM_R_X11Y158_SLICE_X15Y158_DLUT (
.I0(CLBLM_R_X11Y157_SLICE_X15Y157_AQ),
.I1(CLBLM_R_X11Y159_SLICE_X15Y159_AQ),
.I2(CLBLM_L_X12Y158_SLICE_X17Y158_AQ),
.I3(CLBLM_R_X11Y159_SLICE_X14Y159_BQ),
.I4(CLBLM_L_X12Y155_SLICE_X16Y155_BO5),
.I5(CLBLM_L_X12Y158_SLICE_X16Y158_AQ),
.O5(CLBLM_R_X11Y158_SLICE_X15Y158_DO5),
.O6(CLBLM_R_X11Y158_SLICE_X15Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fff3f0f2fff3f)
  ) CLBLM_R_X11Y158_SLICE_X15Y158_CLUT (
.I0(CLBLM_R_X11Y157_SLICE_X15Y157_AQ),
.I1(CLBLM_R_X11Y159_SLICE_X15Y159_AQ),
.I2(CLBLM_L_X8Y157_SLICE_X10Y157_DQ),
.I3(CLBLM_R_X11Y159_SLICE_X14Y159_BQ),
.I4(CLBLM_L_X12Y158_SLICE_X16Y158_AQ),
.I5(CLBLM_L_X12Y158_SLICE_X17Y158_AQ),
.O5(CLBLM_R_X11Y158_SLICE_X15Y158_CO5),
.O6(CLBLM_R_X11Y158_SLICE_X15Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001100100000)
  ) CLBLM_R_X11Y158_SLICE_X15Y158_BLUT (
.I0(CLBLM_R_X11Y159_SLICE_X14Y159_BQ),
.I1(CLBLM_R_X11Y159_SLICE_X15Y159_AQ),
.I2(CLBLM_L_X12Y155_SLICE_X16Y155_BO5),
.I3(CLBLM_L_X12Y158_SLICE_X17Y158_AQ),
.I4(CLBLM_L_X12Y158_SLICE_X16Y158_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y158_SLICE_X15Y158_BO5),
.O6(CLBLM_R_X11Y158_SLICE_X15Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa00f0aaaacccc)
  ) CLBLM_R_X11Y158_SLICE_X15Y158_ALUT (
.I0(CLBLM_L_X12Y152_SLICE_X17Y152_AQ),
.I1(CLBLM_L_X10Y158_SLICE_X13Y158_AQ),
.I2(CLBLM_R_X11Y158_SLICE_X15Y158_AQ),
.I3(CLBLM_R_X11Y158_SLICE_X15Y158_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X11Y159_SLICE_X15Y159_DO5),
.O5(CLBLM_R_X11Y158_SLICE_X15Y158_AO5),
.O6(CLBLM_R_X11Y158_SLICE_X15Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y159_SLICE_X14Y159_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y159_SLICE_X14Y159_AO6),
.Q(CLBLM_R_X11Y159_SLICE_X14Y159_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y159_SLICE_X14Y159_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y159_SLICE_X14Y159_BO6),
.Q(CLBLM_R_X11Y159_SLICE_X14Y159_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y159_SLICE_X14Y159_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y159_SLICE_X14Y159_CO6),
.Q(CLBLM_R_X11Y159_SLICE_X14Y159_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y159_SLICE_X14Y159_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y159_SLICE_X14Y159_DO6),
.Q(CLBLM_R_X11Y159_SLICE_X14Y159_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc30fc30fe32fe32)
  ) CLBLM_R_X11Y159_SLICE_X14Y159_DLUT (
.I0(CLBLM_L_X10Y159_SLICE_X12Y159_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_L_X10Y159_SLICE_X12Y159_CO6),
.I3(CLBLM_L_X12Y152_SLICE_X17Y152_A5Q),
.I4(1'b1),
.I5(CLBLM_L_X8Y159_SLICE_X11Y159_AO6),
.O5(CLBLM_R_X11Y159_SLICE_X14Y159_DO5),
.O6(CLBLM_R_X11Y159_SLICE_X14Y159_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0f00aaaa0f03)
  ) CLBLM_R_X11Y159_SLICE_X14Y159_CLUT (
.I0(CLBLM_R_X11Y157_SLICE_X15Y157_AQ),
.I1(CLBLM_R_X11Y159_SLICE_X15Y159_AQ),
.I2(CLBLM_L_X12Y158_SLICE_X16Y158_AQ),
.I3(CLBLM_R_X11Y159_SLICE_X14Y159_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X12Y158_SLICE_X17Y158_AQ),
.O5(CLBLM_R_X11Y159_SLICE_X14Y159_CO5),
.O6(CLBLM_R_X11Y159_SLICE_X14Y159_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaafeb00000541)
  ) CLBLM_R_X11Y159_SLICE_X14Y159_BLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X11Y159_SLICE_X15Y159_DO6),
.I2(CLBLM_R_X11Y159_SLICE_X14Y159_BQ),
.I3(CLBLM_L_X12Y159_SLICE_X16Y159_BO6),
.I4(RIOB33_X105Y121_IOB_X1Y121_I),
.I5(CLBLM_L_X8Y155_SLICE_X10Y155_CQ),
.O5(CLBLM_R_X11Y159_SLICE_X14Y159_BO5),
.O6(CLBLM_R_X11Y159_SLICE_X14Y159_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hddddddddd8dd8888)
  ) CLBLM_R_X11Y159_SLICE_X14Y159_ALUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X8Y158_SLICE_X11Y158_BQ),
.I2(CLBLM_R_X11Y159_SLICE_X15Y159_CO5),
.I3(CLBLM_R_X11Y158_SLICE_X14Y158_DO6),
.I4(CLBLM_R_X11Y159_SLICE_X14Y159_AQ),
.I5(CLBLM_L_X12Y159_SLICE_X16Y159_BO6),
.O5(CLBLM_R_X11Y159_SLICE_X14Y159_AO5),
.O6(CLBLM_R_X11Y159_SLICE_X14Y159_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y159_SLICE_X15Y159_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y159_SLICE_X15Y159_AO6),
.Q(CLBLM_R_X11Y159_SLICE_X15Y159_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y159_SLICE_X15Y159_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y159_SLICE_X15Y159_BO6),
.Q(CLBLM_R_X11Y159_SLICE_X15Y159_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f1f3f3f40404040)
  ) CLBLM_R_X11Y159_SLICE_X15Y159_DLUT (
.I0(CLBLM_R_X11Y159_SLICE_X14Y159_BQ),
.I1(CLBLM_R_X11Y157_SLICE_X15Y157_AQ),
.I2(CLBLM_L_X12Y155_SLICE_X16Y155_BO5),
.I3(CLBLM_L_X12Y159_SLICE_X17Y159_AO5),
.I4(CLBLM_L_X12Y158_SLICE_X16Y158_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y159_SLICE_X15Y159_DO5),
.O6(CLBLM_R_X11Y159_SLICE_X15Y159_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00cc00dd0f0f0f0e)
  ) CLBLM_R_X11Y159_SLICE_X15Y159_CLUT (
.I0(CLBLM_L_X12Y158_SLICE_X17Y158_AQ),
.I1(CLBLM_R_X11Y159_SLICE_X14Y159_BQ),
.I2(CLBLM_L_X12Y159_SLICE_X17Y159_AO5),
.I3(CLBLM_L_X12Y158_SLICE_X16Y158_AQ),
.I4(CLBLM_R_X11Y159_SLICE_X15Y159_AQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y159_SLICE_X15Y159_CO5),
.O6(CLBLM_R_X11Y159_SLICE_X15Y159_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hafacafa0afa3afa0)
  ) CLBLM_R_X11Y159_SLICE_X15Y159_BLUT (
.I0(CLBLM_L_X12Y150_SLICE_X16Y150_AQ),
.I1(CLBLM_R_X11Y159_SLICE_X15Y159_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y159_SLICE_X12Y159_CO6),
.I4(CLBLM_L_X10Y159_SLICE_X12Y159_DO6),
.I5(CLBLM_L_X10Y159_SLICE_X13Y159_DO6),
.O5(CLBLM_R_X11Y159_SLICE_X15Y159_BO5),
.O6(CLBLM_R_X11Y159_SLICE_X15Y159_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00e2000000e2)
  ) CLBLM_R_X11Y159_SLICE_X15Y159_ALUT (
.I0(CLBLM_R_X11Y159_SLICE_X15Y159_AQ),
.I1(CLBLM_L_X12Y159_SLICE_X17Y159_AO6),
.I2(CLBLM_L_X12Y158_SLICE_X17Y158_AQ),
.I3(RIOB33_X105Y121_IOB_X1Y121_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X7Y153_SLICE_X8Y153_A5Q),
.O5(CLBLM_R_X11Y159_SLICE_X15Y159_AO5),
.O6(CLBLM_R_X11Y159_SLICE_X15Y159_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y160_SLICE_X14Y160_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X11Y160_SLICE_X14Y160_AO6),
.Q(CLBLM_R_X11Y160_SLICE_X14Y160_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y160_SLICE_X14Y160_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y160_SLICE_X14Y160_DO5),
.O6(CLBLM_R_X11Y160_SLICE_X14Y160_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y160_SLICE_X14Y160_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y160_SLICE_X14Y160_CO5),
.O6(CLBLM_R_X11Y160_SLICE_X14Y160_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y160_SLICE_X14Y160_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y160_SLICE_X14Y160_BO5),
.O6(CLBLM_R_X11Y160_SLICE_X14Y160_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffcfc0f0f0c0c)
  ) CLBLM_R_X11Y160_SLICE_X14Y160_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X10Y158_SLICE_X13Y158_CO6),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(1'b1),
.I4(CLBLM_L_X10Y159_SLICE_X12Y159_CO6),
.I5(CLBLM_R_X11Y159_SLICE_X14Y159_AQ),
.O5(CLBLM_R_X11Y160_SLICE_X14Y160_AO5),
.O6(CLBLM_R_X11Y160_SLICE_X14Y160_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y160_SLICE_X15Y160_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y160_SLICE_X15Y160_DO5),
.O6(CLBLM_R_X11Y160_SLICE_X15Y160_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y160_SLICE_X15Y160_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y160_SLICE_X15Y160_CO5),
.O6(CLBLM_R_X11Y160_SLICE_X15Y160_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y160_SLICE_X15Y160_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y160_SLICE_X15Y160_BO5),
.O6(CLBLM_R_X11Y160_SLICE_X15Y160_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y160_SLICE_X15Y160_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y160_SLICE_X15Y160_AO5),
.O6(CLBLM_R_X11Y160_SLICE_X15Y160_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1e1e0f0f0f0f0f0f)
  ) CLBLM_R_X13Y147_SLICE_X18Y147_DLUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_BQ),
.I1(CLBLM_L_X10Y145_SLICE_X13Y145_CQ),
.I2(CLBLM_R_X13Y153_SLICE_X19Y153_CQ),
.I3(1'b1),
.I4(CLBLM_L_X10Y146_SLICE_X12Y146_C5Q),
.I5(CLBLM_L_X10Y146_SLICE_X12Y146_CQ),
.O5(CLBLM_R_X13Y147_SLICE_X18Y147_DO5),
.O6(CLBLM_R_X13Y147_SLICE_X18Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f001f11ffffdfdd)
  ) CLBLM_R_X13Y147_SLICE_X18Y147_CLUT (
.I0(CLBLM_R_X13Y148_SLICE_X18Y148_BO5),
.I1(CLBLM_R_X5Y155_SLICE_X6Y155_DO6),
.I2(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(CLBLM_R_X13Y155_SLICE_X19Y155_AO6),
.I5(CLBLM_L_X12Y147_SLICE_X17Y147_AO6),
.O5(CLBLM_R_X13Y147_SLICE_X18Y147_CO5),
.O6(CLBLM_R_X13Y147_SLICE_X18Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1000efff0a0a0a0a)
  ) CLBLM_R_X13Y147_SLICE_X18Y147_BLUT (
.I0(CLBLM_L_X10Y146_SLICE_X12Y146_C5Q),
.I1(CLBLM_L_X10Y145_SLICE_X13Y145_CQ),
.I2(CLBLM_L_X10Y145_SLICE_X13Y145_BQ),
.I3(CLBLM_L_X10Y146_SLICE_X12Y146_CQ),
.I4(CLBLM_L_X12Y146_SLICE_X16Y146_DQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y147_SLICE_X18Y147_BO5),
.O6(CLBLM_R_X13Y147_SLICE_X18Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff02fdccccffff)
  ) CLBLM_R_X13Y147_SLICE_X18Y147_ALUT (
.I0(CLBLM_L_X10Y146_SLICE_X12Y146_C5Q),
.I1(CLBLM_L_X10Y146_SLICE_X12Y146_CQ),
.I2(CLBLM_L_X10Y145_SLICE_X13Y145_BQ),
.I3(CLBLM_L_X10Y145_SLICE_X12Y145_CQ),
.I4(CLBLM_L_X10Y145_SLICE_X13Y145_CQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y147_SLICE_X18Y147_AO5),
.O6(CLBLM_R_X13Y147_SLICE_X18Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y147_SLICE_X19Y147_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y147_SLICE_X19Y147_DO5),
.O6(CLBLM_R_X13Y147_SLICE_X19Y147_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y147_SLICE_X19Y147_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y147_SLICE_X19Y147_CO5),
.O6(CLBLM_R_X13Y147_SLICE_X19Y147_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y147_SLICE_X19Y147_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y147_SLICE_X19Y147_BO5),
.O6(CLBLM_R_X13Y147_SLICE_X19Y147_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y147_SLICE_X19Y147_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y147_SLICE_X19Y147_AO5),
.O6(CLBLM_R_X13Y147_SLICE_X19Y147_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y148_SLICE_X18Y148_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y148_SLICE_X18Y148_AO6),
.Q(CLBLM_R_X13Y148_SLICE_X18Y148_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y148_SLICE_X18Y148_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y148_SLICE_X18Y148_DO5),
.O6(CLBLM_R_X13Y148_SLICE_X18Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033003300331023)
  ) CLBLM_R_X13Y148_SLICE_X18Y148_CLUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_BQ),
.I1(CLBLM_R_X13Y153_SLICE_X18Y153_CQ),
.I2(CLBLM_L_X10Y145_SLICE_X13Y145_CQ),
.I3(CLBLM_L_X12Y148_SLICE_X16Y148_DO6),
.I4(CLBLM_L_X10Y146_SLICE_X12Y146_C5Q),
.I5(CLBLM_L_X10Y146_SLICE_X12Y146_CQ),
.O5(CLBLM_R_X13Y148_SLICE_X18Y148_CO5),
.O6(CLBLM_R_X13Y148_SLICE_X18Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a080dffffff00)
  ) CLBLM_R_X13Y148_SLICE_X18Y148_BLUT (
.I0(CLBLM_L_X12Y147_SLICE_X17Y147_AO6),
.I1(CLBLM_R_X7Y146_SLICE_X8Y146_DO6),
.I2(CLBLM_R_X13Y148_SLICE_X18Y148_AQ),
.I3(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.I4(CLBLM_R_X13Y148_SLICE_X18Y148_CO6),
.I5(1'b1),
.O5(CLBLM_R_X13Y148_SLICE_X18Y148_BO5),
.O6(CLBLM_R_X13Y148_SLICE_X18Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccc00af50505050)
  ) CLBLM_R_X13Y148_SLICE_X18Y148_ALUT (
.I0(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.I1(CLBLM_R_X13Y153_SLICE_X18Y153_CQ),
.I2(RIOB33_X105Y141_IOB_X1Y142_I),
.I3(CLBLM_R_X13Y148_SLICE_X18Y148_BO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X13Y148_SLICE_X18Y148_AO5),
.O6(CLBLM_R_X13Y148_SLICE_X18Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y148_SLICE_X19Y148_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y148_SLICE_X19Y148_DO5),
.O6(CLBLM_R_X13Y148_SLICE_X19Y148_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y148_SLICE_X19Y148_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y148_SLICE_X19Y148_CO5),
.O6(CLBLM_R_X13Y148_SLICE_X19Y148_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y148_SLICE_X19Y148_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y148_SLICE_X19Y148_BO5),
.O6(CLBLM_R_X13Y148_SLICE_X19Y148_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y148_SLICE_X19Y148_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y148_SLICE_X19Y148_AO5),
.O6(CLBLM_R_X13Y148_SLICE_X19Y148_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y149_SLICE_X18Y149_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y149_SLICE_X19Y149_BO6),
.Q(CLBLM_R_X13Y149_SLICE_X18Y149_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y149_SLICE_X18Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y149_SLICE_X18Y149_AO6),
.Q(CLBLM_R_X13Y149_SLICE_X18Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y149_SLICE_X18Y149_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y149_SLICE_X18Y149_BO6),
.Q(CLBLM_R_X13Y149_SLICE_X18Y149_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y149_SLICE_X18Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y149_SLICE_X18Y149_CO6),
.Q(CLBLM_R_X13Y149_SLICE_X18Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5500550555005504)
  ) CLBLM_R_X13Y149_SLICE_X18Y149_DLUT (
.I0(CLBLM_L_X12Y148_SLICE_X17Y148_AO6),
.I1(CLBLM_R_X5Y155_SLICE_X6Y155_BO6),
.I2(CLBLM_R_X13Y149_SLICE_X19Y149_DO6),
.I3(CLBLM_L_X12Y149_SLICE_X17Y149_DO6),
.I4(CLBLM_L_X12Y156_SLICE_X16Y156_AO6),
.I5(CLBLM_L_X12Y147_SLICE_X17Y147_AO6),
.O5(CLBLM_R_X13Y149_SLICE_X18Y149_DO5),
.O6(CLBLM_R_X13Y149_SLICE_X18Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa30aa30aa30aa30)
  ) CLBLM_R_X13Y149_SLICE_X18Y149_CLUT (
.I0(CLBLM_L_X10Y145_SLICE_X13Y145_BQ),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(CLBLM_L_X12Y151_SLICE_X17Y151_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y149_SLICE_X18Y149_CO5),
.O6(CLBLM_R_X13Y149_SLICE_X18Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa0000ffcc)
  ) CLBLM_R_X13Y149_SLICE_X18Y149_BLUT (
.I0(CLBLM_L_X10Y153_SLICE_X12Y153_AQ),
.I1(CLBLM_R_X13Y149_SLICE_X18Y149_BQ),
.I2(1'b1),
.I3(CLBLM_L_X12Y149_SLICE_X17Y149_AQ),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_DO6),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y149_SLICE_X18Y149_BO5),
.O6(CLBLM_R_X13Y149_SLICE_X18Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00fffc000000fc)
  ) CLBLM_R_X13Y149_SLICE_X18Y149_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y149_SLICE_X18Y149_BQ),
.I2(CLBLM_R_X13Y149_SLICE_X18Y149_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X7Y146_SLICE_X8Y146_DO6),
.I5(CLBLM_R_X13Y151_SLICE_X18Y151_CQ),
.O5(CLBLM_R_X13Y149_SLICE_X18Y149_AO5),
.O6(CLBLM_R_X13Y149_SLICE_X18Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y149_SLICE_X19Y149_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y149_SLICE_X19Y149_AO5),
.Q(CLBLM_R_X13Y149_SLICE_X19Y149_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y149_SLICE_X19Y149_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y149_SLICE_X19Y149_AO6),
.Q(CLBLM_R_X13Y149_SLICE_X19Y149_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y149_SLICE_X19Y149_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X13Y149_SLICE_X19Y149_CO6),
.Q(CLBLM_R_X13Y149_SLICE_X19Y149_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f00000f1f0011)
  ) CLBLM_R_X13Y149_SLICE_X19Y149_DLUT (
.I0(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.I1(CLBLM_R_X13Y148_SLICE_X18Y148_CO6),
.I2(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.I3(CLBLM_R_X5Y155_SLICE_X6Y155_DO6),
.I4(RIOB33_X105Y141_IOB_X1Y142_I),
.I5(CLBLM_R_X13Y155_SLICE_X19Y155_AO6),
.O5(CLBLM_R_X13Y149_SLICE_X19Y149_DO5),
.O6(CLBLM_R_X13Y149_SLICE_X19Y149_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000fe0efe0e)
  ) CLBLM_R_X13Y149_SLICE_X19Y149_CLUT (
.I0(CLBLM_R_X13Y149_SLICE_X18Y149_AQ),
.I1(CLBLM_R_X13Y149_SLICE_X19Y149_CQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y150_SLICE_X16Y150_A5Q),
.I4(1'b1),
.I5(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.O5(CLBLM_R_X13Y149_SLICE_X19Y149_CO5),
.O6(CLBLM_R_X13Y149_SLICE_X19Y149_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8a83aaa2ffffcccc)
  ) CLBLM_R_X13Y149_SLICE_X19Y149_BLUT (
.I0(CLBLM_R_X13Y149_SLICE_X18Y149_A5Q),
.I1(CLBLM_R_X13Y149_SLICE_X19Y149_A5Q),
.I2(CLBLM_R_X13Y149_SLICE_X19Y149_AQ),
.I3(CLBLM_R_X13Y149_SLICE_X18Y149_DO6),
.I4(CLBLM_L_X12Y148_SLICE_X17Y148_AO6),
.I5(1'b1),
.O5(CLBLM_R_X13Y149_SLICE_X19Y149_BO5),
.O6(CLBLM_R_X13Y149_SLICE_X19Y149_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb0b1b0b01c1b0c08)
  ) CLBLM_R_X13Y149_SLICE_X19Y149_ALUT (
.I0(CLBLM_R_X13Y149_SLICE_X18Y149_A5Q),
.I1(CLBLM_R_X13Y149_SLICE_X19Y149_A5Q),
.I2(CLBLM_R_X13Y149_SLICE_X19Y149_AQ),
.I3(CLBLM_R_X13Y149_SLICE_X18Y149_DO6),
.I4(CLBLM_L_X12Y148_SLICE_X17Y148_AO6),
.I5(1'b1),
.O5(CLBLM_R_X13Y149_SLICE_X19Y149_AO5),
.O6(CLBLM_R_X13Y149_SLICE_X19Y149_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y150_SLICE_X18Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y150_SLICE_X18Y150_AO6),
.Q(CLBLM_R_X13Y150_SLICE_X18Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y150_SLICE_X18Y150_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y150_SLICE_X18Y150_BO6),
.Q(CLBLM_R_X13Y150_SLICE_X18Y150_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y150_SLICE_X18Y150_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y150_SLICE_X18Y150_CO6),
.Q(CLBLM_R_X13Y150_SLICE_X18Y150_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h44444444a0a0a0a0)
  ) CLBLM_R_X13Y150_SLICE_X18Y150_DLUT (
.I0(CLBLM_R_X13Y149_SLICE_X18Y149_A5Q),
.I1(CLBLM_R_X13Y149_SLICE_X19Y149_A5Q),
.I2(CLBLM_R_X13Y149_SLICE_X19Y149_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y150_SLICE_X18Y150_DO5),
.O6(CLBLM_R_X13Y150_SLICE_X18Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0e4a0f5a0e4a0f5)
  ) CLBLM_R_X13Y150_SLICE_X18Y150_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.I2(CLBLM_R_X13Y151_SLICE_X18Y151_BQ),
.I3(CLBLM_L_X12Y150_SLICE_X17Y150_DO6),
.I4(RIOB33_X105Y141_IOB_X1Y142_I),
.I5(1'b1),
.O5(CLBLM_R_X13Y150_SLICE_X18Y150_CO5),
.O6(CLBLM_R_X13Y150_SLICE_X18Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hacaacccccc00cccc)
  ) CLBLM_R_X13Y150_SLICE_X18Y150_BLUT (
.I0(CLBLM_R_X13Y150_SLICE_X18Y150_DO6),
.I1(CLBLM_R_X13Y150_SLICE_X18Y150_BQ),
.I2(CLBLM_R_X11Y154_SLICE_X15Y154_DO6),
.I3(CLBLM_R_X13Y149_SLICE_X18Y149_DO6),
.I4(CLBLM_R_X13Y149_SLICE_X19Y149_BO5),
.I5(CLBLM_R_X13Y149_SLICE_X19Y149_AQ),
.O5(CLBLM_R_X13Y150_SLICE_X18Y150_BO5),
.O6(CLBLM_R_X13Y150_SLICE_X18Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccf500f000)
  ) CLBLM_R_X13Y150_SLICE_X18Y150_ALUT (
.I0(RIOB33_X105Y121_IOB_X1Y121_I),
.I1(CLBLM_L_X12Y146_SLICE_X16Y146_DQ),
.I2(CLBLM_R_X13Y150_SLICE_X18Y150_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X12Y149_SLICE_X16Y149_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y150_SLICE_X18Y150_AO5),
.O6(CLBLM_R_X13Y150_SLICE_X18Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y150_SLICE_X19Y150_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y150_SLICE_X19Y150_AO6),
.Q(CLBLM_R_X13Y150_SLICE_X19Y150_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y150_SLICE_X19Y150_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y150_SLICE_X19Y150_DO5),
.O6(CLBLM_R_X13Y150_SLICE_X19Y150_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y150_SLICE_X19Y150_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y150_SLICE_X19Y150_CO5),
.O6(CLBLM_R_X13Y150_SLICE_X19Y150_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y150_SLICE_X19Y150_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y150_SLICE_X19Y150_BO5),
.O6(CLBLM_R_X13Y150_SLICE_X19Y150_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffcc3300fedc3210)
  ) CLBLM_R_X13Y150_SLICE_X19Y150_ALUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X13Y150_SLICE_X19Y150_AQ),
.I3(CLBLL_L_X4Y149_SLICE_X4Y149_BQ),
.I4(CLBLM_R_X7Y148_SLICE_X9Y148_BQ),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X13Y150_SLICE_X19Y150_AO5),
.O6(CLBLM_R_X13Y150_SLICE_X19Y150_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y151_SLICE_X18Y151_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y151_SLICE_X18Y151_AO6),
.Q(CLBLM_R_X13Y151_SLICE_X18Y151_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y151_SLICE_X18Y151_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y151_SLICE_X18Y151_BO6),
.Q(CLBLM_R_X13Y151_SLICE_X18Y151_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y151_SLICE_X18Y151_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y151_SLICE_X18Y151_CO6),
.Q(CLBLM_R_X13Y151_SLICE_X18Y151_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y151_SLICE_X18Y151_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y151_SLICE_X18Y151_DO6),
.Q(CLBLM_R_X13Y151_SLICE_X18Y151_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffa50ffffea40)
  ) CLBLM_R_X13Y151_SLICE_X18Y151_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I2(CLBLM_R_X13Y151_SLICE_X18Y151_DQ),
.I3(CLBLM_R_X11Y151_SLICE_X15Y151_A5Q),
.I4(CLBLM_L_X10Y152_SLICE_X13Y152_DO6),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X13Y151_SLICE_X18Y151_DO5),
.O6(CLBLM_R_X13Y151_SLICE_X18Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h888888888dd88dd8)
  ) CLBLM_R_X13Y151_SLICE_X18Y151_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X12Y149_SLICE_X16Y149_CQ),
.I2(CLBLM_R_X13Y155_SLICE_X18Y155_BQ),
.I3(CLBLM_R_X11Y150_SLICE_X15Y150_AO5),
.I4(1'b1),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X13Y151_SLICE_X18Y151_CO5),
.O6(CLBLM_R_X13Y151_SLICE_X18Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdf80d08f5f00500)
  ) CLBLM_R_X13Y151_SLICE_X18Y151_BLUT (
.I0(CLBLM_R_X11Y149_SLICE_X15Y149_DO6),
.I1(CLBLM_R_X13Y151_SLICE_X18Y151_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X10Y151_SLICE_X12Y151_BQ),
.I4(CLBLM_R_X13Y153_SLICE_X18Y153_AQ),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X13Y151_SLICE_X18Y151_BO5),
.O6(CLBLM_R_X13Y151_SLICE_X18Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf5a0cccc5500)
  ) CLBLM_R_X13Y151_SLICE_X18Y151_ALUT (
.I0(CLBLM_R_X11Y149_SLICE_X15Y149_DO6),
.I1(CLBLM_R_X11Y156_SLICE_X14Y156_BQ),
.I2(CLBLM_R_X13Y151_SLICE_X18Y151_AQ),
.I3(CLBLM_L_X12Y153_SLICE_X16Y153_AQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X13Y151_SLICE_X18Y151_AO5),
.O6(CLBLM_R_X13Y151_SLICE_X18Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y151_SLICE_X19Y151_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y151_SLICE_X19Y151_DO5),
.O6(CLBLM_R_X13Y151_SLICE_X19Y151_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeffeeffeeffee)
  ) CLBLM_R_X13Y151_SLICE_X19Y151_CLUT (
.I0(CLBLM_R_X13Y151_SLICE_X18Y151_AQ),
.I1(CLBLM_R_X13Y152_SLICE_X19Y152_AQ),
.I2(1'b1),
.I3(CLBLM_L_X10Y151_SLICE_X12Y151_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y151_SLICE_X19Y151_CO5),
.O6(CLBLM_R_X13Y151_SLICE_X19Y151_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffeeffffffee)
  ) CLBLM_R_X13Y151_SLICE_X19Y151_BLUT (
.I0(CLBLM_R_X11Y151_SLICE_X14Y151_AQ),
.I1(CLBLM_R_X13Y153_SLICE_X18Y153_BQ),
.I2(1'b1),
.I3(CLBLM_L_X12Y153_SLICE_X16Y153_AQ),
.I4(CLBLM_R_X13Y153_SLICE_X19Y153_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y151_SLICE_X19Y151_BO5),
.O6(CLBLM_R_X13Y151_SLICE_X19Y151_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffff0000000f0)
  ) CLBLM_R_X13Y151_SLICE_X19Y151_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X13Y150_SLICE_X19Y150_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I5(CLBLL_L_X4Y149_SLICE_X4Y149_BQ),
.O5(CLBLM_R_X13Y151_SLICE_X19Y151_AO5),
.O6(CLBLM_R_X13Y151_SLICE_X19Y151_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y152_SLICE_X18Y152_A5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y152_SLICE_X18Y152_BO6),
.Q(CLBLM_R_X13Y152_SLICE_X18Y152_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y152_SLICE_X18Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y152_SLICE_X18Y152_AO6),
.Q(CLBLM_R_X13Y152_SLICE_X18Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y152_SLICE_X18Y152_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y152_SLICE_X18Y152_CO6),
.Q(CLBLM_R_X13Y152_SLICE_X18Y152_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3f0f2f3f3f3f1)
  ) CLBLM_R_X13Y152_SLICE_X18Y152_DLUT (
.I0(CLBLM_R_X13Y154_SLICE_X19Y154_AQ),
.I1(CLBLM_R_X13Y152_SLICE_X19Y152_CO6),
.I2(CLBLM_R_X11Y149_SLICE_X15Y149_DO6),
.I3(CLBLM_R_X5Y155_SLICE_X6Y155_BO6),
.I4(CLBLM_L_X12Y155_SLICE_X16Y155_AO5),
.I5(CLBLM_R_X7Y148_SLICE_X9Y148_BQ),
.O5(CLBLM_R_X13Y152_SLICE_X18Y152_DO5),
.O6(CLBLM_R_X13Y152_SLICE_X18Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haafeaaaa00540000)
  ) CLBLM_R_X13Y152_SLICE_X18Y152_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y152_SLICE_X18Y152_CQ),
.I2(CLBLM_L_X12Y150_SLICE_X17Y150_BQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I5(CLBLM_R_X13Y152_SLICE_X19Y152_BQ),
.O5(CLBLM_R_X13Y152_SLICE_X18Y152_CO5),
.O6(CLBLM_R_X13Y152_SLICE_X18Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff880088f5f5f5f5)
  ) CLBLM_R_X13Y152_SLICE_X18Y152_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X13Y152_SLICE_X18Y152_A5Q),
.I2(CLBLM_R_X5Y155_SLICE_X6Y155_DO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_L_X10Y151_SLICE_X13Y151_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y152_SLICE_X18Y152_BO5),
.O6(CLBLM_R_X13Y152_SLICE_X18Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf5a0cccc5500)
  ) CLBLM_R_X13Y152_SLICE_X18Y152_ALUT (
.I0(CLBLM_R_X11Y149_SLICE_X15Y149_DO6),
.I1(CLBLM_R_X11Y152_SLICE_X14Y152_AQ),
.I2(CLBLM_R_X13Y152_SLICE_X18Y152_AQ),
.I3(CLBLM_R_X11Y152_SLICE_X15Y152_BQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X13Y152_SLICE_X18Y152_AO5),
.O6(CLBLM_R_X13Y152_SLICE_X18Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y152_SLICE_X19Y152_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y152_SLICE_X19Y152_AO6),
.Q(CLBLM_R_X13Y152_SLICE_X19Y152_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y152_SLICE_X19Y152_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y152_SLICE_X19Y152_BO6),
.Q(CLBLM_R_X13Y152_SLICE_X19Y152_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y152_SLICE_X19Y152_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y152_SLICE_X19Y152_DO5),
.O6(CLBLM_R_X13Y152_SLICE_X19Y152_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa000055ba0000)
  ) CLBLM_R_X13Y152_SLICE_X19Y152_CLUT (
.I0(CLBLM_R_X13Y152_SLICE_X18Y152_AQ),
.I1(CLBLM_R_X13Y151_SLICE_X19Y151_CO6),
.I2(CLBLM_L_X12Y152_SLICE_X17Y152_CO6),
.I3(CLBLM_R_X13Y152_SLICE_X19Y152_BQ),
.I4(CLBLM_L_X12Y155_SLICE_X16Y155_AO5),
.I5(CLBLM_R_X13Y151_SLICE_X19Y151_BO6),
.O5(CLBLM_R_X13Y152_SLICE_X19Y152_CO5),
.O6(CLBLM_R_X13Y152_SLICE_X19Y152_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfd0df808f505f000)
  ) CLBLM_R_X13Y152_SLICE_X19Y152_BLUT (
.I0(CLBLM_R_X11Y149_SLICE_X15Y149_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y151_SLICE_X16Y151_BQ),
.I4(CLBLM_R_X13Y152_SLICE_X18Y152_AQ),
.I5(CLBLM_R_X13Y152_SLICE_X19Y152_BQ),
.O5(CLBLM_R_X13Y152_SLICE_X19Y152_BO5),
.O6(CLBLM_R_X13Y152_SLICE_X19Y152_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfddd3111eccc2000)
  ) CLBLM_R_X13Y152_SLICE_X19Y152_ALUT (
.I0(CLBLM_R_X11Y149_SLICE_X15Y149_DO6),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X13Y152_SLICE_X19Y152_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y157_SLICE_X15Y157_BQ),
.I5(CLBLM_R_X11Y152_SLICE_X15Y152_CQ),
.O5(CLBLM_R_X13Y152_SLICE_X19Y152_AO5),
.O6(CLBLM_R_X13Y152_SLICE_X19Y152_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y153_SLICE_X18Y153_C5_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y153_SLICE_X18Y153_CO5),
.Q(CLBLM_R_X13Y153_SLICE_X18Y153_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y153_SLICE_X18Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y153_SLICE_X18Y153_AO6),
.Q(CLBLM_R_X13Y153_SLICE_X18Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y153_SLICE_X18Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y153_SLICE_X18Y153_BO6),
.Q(CLBLM_R_X13Y153_SLICE_X18Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y153_SLICE_X18Y153_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y153_SLICE_X18Y153_CO6),
.Q(CLBLM_R_X13Y153_SLICE_X18Y153_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y153_SLICE_X18Y153_D_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y153_SLICE_X18Y153_DO6),
.Q(CLBLM_R_X13Y153_SLICE_X18Y153_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefefeeedcdcdccc)
  ) CLBLM_R_X13Y153_SLICE_X18Y153_DLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y152_SLICE_X13Y152_DO6),
.I2(CLBLM_R_X13Y153_SLICE_X18Y153_DQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I5(CLBLM_R_X13Y157_SLICE_X18Y157_AQ),
.O5(CLBLM_R_X13Y153_SLICE_X18Y153_DO5),
.O6(CLBLM_R_X13Y153_SLICE_X18Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8d8d8d8ffaa5500)
  ) CLBLM_R_X13Y153_SLICE_X18Y153_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_L_X10Y145_SLICE_X13Y145_CQ),
.I2(CLBLM_L_X10Y154_SLICE_X13Y154_AQ),
.I3(CLBLM_L_X12Y158_SLICE_X17Y158_BQ),
.I4(CLBLM_R_X13Y148_SLICE_X18Y148_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y153_SLICE_X18Y153_CO5),
.O6(CLBLM_R_X13Y153_SLICE_X18Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cf000fa0afa0a)
  ) CLBLM_R_X13Y153_SLICE_X18Y153_BLUT (
.I0(CLBLM_R_X13Y151_SLICE_X18Y151_BQ),
.I1(CLBLM_R_X13Y153_SLICE_X18Y153_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y156_SLICE_X17Y156_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X11Y149_SLICE_X15Y149_DO6),
.O5(CLBLM_R_X13Y153_SLICE_X18Y153_BO5),
.O6(CLBLM_R_X13Y153_SLICE_X18Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffccd80000ccd8)
  ) CLBLM_R_X13Y153_SLICE_X18Y153_ALUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I1(CLBLM_R_X13Y152_SLICE_X18Y152_CQ),
.I2(CLBLM_R_X13Y153_SLICE_X18Y153_AQ),
.I3(RIOB33_X105Y117_IOB_X1Y118_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X13Y154_SLICE_X18Y154_AQ),
.O5(CLBLM_R_X13Y153_SLICE_X18Y153_AO5),
.O6(CLBLM_R_X13Y153_SLICE_X18Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y153_SLICE_X19Y153_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y153_SLICE_X19Y153_AO6),
.Q(CLBLM_R_X13Y153_SLICE_X19Y153_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y153_SLICE_X19Y153_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y153_SLICE_X19Y153_BO6),
.Q(CLBLM_R_X13Y153_SLICE_X19Y153_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y153_SLICE_X19Y153_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y153_SLICE_X19Y153_CO6),
.Q(CLBLM_R_X13Y153_SLICE_X19Y153_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00c300ff0087)
  ) CLBLM_R_X13Y153_SLICE_X19Y153_DLUT (
.I0(CLBLM_R_X13Y155_SLICE_X19Y155_AO6),
.I1(CLBLM_R_X13Y154_SLICE_X19Y154_AQ),
.I2(CLBLM_R_X7Y148_SLICE_X9Y148_BQ),
.I3(CLBLM_R_X13Y152_SLICE_X19Y152_CO6),
.I4(CLBLM_L_X12Y155_SLICE_X16Y155_AO5),
.I5(CLBLM_R_X5Y155_SLICE_X6Y155_DO6),
.O5(CLBLM_R_X13Y153_SLICE_X19Y153_DO5),
.O6(CLBLM_R_X13Y153_SLICE_X19Y153_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaa0000fefe5454)
  ) CLBLM_R_X13Y153_SLICE_X19Y153_CLUT (
.I0(LIOB33_X0Y77_IOB_X0Y77_I),
.I1(CLBLM_R_X13Y153_SLICE_X19Y153_CQ),
.I2(CLBLM_L_X12Y153_SLICE_X17Y153_CQ),
.I3(1'b1),
.I4(CLBLM_L_X8Y155_SLICE_X11Y155_CQ),
.I5(CLBLM_R_X7Y146_SLICE_X8Y146_CO6),
.O5(CLBLM_R_X13Y153_SLICE_X19Y153_CO5),
.O6(CLBLM_R_X13Y153_SLICE_X19Y153_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfc0cfe0efe0e)
  ) CLBLM_R_X13Y153_SLICE_X19Y153_BLUT (
.I0(RIOB33_X105Y141_IOB_X1Y142_I),
.I1(CLBLM_R_X13Y153_SLICE_X19Y153_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y149_SLICE_X16Y149_B5Q),
.I4(1'b1),
.I5(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.O5(CLBLM_R_X13Y153_SLICE_X19Y153_BO5),
.O6(CLBLM_R_X13Y153_SLICE_X19Y153_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffd1110000d111)
  ) CLBLM_R_X13Y153_SLICE_X19Y153_ALUT (
.I0(CLBLM_R_X13Y153_SLICE_X19Y153_DO6),
.I1(CLBLM_R_X11Y149_SLICE_X15Y149_DO6),
.I2(CLBLM_R_X13Y153_SLICE_X19Y153_AQ),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_R_X13Y153_SLICE_X19Y153_BQ),
.O5(CLBLM_R_X13Y153_SLICE_X19Y153_AO5),
.O6(CLBLM_R_X13Y153_SLICE_X19Y153_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y154_SLICE_X18Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y154_SLICE_X18Y154_AO6),
.Q(CLBLM_R_X13Y154_SLICE_X18Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y154_SLICE_X18Y154_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y154_SLICE_X18Y154_BO6),
.Q(CLBLM_R_X13Y154_SLICE_X18Y154_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y154_SLICE_X18Y154_C_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y154_SLICE_X18Y154_CO6),
.Q(CLBLM_R_X13Y154_SLICE_X18Y154_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ff00aa00aa)
  ) CLBLM_R_X13Y154_SLICE_X18Y154_DLUT (
.I0(CLBLM_L_X12Y153_SLICE_X17Y153_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_L_X10Y150_SLICE_X13Y150_BQ),
.I4(1'b1),
.I5(CLBLM_R_X11Y152_SLICE_X15Y152_AQ),
.O5(CLBLM_R_X13Y154_SLICE_X18Y154_DO5),
.O6(CLBLM_R_X13Y154_SLICE_X18Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f0f0aa88)
  ) CLBLM_R_X13Y154_SLICE_X18Y154_CLUT (
.I0(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I1(CLBLM_R_X13Y154_SLICE_X18Y154_CQ),
.I2(CLBLM_L_X12Y151_SLICE_X17Y151_AQ),
.I3(CLBLM_R_X7Y152_SLICE_X9Y152_CO6),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(RIOB33_X105Y117_IOB_X1Y118_I),
.O5(CLBLM_R_X13Y154_SLICE_X18Y154_CO5),
.O6(CLBLM_R_X13Y154_SLICE_X18Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f0eef000f000)
  ) CLBLM_R_X13Y154_SLICE_X18Y154_BLUT (
.I0(CLBLM_R_X13Y148_SLICE_X18Y148_AQ),
.I1(CLBLM_R_X13Y154_SLICE_X18Y154_BQ),
.I2(CLBLM_L_X12Y153_SLICE_X17Y153_AQ),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(RIOB33_X105Y117_IOB_X1Y118_I),
.I5(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.O5(CLBLM_R_X13Y154_SLICE_X18Y154_BO5),
.O6(CLBLM_R_X13Y154_SLICE_X18Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f2f2ff00f2f2)
  ) CLBLM_R_X13Y154_SLICE_X18Y154_ALUT (
.I0(RIOB33_X105Y141_IOB_X1Y142_I),
.I1(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.I2(CLBLM_R_X13Y154_SLICE_X18Y154_AQ),
.I3(CLBLM_L_X8Y154_SLICE_X11Y154_CQ),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X13Y154_SLICE_X18Y154_AO5),
.O6(CLBLM_R_X13Y154_SLICE_X18Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y154_SLICE_X19Y154_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y154_SLICE_X19Y154_AO6),
.Q(CLBLM_R_X13Y154_SLICE_X19Y154_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y154_SLICE_X19Y154_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y154_SLICE_X19Y154_DO5),
.O6(CLBLM_R_X13Y154_SLICE_X19Y154_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y154_SLICE_X19Y154_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y154_SLICE_X19Y154_CO5),
.O6(CLBLM_R_X13Y154_SLICE_X19Y154_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y154_SLICE_X19Y154_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y154_SLICE_X19Y154_BO5),
.O6(CLBLM_R_X13Y154_SLICE_X19Y154_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffafcf80f0a0c08)
  ) CLBLM_R_X13Y154_SLICE_X19Y154_ALUT (
.I0(CLBLM_R_X13Y154_SLICE_X19Y154_AQ),
.I1(RIOB33_X105Y117_IOB_X1Y118_I),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X13Y154_SLICE_X18Y154_BQ),
.I4(CLBLM_R_X7Y149_SLICE_X9Y149_AQ),
.I5(CLBLM_L_X10Y155_SLICE_X13Y155_A5Q),
.O5(CLBLM_R_X13Y154_SLICE_X19Y154_AO5),
.O6(CLBLM_R_X13Y154_SLICE_X19Y154_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y155_SLICE_X18Y155_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y155_SLICE_X18Y155_AO6),
.Q(CLBLM_R_X13Y155_SLICE_X18Y155_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y155_SLICE_X18Y155_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y155_SLICE_X18Y155_BO6),
.Q(CLBLM_R_X13Y155_SLICE_X18Y155_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff000000ff)
  ) CLBLM_R_X13Y155_SLICE_X18Y155_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.O5(CLBLM_R_X13Y155_SLICE_X18Y155_DO5),
.O6(CLBLM_R_X13Y155_SLICE_X18Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000fcfc0000ffaa)
  ) CLBLM_R_X13Y155_SLICE_X18Y155_CLUT (
.I0(CLBLM_R_X11Y154_SLICE_X14Y154_AQ),
.I1(CLBLM_R_X13Y151_SLICE_X18Y151_DQ),
.I2(CLBLM_R_X13Y154_SLICE_X18Y154_CQ),
.I3(CLBLM_R_X7Y149_SLICE_X8Y149_AQ),
.I4(CLBLM_L_X10Y150_SLICE_X13Y150_BQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y155_SLICE_X18Y155_CO5),
.O6(CLBLM_R_X13Y155_SLICE_X18Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc05050a0a)
  ) CLBLM_R_X13Y155_SLICE_X18Y155_BLUT (
.I0(CLBLM_L_X12Y152_SLICE_X17Y152_BO5),
.I1(CLBLM_L_X12Y156_SLICE_X17Y156_AQ),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(1'b1),
.I4(CLBLM_L_X8Y155_SLICE_X11Y155_CQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y155_SLICE_X18Y155_BO5),
.O6(CLBLM_R_X13Y155_SLICE_X18Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hce02cc00cd01cc00)
  ) CLBLM_R_X13Y155_SLICE_X18Y155_ALUT (
.I0(CLBLM_R_X13Y155_SLICE_X18Y155_AQ),
.I1(LIOB33_X0Y77_IOB_X0Y77_I),
.I2(CLBLM_R_X7Y153_SLICE_X8Y153_AQ),
.I3(CLBLM_L_X12Y158_SLICE_X17Y158_BQ),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X12Y155_SLICE_X16Y155_AO6),
.O5(CLBLM_R_X13Y155_SLICE_X18Y155_AO5),
.O6(CLBLM_R_X13Y155_SLICE_X18Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y155_SLICE_X19Y155_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y155_SLICE_X19Y155_DO5),
.O6(CLBLM_R_X13Y155_SLICE_X19Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y155_SLICE_X19Y155_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y155_SLICE_X19Y155_CO5),
.O6(CLBLM_R_X13Y155_SLICE_X19Y155_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y155_SLICE_X19Y155_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y155_SLICE_X19Y155_BO5),
.O6(CLBLM_R_X13Y155_SLICE_X19Y155_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000005050)
  ) CLBLM_R_X13Y155_SLICE_X19Y155_ALUT (
.I0(RIOB33_X105Y135_IOB_X1Y136_I),
.I1(1'b1),
.I2(RIOB33_X105Y131_IOB_X1Y131_I),
.I3(1'b1),
.I4(CLBLL_L_X4Y158_SLICE_X4Y158_AO6),
.I5(RIOB33_X105Y135_IOB_X1Y135_I),
.O5(CLBLM_R_X13Y155_SLICE_X19Y155_AO5),
.O6(CLBLM_R_X13Y155_SLICE_X19Y155_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y156_SLICE_X18Y156_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y156_SLICE_X18Y156_AO6),
.Q(CLBLM_R_X13Y156_SLICE_X18Y156_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001000180008000)
  ) CLBLM_R_X13Y156_SLICE_X18Y156_DLUT (
.I0(CLBLM_L_X12Y157_SLICE_X17Y157_BQ),
.I1(CLBLM_R_X11Y157_SLICE_X14Y157_AQ),
.I2(CLBLM_L_X12Y156_SLICE_X17Y156_AQ),
.I3(CLBLM_L_X8Y154_SLICE_X10Y154_AQ),
.I4(1'b1),
.I5(CLBLM_L_X12Y158_SLICE_X16Y158_CO5),
.O5(CLBLM_R_X13Y156_SLICE_X18Y156_DO5),
.O6(CLBLM_R_X13Y156_SLICE_X18Y156_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffe7fffffff)
  ) CLBLM_R_X13Y156_SLICE_X18Y156_CLUT (
.I0(CLBLM_L_X12Y157_SLICE_X17Y157_BQ),
.I1(CLBLM_R_X11Y157_SLICE_X14Y157_AQ),
.I2(CLBLM_R_X11Y158_SLICE_X14Y158_AQ),
.I3(CLBLM_L_X8Y154_SLICE_X10Y154_AQ),
.I4(CLBLM_L_X12Y156_SLICE_X17Y156_AQ),
.I5(CLBLM_L_X12Y158_SLICE_X16Y158_CO5),
.O5(CLBLM_R_X13Y156_SLICE_X18Y156_CO5),
.O6(CLBLM_R_X13Y156_SLICE_X18Y156_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f070f0f0008)
  ) CLBLM_R_X13Y156_SLICE_X18Y156_BLUT (
.I0(CLBLM_R_X13Y156_SLICE_X18Y156_DO6),
.I1(CLBLM_L_X12Y157_SLICE_X16Y157_BQ),
.I2(CLBLM_R_X11Y159_SLICE_X15Y159_CO5),
.I3(CLBLM_L_X12Y158_SLICE_X16Y158_BO5),
.I4(CLBLM_R_X11Y158_SLICE_X15Y158_DO6),
.I5(CLBLM_R_X11Y158_SLICE_X14Y158_AQ),
.O5(CLBLM_R_X13Y156_SLICE_X18Y156_BO5),
.O6(CLBLM_R_X13Y156_SLICE_X18Y156_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f0f0fcfc)
  ) CLBLM_R_X13Y156_SLICE_X18Y156_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y141_IOB_X1Y142_I),
.I2(CLBLM_R_X13Y156_SLICE_X18Y156_AQ),
.I3(CLBLM_R_X13Y157_SLICE_X19Y157_AQ),
.I4(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.I5(LIOB33_X0Y77_IOB_X0Y77_I),
.O5(CLBLM_R_X13Y156_SLICE_X18Y156_AO5),
.O6(CLBLM_R_X13Y156_SLICE_X18Y156_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y156_SLICE_X19Y156_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y156_SLICE_X19Y156_AO6),
.Q(CLBLM_R_X13Y156_SLICE_X19Y156_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y156_SLICE_X19Y156_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y156_SLICE_X19Y156_DO5),
.O6(CLBLM_R_X13Y156_SLICE_X19Y156_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y156_SLICE_X19Y156_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y156_SLICE_X19Y156_CO5),
.O6(CLBLM_R_X13Y156_SLICE_X19Y156_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y156_SLICE_X19Y156_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y156_SLICE_X19Y156_BO5),
.O6(CLBLM_R_X13Y156_SLICE_X19Y156_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf5f0ccccf5f0)
  ) CLBLM_R_X13Y156_SLICE_X19Y156_ALUT (
.I0(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.I1(CLBLM_R_X7Y154_SLICE_X8Y154_BQ),
.I2(CLBLM_R_X13Y156_SLICE_X19Y156_AQ),
.I3(RIOB33_X105Y141_IOB_X1Y142_I),
.I4(LIOB33_X0Y77_IOB_X0Y77_I),
.I5(1'b1),
.O5(CLBLM_R_X13Y156_SLICE_X19Y156_AO5),
.O6(CLBLM_R_X13Y156_SLICE_X19Y156_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y157_SLICE_X18Y157_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(LIOB33_X0Y77_IOB_X0Y77_I),
.D(CLBLM_R_X11Y158_SLICE_X14Y158_BQ),
.Q(CLBLM_R_X13Y157_SLICE_X18Y157_AQ),
.R(CLBLM_R_X13Y155_SLICE_X18Y155_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffff7fffffff)
  ) CLBLM_R_X13Y157_SLICE_X18Y157_DLUT (
.I0(CLBLM_R_X11Y158_SLICE_X14Y158_AQ),
.I1(CLBLM_R_X13Y158_SLICE_X18Y158_BQ),
.I2(CLBLM_R_X13Y159_SLICE_X18Y159_DO6),
.I3(CLBLM_R_X11Y157_SLICE_X15Y157_BQ),
.I4(CLBLM_R_X11Y157_SLICE_X14Y157_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y157_SLICE_X18Y157_DO5),
.O6(CLBLM_R_X13Y157_SLICE_X18Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aa55aa556a5566)
  ) CLBLM_R_X13Y157_SLICE_X18Y157_CLUT (
.I0(CLBLM_R_X13Y157_SLICE_X19Y157_AQ),
.I1(CLBLM_R_X11Y157_SLICE_X14Y157_BQ),
.I2(CLBLM_R_X13Y157_SLICE_X19Y157_BO6),
.I3(CLBLM_R_X11Y158_SLICE_X15Y158_DO6),
.I4(CLBLM_R_X13Y157_SLICE_X18Y157_DO6),
.I5(CLBLM_L_X12Y158_SLICE_X16Y158_BO5),
.O5(CLBLM_R_X13Y157_SLICE_X18Y157_CO5),
.O6(CLBLM_R_X13Y157_SLICE_X18Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3331333333233333)
  ) CLBLM_R_X13Y157_SLICE_X18Y157_BLUT (
.I0(CLBLM_L_X12Y156_SLICE_X17Y156_AQ),
.I1(CLBLM_R_X11Y158_SLICE_X15Y158_DO6),
.I2(CLBLM_L_X12Y158_SLICE_X16Y158_CO5),
.I3(CLBLM_L_X12Y158_SLICE_X16Y158_BO5),
.I4(CLBLM_L_X12Y156_SLICE_X17Y156_BQ),
.I5(CLBLM_L_X8Y154_SLICE_X10Y154_AQ),
.O5(CLBLM_R_X13Y157_SLICE_X18Y157_BO5),
.O6(CLBLM_R_X13Y157_SLICE_X18Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafa0a0affff00ff)
  ) CLBLM_R_X13Y157_SLICE_X18Y157_ALUT (
.I0(CLBLM_L_X12Y157_SLICE_X16Y157_A5Q),
.I1(1'b1),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(RIOB33_X105Y143_IOB_X1Y143_I),
.I4(CLBLM_L_X12Y156_SLICE_X16Y156_AQ),
.I5(1'b1),
.O5(CLBLM_R_X13Y157_SLICE_X18Y157_AO5),
.O6(CLBLM_R_X13Y157_SLICE_X18Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y157_SLICE_X19Y157_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y157_SLICE_X19Y157_AO6),
.Q(CLBLM_R_X13Y157_SLICE_X19Y157_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y157_SLICE_X19Y157_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y157_SLICE_X19Y157_DO5),
.O6(CLBLM_R_X13Y157_SLICE_X19Y157_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y157_SLICE_X19Y157_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y157_SLICE_X19Y157_CO5),
.O6(CLBLM_R_X13Y157_SLICE_X19Y157_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000202)
  ) CLBLM_R_X13Y157_SLICE_X19Y157_BLUT (
.I0(CLBLM_R_X13Y159_SLICE_X18Y159_CO6),
.I1(CLBLM_R_X11Y157_SLICE_X15Y157_BQ),
.I2(CLBLM_R_X11Y157_SLICE_X14Y157_AQ),
.I3(1'b1),
.I4(CLBLM_R_X11Y158_SLICE_X14Y158_AQ),
.I5(CLBLM_R_X13Y158_SLICE_X18Y158_BQ),
.O5(CLBLM_R_X13Y157_SLICE_X19Y157_BO5),
.O6(CLBLM_R_X13Y157_SLICE_X19Y157_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aafcaa00aafc)
  ) CLBLM_R_X13Y157_SLICE_X19Y157_ALUT (
.I0(CLBLM_R_X13Y154_SLICE_X18Y154_CQ),
.I1(CLBLM_R_X11Y158_SLICE_X14Y158_DO5),
.I2(CLBLM_R_X13Y157_SLICE_X18Y157_CO6),
.I3(LIOB33_X0Y77_IOB_X0Y77_I),
.I4(CLBLM_R_X11Y159_SLICE_X15Y159_CO5),
.I5(1'b1),
.O5(CLBLM_R_X13Y157_SLICE_X19Y157_AO5),
.O6(CLBLM_R_X13Y157_SLICE_X19Y157_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y158_SLICE_X18Y158_A_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y158_SLICE_X18Y158_AO6),
.Q(CLBLM_R_X13Y158_SLICE_X18Y158_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X13Y158_SLICE_X18Y158_B_FDRE (
.C(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O),
.CE(1'b1),
.D(CLBLM_R_X13Y158_SLICE_X18Y158_BO6),
.Q(CLBLM_R_X13Y158_SLICE_X18Y158_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ffff2700)
  ) CLBLM_R_X13Y158_SLICE_X18Y158_DLUT (
.I0(CLBLM_R_X11Y157_SLICE_X15Y157_BQ),
.I1(CLBLM_R_X13Y158_SLICE_X19Y158_AO6),
.I2(CLBLM_R_X13Y158_SLICE_X19Y158_BO6),
.I3(CLBLM_R_X11Y158_SLICE_X14Y158_BQ),
.I4(CLBLM_R_X11Y158_SLICE_X15Y158_DO6),
.I5(CLBLM_L_X12Y158_SLICE_X16Y158_BO5),
.O5(CLBLM_R_X13Y158_SLICE_X18Y158_DO5),
.O6(CLBLM_R_X13Y158_SLICE_X18Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333cccc3333666c)
  ) CLBLM_R_X13Y158_SLICE_X18Y158_CLUT (
.I0(CLBLM_R_X11Y157_SLICE_X14Y157_CQ),
.I1(CLBLM_R_X13Y158_SLICE_X18Y158_AQ),
.I2(CLBLM_R_X13Y159_SLICE_X18Y159_BO6),
.I3(CLBLM_R_X13Y159_SLICE_X18Y159_AO6),
.I4(CLBLM_R_X11Y158_SLICE_X15Y158_DO6),
.I5(CLBLM_L_X12Y158_SLICE_X16Y158_BO5),
.O5(CLBLM_R_X13Y158_SLICE_X18Y158_CO5),
.O6(CLBLM_R_X13Y158_SLICE_X18Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0fff600000f06)
  ) CLBLM_R_X13Y158_SLICE_X18Y158_BLUT (
.I0(CLBLM_R_X13Y158_SLICE_X18Y158_DO6),
.I1(CLBLM_R_X13Y158_SLICE_X18Y158_BQ),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_R_X11Y158_SLICE_X14Y158_DO5),
.I4(CLBLM_R_X11Y159_SLICE_X15Y159_CO5),
.I5(CLBLM_L_X10Y158_SLICE_X13Y158_BQ),
.O5(CLBLM_R_X13Y158_SLICE_X18Y158_BO5),
.O6(CLBLM_R_X13Y158_SLICE_X18Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000ff0ff000fc0c)
  ) CLBLM_R_X13Y158_SLICE_X18Y158_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y158_SLICE_X14Y158_DO5),
.I2(LIOB33_X0Y77_IOB_X0Y77_I),
.I3(CLBLM_L_X12Y158_SLICE_X16Y158_AQ),
.I4(CLBLM_R_X11Y159_SLICE_X15Y159_CO5),
.I5(CLBLM_R_X13Y158_SLICE_X18Y158_CO6),
.O5(CLBLM_R_X13Y158_SLICE_X18Y158_AO5),
.O6(CLBLM_R_X13Y158_SLICE_X18Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y158_SLICE_X19Y158_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y158_SLICE_X19Y158_DO5),
.O6(CLBLM_R_X13Y158_SLICE_X19Y158_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y158_SLICE_X19Y158_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y158_SLICE_X19Y158_CO5),
.O6(CLBLM_R_X13Y158_SLICE_X19Y158_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffffffffffb)
  ) CLBLM_R_X13Y158_SLICE_X19Y158_BLUT (
.I0(CLBLM_L_X12Y156_SLICE_X17Y156_AQ),
.I1(CLBLM_L_X12Y158_SLICE_X16Y158_CO5),
.I2(CLBLM_L_X12Y157_SLICE_X17Y157_BQ),
.I3(CLBLM_L_X8Y154_SLICE_X10Y154_AQ),
.I4(CLBLM_R_X11Y158_SLICE_X14Y158_AQ),
.I5(CLBLM_R_X11Y157_SLICE_X14Y157_AQ),
.O5(CLBLM_R_X13Y158_SLICE_X19Y158_BO5),
.O6(CLBLM_R_X13Y158_SLICE_X19Y158_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfffffffffffffff)
  ) CLBLM_R_X13Y158_SLICE_X19Y158_ALUT (
.I0(CLBLM_L_X12Y156_SLICE_X17Y156_AQ),
.I1(CLBLM_L_X12Y158_SLICE_X16Y158_CO5),
.I2(CLBLM_L_X12Y157_SLICE_X17Y157_BQ),
.I3(CLBLM_L_X8Y154_SLICE_X10Y154_AQ),
.I4(CLBLM_R_X11Y158_SLICE_X14Y158_AQ),
.I5(CLBLM_R_X11Y157_SLICE_X14Y157_AQ),
.O5(CLBLM_R_X13Y158_SLICE_X19Y158_AO5),
.O6(CLBLM_R_X13Y158_SLICE_X19Y158_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0020a0a000000000)
  ) CLBLM_R_X13Y159_SLICE_X18Y159_DLUT (
.I0(CLBLM_L_X12Y157_SLICE_X17Y157_BQ),
.I1(CLBLM_L_X12Y158_SLICE_X17Y158_AQ),
.I2(CLBLM_L_X12Y156_SLICE_X17Y156_AQ),
.I3(CLBLM_L_X12Y158_SLICE_X16Y158_AQ),
.I4(CLBLM_R_X11Y159_SLICE_X15Y159_AQ),
.I5(CLBLM_L_X8Y154_SLICE_X10Y154_AQ),
.O5(CLBLM_R_X13Y159_SLICE_X18Y159_DO5),
.O6(CLBLM_R_X13Y159_SLICE_X18Y159_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000005040000)
  ) CLBLM_R_X13Y159_SLICE_X18Y159_CLUT (
.I0(CLBLM_L_X12Y157_SLICE_X17Y157_BQ),
.I1(CLBLM_L_X12Y158_SLICE_X17Y158_AQ),
.I2(CLBLM_L_X12Y156_SLICE_X17Y156_AQ),
.I3(CLBLM_L_X12Y158_SLICE_X16Y158_AQ),
.I4(CLBLM_R_X11Y159_SLICE_X15Y159_AQ),
.I5(CLBLM_L_X8Y154_SLICE_X10Y154_AQ),
.O5(CLBLM_R_X13Y159_SLICE_X18Y159_CO5),
.O6(CLBLM_R_X13Y159_SLICE_X18Y159_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000000000)
  ) CLBLM_R_X13Y159_SLICE_X18Y159_BLUT (
.I0(CLBLM_R_X13Y159_SLICE_X18Y159_DO6),
.I1(CLBLM_R_X11Y157_SLICE_X15Y157_BQ),
.I2(CLBLM_R_X11Y158_SLICE_X14Y158_AQ),
.I3(CLBLM_R_X13Y158_SLICE_X18Y158_BQ),
.I4(CLBLM_R_X13Y157_SLICE_X19Y157_AQ),
.I5(CLBLM_R_X11Y157_SLICE_X14Y157_AQ),
.O5(CLBLM_R_X13Y159_SLICE_X18Y159_BO5),
.O6(CLBLM_R_X13Y159_SLICE_X18Y159_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000100000000)
  ) CLBLM_R_X13Y159_SLICE_X18Y159_ALUT (
.I0(CLBLM_R_X11Y157_SLICE_X14Y157_AQ),
.I1(CLBLM_R_X13Y158_SLICE_X18Y158_BQ),
.I2(CLBLM_R_X11Y158_SLICE_X14Y158_AQ),
.I3(CLBLM_R_X11Y157_SLICE_X15Y157_BQ),
.I4(CLBLM_R_X13Y157_SLICE_X19Y157_AQ),
.I5(CLBLM_R_X13Y159_SLICE_X18Y159_CO6),
.O5(CLBLM_R_X13Y159_SLICE_X18Y159_AO5),
.O6(CLBLM_R_X13Y159_SLICE_X18Y159_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y159_SLICE_X19Y159_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y159_SLICE_X19Y159_DO5),
.O6(CLBLM_R_X13Y159_SLICE_X19Y159_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y159_SLICE_X19Y159_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y159_SLICE_X19Y159_CO5),
.O6(CLBLM_R_X13Y159_SLICE_X19Y159_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y159_SLICE_X19Y159_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y159_SLICE_X19Y159_BO5),
.O6(CLBLM_R_X13Y159_SLICE_X19Y159_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X13Y159_SLICE_X19Y159_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X13Y159_SLICE_X19Y159_AO5),
.O6(CLBLM_R_X13Y159_SLICE_X19Y159_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y141_SLICE_X162Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y141_SLICE_X162Y141_DO5),
.O6(CLBLM_R_X103Y141_SLICE_X162Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y141_SLICE_X162Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y141_SLICE_X162Y141_CO5),
.O6(CLBLM_R_X103Y141_SLICE_X162Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y141_SLICE_X162Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y141_SLICE_X162Y141_BO5),
.O6(CLBLM_R_X103Y141_SLICE_X162Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y141_SLICE_X162Y141_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y141_SLICE_X162Y141_AO5),
.O6(CLBLM_R_X103Y141_SLICE_X162Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y141_SLICE_X163Y141_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y141_SLICE_X163Y141_DO5),
.O6(CLBLM_R_X103Y141_SLICE_X163Y141_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y141_SLICE_X163Y141_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y141_SLICE_X163Y141_CO5),
.O6(CLBLM_R_X103Y141_SLICE_X163Y141_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y141_SLICE_X163Y141_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y141_SLICE_X163Y141_BO5),
.O6(CLBLM_R_X103Y141_SLICE_X163Y141_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha000a00088880000)
  ) CLBLM_R_X103Y141_SLICE_X163Y141_ALUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(RIOB33_X105Y139_IOB_X1Y140_I),
.I2(RIOB33_X105Y139_IOB_X1Y139_I),
.I3(RIOB33_X105Y137_IOB_X1Y138_I),
.I4(RIOB33_X105Y141_IOB_X1Y141_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y141_SLICE_X163Y141_AO5),
.O6(CLBLM_R_X103Y141_SLICE_X163Y141_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_DO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_CO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_BO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X162Y169_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X162Y169_AO5),
.O6(CLBLM_R_X103Y169_SLICE_X162Y169_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_DO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_CO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_BO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0ffffccccffff)
  ) CLBLM_R_X103Y169_SLICE_X163Y169_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y156_SLICE_X15Y156_BQ),
.I2(CLBLM_L_X12Y155_SLICE_X16Y155_AQ),
.I3(1'b1),
.I4(RIOB33_X105Y143_IOB_X1Y143_I),
.I5(1'b1),
.O5(CLBLM_R_X103Y169_SLICE_X163Y169_AO5),
.O6(CLBLM_R_X103Y169_SLICE_X163Y169_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X162Y172_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X162Y172_DO5),
.O6(CLBLM_R_X103Y172_SLICE_X162Y172_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X162Y172_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X162Y172_CO5),
.O6(CLBLM_R_X103Y172_SLICE_X162Y172_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X162Y172_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X162Y172_BO5),
.O6(CLBLM_R_X103Y172_SLICE_X162Y172_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X162Y172_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X162Y172_AO5),
.O6(CLBLM_R_X103Y172_SLICE_X162Y172_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X163Y172_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X163Y172_DO5),
.O6(CLBLM_R_X103Y172_SLICE_X163Y172_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X163Y172_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X163Y172_CO5),
.O6(CLBLM_R_X103Y172_SLICE_X163Y172_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y172_SLICE_X163Y172_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X163Y172_BO5),
.O6(CLBLM_R_X103Y172_SLICE_X163Y172_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fff0ffffff00ff)
  ) CLBLM_R_X103Y172_SLICE_X163Y172_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X13Y156_SLICE_X18Y156_AQ),
.I3(RIOB33_X105Y143_IOB_X1Y143_I),
.I4(CLBLM_L_X12Y156_SLICE_X16Y156_BQ),
.I5(1'b1),
.O5(CLBLM_R_X103Y172_SLICE_X163Y172_AO5),
.O6(CLBLM_R_X103Y172_SLICE_X163Y172_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_DO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_CO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_BO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X162Y174_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X162Y174_AO5),
.O6(CLBLM_R_X103Y174_SLICE_X162Y174_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_DO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_CO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_BO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcfcfcfcfffff0f0f)
  ) CLBLM_R_X103Y174_SLICE_X163Y174_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X13Y153_SLICE_X19Y153_BQ),
.I2(RIOB33_X105Y143_IOB_X1Y143_I),
.I3(1'b1),
.I4(CLBLM_R_X13Y156_SLICE_X19Y156_AQ),
.I5(1'b1),
.O5(CLBLM_R_X103Y174_SLICE_X163Y174_AO5),
.O6(CLBLM_R_X103Y174_SLICE_X163Y174_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_DO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_CO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_BO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X162Y177_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X162Y177_AO5),
.O6(CLBLM_R_X103Y177_SLICE_X162Y177_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_DO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_CO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_BO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5f5f5f5ffff5555)
  ) CLBLM_R_X103Y177_SLICE_X163Y177_ALUT (
.I0(RIOB33_X105Y143_IOB_X1Y143_I),
.I1(1'b1),
.I2(CLBLM_R_X13Y154_SLICE_X18Y154_AQ),
.I3(1'b1),
.I4(CLBLM_R_X13Y157_SLICE_X18Y157_AQ),
.I5(1'b1),
.O5(CLBLM_R_X103Y177_SLICE_X163Y177_AO5),
.O6(CLBLM_R_X103Y177_SLICE_X163Y177_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(LIOB33_X0Y77_IOB_X0Y78_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y51_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y51_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y51_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y51_IOB_X0Y52_IBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_IPAD),
.O(LIOB33_X0Y51_IOB_X0Y52_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y53_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y53_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y53_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y53_IOB_X0Y54_IBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_IPAD),
.O(LIOB33_X0Y53_IOB_X0Y54_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y55_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y55_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y55_IOB_X0Y56_IBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_IPAD),
.O(LIOB33_X0Y55_IOB_X0Y56_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y57_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y57_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y57_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y57_IOB_X0Y58_IBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_IPAD),
.O(LIOB33_X0Y57_IOB_X0Y58_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y59_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y59_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y59_IOB_X0Y60_IBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_IPAD),
.O(LIOB33_X0Y59_IOB_X0Y60_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y61_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y61_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y61_IOB_X0Y62_IBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_IPAD),
.O(LIOB33_X0Y61_IOB_X0Y62_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y63_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y63_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y63_IOB_X0Y64_IBUF (
.I(LIOB33_X0Y63_IOB_X0Y64_IPAD),
.O(LIOB33_X0Y63_IOB_X0Y64_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y65_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y65_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y65_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y65_IOB_X0Y66_IBUF (
.I(LIOB33_X0Y65_IOB_X0Y66_IPAD),
.O(LIOB33_X0Y65_IOB_X0Y66_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y67_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y67_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y67_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y67_IOB_X0Y68_IBUF (
.I(LIOB33_X0Y67_IOB_X0Y68_IPAD),
.O(LIOB33_X0Y67_IOB_X0Y68_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y69_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y69_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y69_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y69_IOB_X0Y70_IBUF (
.I(LIOB33_X0Y69_IOB_X0Y70_IPAD),
.O(LIOB33_X0Y69_IOB_X0Y70_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y71_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y71_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y71_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y71_IOB_X0Y72_IBUF (
.I(LIOB33_X0Y71_IOB_X0Y72_IPAD),
.O(LIOB33_X0Y71_IOB_X0Y72_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y73_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y73_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y73_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y73_IOB_X0Y74_IBUF (
.I(LIOB33_X0Y73_IOB_X0Y74_IPAD),
.O(LIOB33_X0Y73_IOB_X0Y74_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y75_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y75_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y75_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y75_IOB_X0Y76_IBUF (
.I(LIOB33_X0Y75_IOB_X0Y76_IPAD),
.O(LIOB33_X0Y75_IOB_X0Y76_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y77_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y77_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y77_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y77_IOB_X0Y78_IBUF (
.I(LIOB33_X0Y77_IOB_X0Y78_IPAD),
.O(LIOB33_X0Y77_IOB_X0Y78_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y79_IOB_X0Y79_IBUF (
.I(LIOB33_X0Y79_IOB_X0Y79_IPAD),
.O(LIOB33_X0Y79_IOB_X0Y79_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y79_IOB_X0Y80_OBUF (
.I(CLBLL_L_X2Y140_SLICE_X0Y140_AO6),
.O(LIOB33_X0Y79_IOB_X0Y80_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y101_OBUF (
.I(CLBLL_L_X2Y139_SLICE_X0Y139_AO6),
.O(LIOB33_X0Y101_IOB_X0Y101_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y101_IOB_X0Y102_OBUF (
.I(CLBLL_L_X2Y139_SLICE_X0Y139_AO5),
.O(LIOB33_X0Y101_IOB_X0Y102_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y103_OBUF (
.I(CLBLL_L_X2Y139_SLICE_X0Y139_BO6),
.O(LIOB33_X0Y103_IOB_X0Y103_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y103_IOB_X0Y104_OBUF (
.I(CLBLL_L_X2Y139_SLICE_X0Y139_BO5),
.O(LIOB33_X0Y103_IOB_X0Y104_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y105_OBUF (
.I(CLBLL_L_X2Y140_SLICE_X0Y140_BO6),
.O(LIOB33_X0Y105_IOB_X0Y105_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y105_IOB_X0Y106_OBUF (
.I(CLBLL_L_X2Y140_SLICE_X0Y140_BO5),
.O(LIOB33_X0Y105_IOB_X0Y106_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y107_OBUF (
.I(CLBLM_R_X3Y142_SLICE_X3Y142_CO6),
.O(LIOB33_X0Y107_IOB_X0Y107_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y107_IOB_X0Y108_OBUF (
.I(CLBLM_R_X3Y151_SLICE_X3Y151_BO6),
.O(LIOB33_X0Y107_IOB_X0Y108_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y109_OBUF (
.I(CLBLM_R_X3Y142_SLICE_X3Y142_DO6),
.O(LIOB33_X0Y109_IOB_X0Y109_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y109_IOB_X0Y110_OBUF (
.I(CLBLM_R_X3Y142_SLICE_X3Y142_BO6),
.O(LIOB33_X0Y109_IOB_X0Y110_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y111_OBUF (
.I(1'b0),
.O(LIOB33_X0Y111_IOB_X0Y111_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y112_OBUF (
.I(CLBLM_L_X12Y151_SLICE_X16Y151_C5Q),
.O(LIOB33_X0Y111_IOB_X0Y112_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y113_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_I),
.O(LIOB33_X0Y113_IOB_X0Y113_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y113_IOB_X0Y114_OBUF (
.I(CLBLM_L_X8Y146_SLICE_X10Y146_BQ),
.O(LIOB33_X0Y113_IOB_X0Y114_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y115_OBUF (
.I(CLBLM_L_X12Y151_SLICE_X16Y151_CQ),
.O(LIOB33_X0Y115_IOB_X0Y115_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y115_IOB_X0Y116_OBUF (
.I(CLBLM_R_X11Y144_SLICE_X15Y144_AQ),
.O(LIOB33_X0Y115_IOB_X0Y116_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y117_OBUF (
.I(CLBLM_R_X5Y147_SLICE_X7Y147_CQ),
.O(LIOB33_X0Y117_IOB_X0Y117_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y118_OBUF (
.I(CLBLM_R_X5Y148_SLICE_X7Y148_BQ),
.O(LIOB33_X0Y117_IOB_X0Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUF (
.I(CLBLM_R_X11Y149_SLICE_X15Y149_AQ),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUF (
.I(CLBLM_L_X12Y149_SLICE_X16Y149_BQ),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUF (
.I(CLBLM_R_X11Y144_SLICE_X15Y144_A5Q),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUF (
.I(CLBLL_L_X4Y149_SLICE_X5Y149_A5Q),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUF (
.I(CLBLM_L_X8Y146_SLICE_X10Y146_B5Q),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(CLBLM_R_X5Y148_SLICE_X7Y148_B5Q),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y125_OBUF (
.I(CLBLM_L_X8Y154_SLICE_X10Y154_C5Q),
.O(LIOB33_X0Y125_IOB_X0Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y126_OBUF (
.I(CLBLL_L_X4Y147_SLICE_X5Y147_AQ),
.O(LIOB33_X0Y125_IOB_X0Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y127_OBUF (
.I(CLBLL_L_X4Y152_SLICE_X4Y152_AQ),
.O(LIOB33_X0Y127_IOB_X0Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y128_OBUF (
.I(CLBLM_R_X3Y151_SLICE_X2Y151_AQ),
.O(LIOB33_X0Y127_IOB_X0Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y129_OBUF (
.I(CLBLL_L_X4Y151_SLICE_X5Y151_CQ),
.O(LIOB33_X0Y129_IOB_X0Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y130_OBUF (
.I(CLBLL_L_X52Y126_SLICE_X78Y126_AO6),
.O(LIOB33_X0Y129_IOB_X0Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y131_OBUF (
.I(CLBLM_L_X10Y144_SLICE_X12Y144_AO5),
.O(LIOB33_X0Y131_IOB_X0Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y132_OBUF (
.I(CLBLM_L_X10Y144_SLICE_X12Y144_AQ),
.O(LIOB33_X0Y131_IOB_X0Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y133_OBUF (
.I(CLBLM_R_X5Y146_SLICE_X6Y146_A5Q),
.O(LIOB33_X0Y133_IOB_X0Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y134_OBUF (
.I(CLBLM_R_X7Y145_SLICE_X8Y145_AQ),
.O(LIOB33_X0Y133_IOB_X0Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y135_OBUF (
.I(CLBLM_R_X5Y146_SLICE_X6Y146_AQ),
.O(LIOB33_X0Y135_IOB_X0Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUF (
.I(CLBLM_R_X7Y144_SLICE_X8Y144_AQ),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUF (
.I(CLBLM_R_X5Y144_SLICE_X6Y144_BQ),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUF (
.I(CLBLM_R_X5Y146_SLICE_X6Y146_BQ),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUF (
.I(CLBLM_R_X5Y144_SLICE_X6Y144_AQ),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUF (
.I(CLBLL_L_X4Y147_SLICE_X5Y147_BQ),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y141_OBUF (
.I(CLBLM_R_X5Y147_SLICE_X6Y147_AQ),
.O(LIOB33_X0Y141_IOB_X0Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y142_OBUF (
.I(LIOB33_X0Y53_IOB_X0Y54_I),
.O(LIOB33_X0Y141_IOB_X0Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y143_IOB_X0Y143_OBUF (
.I(LIOB33_X0Y55_IOB_X0Y55_I),
.O(LIOB33_X0Y143_IOB_X0Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y145_OBUF (
.I(LIOB33_X0Y57_IOB_X0Y58_I),
.O(LIOB33_X0Y145_IOB_X0Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y146_OBUF (
.I(LIOB33_X0Y59_IOB_X0Y59_I),
.O(LIOB33_X0Y145_IOB_X0Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y147_OBUF (
.I(LIOB33_X0Y71_IOB_X0Y71_I),
.O(LIOB33_X0Y147_IOB_X0Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y148_OBUF (
.I(LIOB33_X0Y61_IOB_X0Y61_I),
.O(LIOB33_X0Y147_IOB_X0Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y151_OBUF (
.I(LIOB33_X0Y65_IOB_X0Y65_I),
.O(LIOB33_X0Y151_IOB_X0Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y151_IOB_X0Y152_OBUF (
.I(LIOB33_X0Y65_IOB_X0Y66_I),
.O(LIOB33_X0Y151_IOB_X0Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y153_OBUF (
.I(LIOB33_X0Y67_IOB_X0Y67_I),
.O(LIOB33_X0Y153_IOB_X0Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y153_IOB_X0Y154_OBUF (
.I(LIOB33_X0Y67_IOB_X0Y68_I),
.O(LIOB33_X0Y153_IOB_X0Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y155_OBUF (
.I(LIOB33_X0Y69_IOB_X0Y70_I),
.O(LIOB33_X0Y155_IOB_X0Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y155_IOB_X0Y156_OBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_I),
.O(LIOB33_X0Y155_IOB_X0Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y157_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_I),
.O(LIOB33_X0Y157_IOB_X0Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y157_IOB_X0Y158_OBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_I),
.O(LIOB33_X0Y157_IOB_X0Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y159_OBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_I),
.O(LIOB33_X0Y159_IOB_X0Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y159_IOB_X0Y160_OBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_I),
.O(LIOB33_X0Y159_IOB_X0Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y161_OBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_I),
.O(LIOB33_X0Y161_IOB_X0Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y161_IOB_X0Y162_OBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_I),
.O(LIOB33_X0Y161_IOB_X0Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y163_OBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_I),
.O(LIOB33_X0Y163_IOB_X0Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y163_IOB_X0Y164_OBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_I),
.O(LIOB33_X0Y163_IOB_X0Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y165_OBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_I),
.O(LIOB33_X0Y165_IOB_X0Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y165_IOB_X0Y166_OBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_I),
.O(LIOB33_X0Y165_IOB_X0Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y167_OBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_I),
.O(LIOB33_X0Y167_IOB_X0Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y167_IOB_X0Y168_OBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_I),
.O(LIOB33_X0Y167_IOB_X0Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y169_OBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_I),
.O(LIOB33_X0Y169_IOB_X0Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y169_IOB_X0Y170_OBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.O(LIOB33_X0Y169_IOB_X0Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y171_OBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.O(LIOB33_X0Y171_IOB_X0Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y171_IOB_X0Y172_OBUF (
.I(CLBLM_R_X103Y141_SLICE_X163Y141_AO6),
.O(LIOB33_X0Y171_IOB_X0Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y173_OBUF (
.I(CLBLM_R_X103Y141_SLICE_X163Y141_AO5),
.O(LIOB33_X0Y173_IOB_X0Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y173_IOB_X0Y174_OBUF (
.I(CLBLM_L_X10Y163_SLICE_X13Y163_AO6),
.O(LIOB33_X0Y173_IOB_X0Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y175_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_I),
.O(LIOB33_X0Y175_IOB_X0Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y175_IOB_X0Y176_OBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_I),
.O(LIOB33_X0Y175_IOB_X0Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y177_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_I),
.O(LIOB33_X0Y177_IOB_X0Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y177_IOB_X0Y178_OBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_I),
.O(LIOB33_X0Y177_IOB_X0Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y179_OBUF (
.I(RIOB33_X105Y131_IOB_X1Y131_I),
.O(LIOB33_X0Y179_IOB_X0Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y179_IOB_X0Y180_OBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_I),
.O(LIOB33_X0Y179_IOB_X0Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y181_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_I),
.O(LIOB33_X0Y181_IOB_X0Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y181_IOB_X0Y182_OBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_I),
.O(LIOB33_X0Y181_IOB_X0Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y183_OBUF (
.I(RIOB33_X105Y135_IOB_X1Y135_I),
.O(LIOB33_X0Y183_IOB_X0Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y183_IOB_X0Y184_OBUF (
.I(RIOB33_X105Y135_IOB_X1Y136_I),
.O(LIOB33_X0Y183_IOB_X0Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y185_OBUF (
.I(RIOB33_X105Y137_IOB_X1Y137_I),
.O(LIOB33_X0Y185_IOB_X0Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y185_IOB_X0Y186_OBUF (
.I(RIOB33_X105Y143_IOB_X1Y143_I),
.O(LIOB33_X0Y185_IOB_X0Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y187_OBUF (
.I(RIOB33_X105Y143_IOB_X1Y144_I),
.O(LIOB33_X0Y187_IOB_X0Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y187_IOB_X0Y188_OBUF (
.I(RIOB33_X105Y145_IOB_X1Y145_I),
.O(LIOB33_X0Y187_IOB_X0Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y189_OBUF (
.I(RIOB33_X105Y145_IOB_X1Y146_I),
.O(LIOB33_X0Y189_IOB_X0Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y189_IOB_X0Y190_OBUF (
.I(RIOB33_X105Y147_IOB_X1Y147_I),
.O(LIOB33_X0Y189_IOB_X0Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y191_OBUF (
.I(RIOB33_X105Y147_IOB_X1Y148_I),
.O(LIOB33_X0Y191_IOB_X0Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y191_IOB_X0Y192_OBUF (
.I(LIOB33_X0Y51_IOB_X0Y52_I),
.O(LIOB33_X0Y191_IOB_X0Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y193_OBUF (
.I(LIOB33_X0Y55_IOB_X0Y56_I),
.O(LIOB33_X0Y193_IOB_X0Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y193_IOB_X0Y194_OBUF (
.I(LIOB33_X0Y59_IOB_X0Y60_I),
.O(LIOB33_X0Y193_IOB_X0Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y195_OBUF (
.I(LIOB33_X0Y63_IOB_X0Y64_I),
.O(LIOB33_X0Y195_IOB_X0Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y195_IOB_X0Y196_OBUF (
.I(LIOB33_X0Y69_IOB_X0Y69_I),
.O(LIOB33_X0Y195_IOB_X0Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y197_OBUF (
.I(LIOB33_X0Y71_IOB_X0Y72_I),
.O(LIOB33_X0Y197_IOB_X0Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y197_IOB_X0Y198_OBUF (
.I(LIOB33_X0Y73_IOB_X0Y73_I),
.O(LIOB33_X0Y197_IOB_X0Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y50_IOB_X0Y50_IBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_IPAD),
.O(LIOB33_SING_X0Y50_IOB_X0Y50_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y100_IOB_X0Y100_OBUF (
.I(CLBLL_L_X2Y140_SLICE_X0Y140_AO5),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_OBUF (
.I(LIOB33_X0Y61_IOB_X0Y62_I),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y150_IOB_X0Y150_OBUF (
.I(LIOB33_X0Y63_IOB_X0Y63_I),
.O(LIOB33_SING_X0Y150_IOB_X0Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y199_IOB_X0Y199_OBUF (
.I(LIOB33_X0Y73_IOB_X0Y74_I),
.O(LIOB33_SING_X0Y199_IOB_X0Y199_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y101_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y102_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y103_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y104_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y105_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y105_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y106_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y107_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y108_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y109_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y110_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y111_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y112_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y113_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y114_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y114_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y115_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y115_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y115_IOB_X1Y116_IBUF (
.I(RIOB33_X105Y115_IOB_X1Y116_IPAD),
.O(RIOB33_X105Y115_IOB_X1Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y117_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y117_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y117_IOB_X1Y118_IBUF (
.I(RIOB33_X105Y117_IOB_X1Y118_IPAD),
.O(RIOB33_X105Y117_IOB_X1Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y119_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y119_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y119_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y119_IOB_X1Y120_IBUF (
.I(RIOB33_X105Y119_IOB_X1Y120_IPAD),
.O(RIOB33_X105Y119_IOB_X1Y120_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y121_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y121_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y121_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y121_IOB_X1Y122_IBUF (
.I(RIOB33_X105Y121_IOB_X1Y122_IPAD),
.O(RIOB33_X105Y121_IOB_X1Y122_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y123_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y123_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y123_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y123_IOB_X1Y124_IBUF (
.I(RIOB33_X105Y123_IOB_X1Y124_IPAD),
.O(RIOB33_X105Y123_IOB_X1Y124_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y125_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y125_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y125_IOB_X1Y126_IBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_IPAD),
.O(RIOB33_X105Y125_IOB_X1Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y127_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y127_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y127_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y127_IOB_X1Y128_IBUF (
.I(RIOB33_X105Y127_IOB_X1Y128_IPAD),
.O(RIOB33_X105Y127_IOB_X1Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y129_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y129_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y129_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y129_IOB_X1Y130_IBUF (
.I(RIOB33_X105Y129_IOB_X1Y130_IPAD),
.O(RIOB33_X105Y129_IOB_X1Y130_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y131_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y131_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y131_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y131_IOB_X1Y132_IBUF (
.I(RIOB33_X105Y131_IOB_X1Y132_IPAD),
.O(RIOB33_X105Y131_IOB_X1Y132_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y133_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y133_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y133_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y133_IOB_X1Y134_IBUF (
.I(RIOB33_X105Y133_IOB_X1Y134_IPAD),
.O(RIOB33_X105Y133_IOB_X1Y134_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y135_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y135_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y135_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y135_IOB_X1Y136_IBUF (
.I(RIOB33_X105Y135_IOB_X1Y136_IPAD),
.O(RIOB33_X105Y135_IOB_X1Y136_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y137_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y137_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y137_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y137_IOB_X1Y138_IBUF (
.I(RIOB33_X105Y137_IOB_X1Y138_IPAD),
.O(RIOB33_X105Y137_IOB_X1Y138_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y139_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y139_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y139_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y139_IOB_X1Y140_IBUF (
.I(RIOB33_X105Y139_IOB_X1Y140_IPAD),
.O(RIOB33_X105Y139_IOB_X1Y140_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y141_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y141_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y141_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y141_IOB_X1Y142_IBUF (
.I(RIOB33_X105Y141_IOB_X1Y142_IPAD),
.O(RIOB33_X105Y141_IOB_X1Y142_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y143_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y143_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y143_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y143_IOB_X1Y144_IBUF (
.I(RIOB33_X105Y143_IOB_X1Y144_IPAD),
.O(RIOB33_X105Y143_IOB_X1Y144_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y145_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y145_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y145_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y145_IOB_X1Y146_IBUF (
.I(RIOB33_X105Y145_IOB_X1Y146_IPAD),
.O(RIOB33_X105Y145_IOB_X1Y146_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y147_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y147_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y147_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y147_IOB_X1Y148_IBUF (
.I(RIOB33_X105Y147_IOB_X1Y148_IPAD),
.O(RIOB33_X105Y147_IOB_X1Y148_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y151_OBUF (
.I(LIOB33_X0Y75_IOB_X0Y76_I),
.O(RIOB33_X105Y151_IOB_X1Y151_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y151_IOB_X1Y152_OBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O(RIOB33_X105Y151_IOB_X1Y152_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y153_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_I),
.O(RIOB33_X105Y153_IOB_X1Y153_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y153_IOB_X1Y154_OBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_I),
.O(RIOB33_X105Y153_IOB_X1Y154_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y155_OBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_I),
.O(RIOB33_X105Y155_IOB_X1Y155_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y155_IOB_X1Y156_OBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_I),
.O(RIOB33_X105Y155_IOB_X1Y156_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y157_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y126_I),
.O(RIOB33_X105Y157_IOB_X1Y157_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y157_IOB_X1Y158_OBUF (
.I(CLBLL_L_X36Y150_SLICE_X54Y150_AO6),
.O(RIOB33_X105Y157_IOB_X1Y158_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y159_OBUF (
.I(CLBLM_R_X13Y154_SLICE_X18Y154_DO6),
.O(RIOB33_X105Y159_IOB_X1Y159_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y159_IOB_X1Y160_OBUF (
.I(CLBLM_R_X13Y155_SLICE_X18Y155_CO6),
.O(RIOB33_X105Y159_IOB_X1Y160_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y161_OBUF (
.I(CLBLM_R_X13Y155_SLICE_X18Y155_CO5),
.O(RIOB33_X105Y161_IOB_X1Y161_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y161_IOB_X1Y162_OBUF (
.I(CLBLM_L_X12Y155_SLICE_X17Y155_DO6),
.O(RIOB33_X105Y161_IOB_X1Y162_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y163_OBUF (
.I(CLBLM_L_X12Y155_SLICE_X17Y155_DO5),
.O(RIOB33_X105Y163_IOB_X1Y163_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y163_IOB_X1Y164_OBUF (
.I(CLBLM_R_X7Y149_SLICE_X9Y149_DO5),
.O(RIOB33_X105Y163_IOB_X1Y164_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y165_OBUF (
.I(RIOB33_X105Y125_IOB_X1Y125_I),
.O(RIOB33_X105Y165_IOB_X1Y165_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y165_IOB_X1Y166_OBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_I),
.O(RIOB33_X105Y165_IOB_X1Y166_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y167_OBUF (
.I(LIOB33_SING_X0Y50_IOB_X0Y50_I),
.O(RIOB33_X105Y167_IOB_X1Y167_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y167_IOB_X1Y168_OBUF (
.I(CLBLM_L_X10Y163_SLICE_X13Y163_AO6),
.O(RIOB33_X105Y167_IOB_X1Y168_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y169_OBUF (
.I(CLBLM_R_X103Y169_SLICE_X163Y169_AO6),
.O(RIOB33_X105Y169_IOB_X1Y169_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y169_IOB_X1Y170_OBUF (
.I(CLBLM_R_X103Y169_SLICE_X163Y169_AO5),
.O(RIOB33_X105Y169_IOB_X1Y170_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y171_OBUF (
.I(CLBLM_L_X12Y159_SLICE_X16Y159_CO6),
.O(RIOB33_X105Y171_IOB_X1Y171_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y171_IOB_X1Y172_OBUF (
.I(CLBLM_R_X103Y172_SLICE_X163Y172_AO6),
.O(RIOB33_X105Y171_IOB_X1Y172_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y173_OBUF (
.I(CLBLM_R_X103Y172_SLICE_X163Y172_AO5),
.O(RIOB33_X105Y173_IOB_X1Y173_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y173_IOB_X1Y174_OBUF (
.I(CLBLM_R_X103Y174_SLICE_X163Y174_AO6),
.O(RIOB33_X105Y173_IOB_X1Y174_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y175_OBUF (
.I(CLBLM_R_X13Y157_SLICE_X18Y157_AO5),
.O(RIOB33_X105Y175_IOB_X1Y175_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y175_IOB_X1Y176_OBUF (
.I(CLBLM_R_X103Y174_SLICE_X163Y174_AO5),
.O(RIOB33_X105Y175_IOB_X1Y176_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y177_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_AO6),
.O(RIOB33_X105Y177_IOB_X1Y177_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y177_IOB_X1Y178_OBUF (
.I(CLBLM_R_X103Y177_SLICE_X163Y177_AO5),
.O(RIOB33_X105Y177_IOB_X1Y178_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y179_OBUF (
.I(CLBLM_L_X12Y159_SLICE_X16Y159_AO5),
.O(RIOB33_X105Y179_IOB_X1Y179_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y179_IOB_X1Y180_OBUF (
.I(CLBLM_R_X13Y154_SLICE_X18Y154_DO6),
.O(RIOB33_X105Y179_IOB_X1Y180_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y181_OBUF (
.I(CLBLM_R_X13Y155_SLICE_X18Y155_CO6),
.O(RIOB33_X105Y181_IOB_X1Y181_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y181_IOB_X1Y182_OBUF (
.I(CLBLM_R_X13Y155_SLICE_X18Y155_CO5),
.O(RIOB33_X105Y181_IOB_X1Y182_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y183_OBUF (
.I(CLBLM_L_X12Y155_SLICE_X17Y155_DO6),
.O(RIOB33_X105Y183_IOB_X1Y183_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y183_IOB_X1Y184_OBUF (
.I(CLBLM_L_X12Y155_SLICE_X17Y155_DO5),
.O(RIOB33_X105Y183_IOB_X1Y184_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y185_OBUF (
.I(CLBLM_R_X7Y149_SLICE_X9Y149_DO5),
.O(RIOB33_X105Y185_IOB_X1Y185_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y185_IOB_X1Y186_OBUF (
.I(CLBLM_R_X13Y154_SLICE_X18Y154_AQ),
.O(RIOB33_X105Y185_IOB_X1Y186_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y187_OBUF (
.I(CLBLM_L_X12Y155_SLICE_X16Y155_AQ),
.O(RIOB33_X105Y187_IOB_X1Y187_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y187_IOB_X1Y188_OBUF (
.I(CLBLM_R_X11Y156_SLICE_X15Y156_BQ),
.O(RIOB33_X105Y187_IOB_X1Y188_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y189_OBUF (
.I(CLBLM_L_X12Y159_SLICE_X16Y159_BQ),
.O(RIOB33_X105Y189_IOB_X1Y189_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y189_IOB_X1Y190_OBUF (
.I(CLBLM_R_X13Y156_SLICE_X18Y156_AQ),
.O(RIOB33_X105Y189_IOB_X1Y190_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y191_OBUF (
.I(CLBLM_L_X12Y156_SLICE_X16Y156_BQ),
.O(RIOB33_X105Y191_IOB_X1Y191_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y191_IOB_X1Y192_OBUF (
.I(CLBLM_R_X13Y153_SLICE_X19Y153_BQ),
.O(RIOB33_X105Y191_IOB_X1Y192_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y193_OBUF (
.I(CLBLM_L_X12Y156_SLICE_X16Y156_AQ),
.O(RIOB33_X105Y193_IOB_X1Y193_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y193_IOB_X1Y194_OBUF (
.I(CLBLM_R_X13Y156_SLICE_X19Y156_AQ),
.O(RIOB33_X105Y193_IOB_X1Y194_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y195_OBUF (
.I(CLBLM_R_X13Y157_SLICE_X18Y157_AQ),
.O(RIOB33_X105Y195_IOB_X1Y195_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y195_IOB_X1Y196_OBUF (
.I(CLBLM_L_X12Y159_SLICE_X16Y159_AQ),
.O(RIOB33_X105Y195_IOB_X1Y196_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y197_OBUF (
.I(CLBLM_L_X16Y156_SLICE_X22Y156_AO5),
.O(RIOB33_X105Y197_IOB_X1Y197_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_X105Y197_IOB_X1Y198_OBUF (
.I(CLBLM_L_X16Y156_SLICE_X22Y156_AO5),
.O(RIOB33_X105Y197_IOB_X1Y198_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y100_IOB_X1Y100_IBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_IPAD),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y149_IOB_X1Y149_IBUF (
.I(RIOB33_SING_X105Y149_IOB_X1Y149_IPAD),
.O(RIOB33_SING_X105Y149_IOB_X1Y149_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y150_IOB_X1Y150_OBUF (
.I(LIOB33_X0Y75_IOB_X0Y75_I),
.O(RIOB33_SING_X105Y150_IOB_X1Y150_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) RIOB33_SING_X105Y199_IOB_X1Y199_OBUF (
.I(CLBLM_R_X13Y156_SLICE_X19Y156_AQ),
.O(RIOB33_SING_X105Y199_IOB_X1Y199_OPAD)
  );
  assign CLBLL_L_X2Y139_SLICE_X0Y139_A = CLBLL_L_X2Y139_SLICE_X0Y139_AO6;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_B = CLBLL_L_X2Y139_SLICE_X0Y139_BO6;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_C = CLBLL_L_X2Y139_SLICE_X0Y139_CO6;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_D = CLBLL_L_X2Y139_SLICE_X0Y139_DO6;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_AMUX = CLBLL_L_X2Y139_SLICE_X0Y139_AO5;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_BMUX = CLBLL_L_X2Y139_SLICE_X0Y139_BO5;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_A = CLBLL_L_X2Y139_SLICE_X1Y139_AO6;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_B = CLBLL_L_X2Y139_SLICE_X1Y139_BO6;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_C = CLBLL_L_X2Y139_SLICE_X1Y139_CO6;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_D = CLBLL_L_X2Y139_SLICE_X1Y139_DO6;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_A = CLBLL_L_X2Y140_SLICE_X0Y140_AO6;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_B = CLBLL_L_X2Y140_SLICE_X0Y140_BO6;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_C = CLBLL_L_X2Y140_SLICE_X0Y140_CO6;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_D = CLBLL_L_X2Y140_SLICE_X0Y140_DO6;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_AMUX = CLBLL_L_X2Y140_SLICE_X0Y140_AO5;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_BMUX = CLBLL_L_X2Y140_SLICE_X0Y140_BO5;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_A = CLBLL_L_X2Y140_SLICE_X1Y140_AO6;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_B = CLBLL_L_X2Y140_SLICE_X1Y140_BO6;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_C = CLBLL_L_X2Y140_SLICE_X1Y140_CO6;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_D = CLBLL_L_X2Y140_SLICE_X1Y140_DO6;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_A = CLBLL_L_X2Y153_SLICE_X0Y153_AO6;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_B = CLBLL_L_X2Y153_SLICE_X0Y153_BO6;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_C = CLBLL_L_X2Y153_SLICE_X0Y153_CO6;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_D = CLBLL_L_X2Y153_SLICE_X0Y153_DO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_A = CLBLL_L_X2Y153_SLICE_X1Y153_AO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_B = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_C = CLBLL_L_X2Y153_SLICE_X1Y153_CO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_D = CLBLL_L_X2Y153_SLICE_X1Y153_DO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_AMUX = CLBLL_L_X2Y153_SLICE_X1Y153_AO5;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_A = CLBLL_L_X2Y154_SLICE_X0Y154_AO6;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_B = CLBLL_L_X2Y154_SLICE_X0Y154_BO6;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_C = CLBLL_L_X2Y154_SLICE_X0Y154_CO6;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_D = CLBLL_L_X2Y154_SLICE_X0Y154_DO6;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_A = CLBLL_L_X2Y154_SLICE_X1Y154_AO6;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_B = CLBLL_L_X2Y154_SLICE_X1Y154_BO6;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_C = CLBLL_L_X2Y154_SLICE_X1Y154_CO6;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_D = CLBLL_L_X2Y154_SLICE_X1Y154_DO6;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_AMUX = CLBLL_L_X2Y154_SLICE_X1Y154_AO5;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_A = CLBLL_L_X2Y155_SLICE_X0Y155_AO6;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_B = CLBLL_L_X2Y155_SLICE_X0Y155_BO6;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_C = CLBLL_L_X2Y155_SLICE_X0Y155_CO6;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_D = CLBLL_L_X2Y155_SLICE_X0Y155_DO6;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_A = CLBLL_L_X2Y155_SLICE_X1Y155_AO6;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_B = CLBLL_L_X2Y155_SLICE_X1Y155_BO6;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_C = CLBLL_L_X2Y155_SLICE_X1Y155_CO6;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_D = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_AMUX = CLBLL_L_X2Y155_SLICE_X1Y155_AO5;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_BMUX = CLBLL_L_X2Y155_SLICE_X1Y155_BO5;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_CMUX = CLBLL_L_X2Y155_SLICE_X1Y155_CO5;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A = CLBLL_L_X4Y146_SLICE_X4Y146_AO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B = CLBLL_L_X4Y146_SLICE_X4Y146_BO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C = CLBLL_L_X4Y146_SLICE_X4Y146_CO6;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D = CLBLL_L_X4Y146_SLICE_X4Y146_DO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A = CLBLL_L_X4Y146_SLICE_X5Y146_AO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B = CLBLL_L_X4Y146_SLICE_X5Y146_BO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C = CLBLL_L_X4Y146_SLICE_X5Y146_CO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D = CLBLL_L_X4Y146_SLICE_X5Y146_DO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_AMUX = CLBLL_L_X4Y146_SLICE_X5Y146_AO5;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A = CLBLL_L_X4Y147_SLICE_X4Y147_AO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B = CLBLL_L_X4Y147_SLICE_X4Y147_BO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C = CLBLL_L_X4Y147_SLICE_X4Y147_CO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D = CLBLL_L_X4Y147_SLICE_X4Y147_DO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A = CLBLL_L_X4Y147_SLICE_X5Y147_AO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B = CLBLL_L_X4Y147_SLICE_X5Y147_BO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C = CLBLL_L_X4Y147_SLICE_X5Y147_CO6;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D = CLBLL_L_X4Y147_SLICE_X5Y147_DO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A = CLBLL_L_X4Y148_SLICE_X4Y148_AO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B = CLBLL_L_X4Y148_SLICE_X4Y148_BO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C = CLBLL_L_X4Y148_SLICE_X4Y148_CO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D = CLBLL_L_X4Y148_SLICE_X4Y148_DO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_BMUX = CLBLL_L_X4Y148_SLICE_X4Y148_BO5;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A = CLBLL_L_X4Y148_SLICE_X5Y148_AO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B = CLBLL_L_X4Y148_SLICE_X5Y148_BO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C = CLBLL_L_X4Y148_SLICE_X5Y148_CO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D = CLBLL_L_X4Y148_SLICE_X5Y148_DO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A = CLBLL_L_X4Y149_SLICE_X4Y149_AO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B = CLBLL_L_X4Y149_SLICE_X4Y149_BO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C = CLBLL_L_X4Y149_SLICE_X4Y149_CO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D = CLBLL_L_X4Y149_SLICE_X4Y149_DO6;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_AMUX = CLBLL_L_X4Y149_SLICE_X4Y149_A5Q;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A = CLBLL_L_X4Y149_SLICE_X5Y149_AO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B = CLBLL_L_X4Y149_SLICE_X5Y149_BO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C = CLBLL_L_X4Y149_SLICE_X5Y149_CO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D = CLBLL_L_X4Y149_SLICE_X5Y149_DO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_AMUX = CLBLL_L_X4Y149_SLICE_X5Y149_A5Q;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_BMUX = CLBLL_L_X4Y149_SLICE_X5Y149_BO5;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_CMUX = CLBLL_L_X4Y149_SLICE_X5Y149_CO5;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_DMUX = CLBLL_L_X4Y149_SLICE_X5Y149_DO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A = CLBLL_L_X4Y150_SLICE_X4Y150_AO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B = CLBLL_L_X4Y150_SLICE_X4Y150_BO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C = CLBLL_L_X4Y150_SLICE_X4Y150_CO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A = CLBLL_L_X4Y150_SLICE_X5Y150_AO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B = CLBLL_L_X4Y150_SLICE_X5Y150_BO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C = CLBLL_L_X4Y150_SLICE_X5Y150_CO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D = CLBLL_L_X4Y150_SLICE_X5Y150_DO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_CMUX = CLBLL_L_X4Y150_SLICE_X5Y150_C5Q;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_DMUX = CLBLL_L_X4Y150_SLICE_X5Y150_D5Q;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A = CLBLL_L_X4Y151_SLICE_X4Y151_AO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B = CLBLL_L_X4Y151_SLICE_X4Y151_BO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C = CLBLL_L_X4Y151_SLICE_X4Y151_CO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D = CLBLL_L_X4Y151_SLICE_X4Y151_DO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_CMUX = CLBLL_L_X4Y151_SLICE_X4Y151_C5Q;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_DMUX = CLBLL_L_X4Y151_SLICE_X4Y151_D5Q;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A = CLBLL_L_X4Y151_SLICE_X5Y151_AO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B = CLBLL_L_X4Y151_SLICE_X5Y151_BO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C = CLBLL_L_X4Y151_SLICE_X5Y151_CO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D = CLBLL_L_X4Y151_SLICE_X5Y151_DO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A = CLBLL_L_X4Y152_SLICE_X4Y152_AO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B = CLBLL_L_X4Y152_SLICE_X4Y152_BO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C = CLBLL_L_X4Y152_SLICE_X4Y152_CO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D = CLBLL_L_X4Y152_SLICE_X4Y152_DO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A = CLBLL_L_X4Y152_SLICE_X5Y152_AO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B = CLBLL_L_X4Y152_SLICE_X5Y152_BO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C = CLBLL_L_X4Y152_SLICE_X5Y152_CO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D = CLBLL_L_X4Y152_SLICE_X5Y152_DO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_DMUX = CLBLL_L_X4Y152_SLICE_X5Y152_DO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_A = CLBLL_L_X4Y153_SLICE_X4Y153_AO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_B = CLBLL_L_X4Y153_SLICE_X4Y153_BO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_C = CLBLL_L_X4Y153_SLICE_X4Y153_CO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_D = CLBLL_L_X4Y153_SLICE_X4Y153_DO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_A = CLBLL_L_X4Y153_SLICE_X5Y153_AO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_B = CLBLL_L_X4Y153_SLICE_X5Y153_BO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_C = CLBLL_L_X4Y153_SLICE_X5Y153_CO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_D = CLBLL_L_X4Y153_SLICE_X5Y153_DO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_DMUX = CLBLL_L_X4Y153_SLICE_X5Y153_DO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_A = CLBLL_L_X4Y154_SLICE_X4Y154_AO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_B = CLBLL_L_X4Y154_SLICE_X4Y154_BO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_C = CLBLL_L_X4Y154_SLICE_X4Y154_CO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_D = CLBLL_L_X4Y154_SLICE_X4Y154_DO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_DMUX = CLBLL_L_X4Y154_SLICE_X4Y154_DO6;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_A = CLBLL_L_X4Y154_SLICE_X5Y154_AO6;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_B = CLBLL_L_X4Y154_SLICE_X5Y154_BO6;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_C = CLBLL_L_X4Y154_SLICE_X5Y154_CO6;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_D = CLBLL_L_X4Y154_SLICE_X5Y154_DO6;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_A = CLBLL_L_X4Y155_SLICE_X4Y155_AO6;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_B = CLBLL_L_X4Y155_SLICE_X4Y155_BO6;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_C = CLBLL_L_X4Y155_SLICE_X4Y155_CO6;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_D = CLBLL_L_X4Y155_SLICE_X4Y155_DO6;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_A = CLBLL_L_X4Y155_SLICE_X5Y155_AO6;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_B = CLBLL_L_X4Y155_SLICE_X5Y155_BO6;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_C = CLBLL_L_X4Y155_SLICE_X5Y155_CO6;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_D = CLBLL_L_X4Y155_SLICE_X5Y155_DO6;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_AMUX = CLBLL_L_X4Y155_SLICE_X5Y155_A5Q;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_A = CLBLL_L_X4Y156_SLICE_X4Y156_AO6;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_B = CLBLL_L_X4Y156_SLICE_X4Y156_BO6;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_C = CLBLL_L_X4Y156_SLICE_X4Y156_CO6;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_D = CLBLL_L_X4Y156_SLICE_X4Y156_DO6;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_AMUX = CLBLL_L_X4Y156_SLICE_X4Y156_AO5;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_BMUX = CLBLL_L_X4Y156_SLICE_X4Y156_BO5;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_CMUX = CLBLL_L_X4Y156_SLICE_X4Y156_CO5;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_A = CLBLL_L_X4Y156_SLICE_X5Y156_AO6;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_B = CLBLL_L_X4Y156_SLICE_X5Y156_BO6;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_C = CLBLL_L_X4Y156_SLICE_X5Y156_CO6;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_D = CLBLL_L_X4Y156_SLICE_X5Y156_DO6;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_CMUX = CLBLL_L_X4Y156_SLICE_X5Y156_CO6;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_DMUX = CLBLL_L_X4Y156_SLICE_X5Y156_DO6;
  assign CLBLL_L_X4Y157_SLICE_X4Y157_A = CLBLL_L_X4Y157_SLICE_X4Y157_AO6;
  assign CLBLL_L_X4Y157_SLICE_X4Y157_B = CLBLL_L_X4Y157_SLICE_X4Y157_BO6;
  assign CLBLL_L_X4Y157_SLICE_X4Y157_C = CLBLL_L_X4Y157_SLICE_X4Y157_CO6;
  assign CLBLL_L_X4Y157_SLICE_X4Y157_D = CLBLL_L_X4Y157_SLICE_X4Y157_DO6;
  assign CLBLL_L_X4Y157_SLICE_X4Y157_AMUX = CLBLL_L_X4Y157_SLICE_X4Y157_AO5;
  assign CLBLL_L_X4Y157_SLICE_X4Y157_BMUX = CLBLL_L_X4Y157_SLICE_X4Y157_BO5;
  assign CLBLL_L_X4Y157_SLICE_X4Y157_CMUX = CLBLL_L_X4Y157_SLICE_X4Y157_CO5;
  assign CLBLL_L_X4Y157_SLICE_X5Y157_A = CLBLL_L_X4Y157_SLICE_X5Y157_AO6;
  assign CLBLL_L_X4Y157_SLICE_X5Y157_B = CLBLL_L_X4Y157_SLICE_X5Y157_BO6;
  assign CLBLL_L_X4Y157_SLICE_X5Y157_C = CLBLL_L_X4Y157_SLICE_X5Y157_CO6;
  assign CLBLL_L_X4Y157_SLICE_X5Y157_D = CLBLL_L_X4Y157_SLICE_X5Y157_DO6;
  assign CLBLL_L_X4Y157_SLICE_X5Y157_AMUX = CLBLL_L_X4Y157_SLICE_X5Y157_AO5;
  assign CLBLL_L_X4Y158_SLICE_X4Y158_A = CLBLL_L_X4Y158_SLICE_X4Y158_AO6;
  assign CLBLL_L_X4Y158_SLICE_X4Y158_B = CLBLL_L_X4Y158_SLICE_X4Y158_BO6;
  assign CLBLL_L_X4Y158_SLICE_X4Y158_C = CLBLL_L_X4Y158_SLICE_X4Y158_CO6;
  assign CLBLL_L_X4Y158_SLICE_X4Y158_D = CLBLL_L_X4Y158_SLICE_X4Y158_DO6;
  assign CLBLL_L_X4Y158_SLICE_X5Y158_A = CLBLL_L_X4Y158_SLICE_X5Y158_AO6;
  assign CLBLL_L_X4Y158_SLICE_X5Y158_B = CLBLL_L_X4Y158_SLICE_X5Y158_BO6;
  assign CLBLL_L_X4Y158_SLICE_X5Y158_C = CLBLL_L_X4Y158_SLICE_X5Y158_CO6;
  assign CLBLL_L_X4Y158_SLICE_X5Y158_D = CLBLL_L_X4Y158_SLICE_X5Y158_DO6;
  assign CLBLL_L_X36Y150_SLICE_X54Y150_A = CLBLL_L_X36Y150_SLICE_X54Y150_AO6;
  assign CLBLL_L_X36Y150_SLICE_X54Y150_B = CLBLL_L_X36Y150_SLICE_X54Y150_BO6;
  assign CLBLL_L_X36Y150_SLICE_X54Y150_C = CLBLL_L_X36Y150_SLICE_X54Y150_CO6;
  assign CLBLL_L_X36Y150_SLICE_X54Y150_D = CLBLL_L_X36Y150_SLICE_X54Y150_DO6;
  assign CLBLL_L_X36Y150_SLICE_X55Y150_A = CLBLL_L_X36Y150_SLICE_X55Y150_AO6;
  assign CLBLL_L_X36Y150_SLICE_X55Y150_B = CLBLL_L_X36Y150_SLICE_X55Y150_BO6;
  assign CLBLL_L_X36Y150_SLICE_X55Y150_C = CLBLL_L_X36Y150_SLICE_X55Y150_CO6;
  assign CLBLL_L_X36Y150_SLICE_X55Y150_D = CLBLL_L_X36Y150_SLICE_X55Y150_DO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B = CLBLL_L_X52Y126_SLICE_X78Y126_BO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C = CLBLL_L_X52Y126_SLICE_X78Y126_CO6;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D = CLBLL_L_X52Y126_SLICE_X78Y126_DO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A = CLBLL_L_X52Y126_SLICE_X79Y126_AO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B = CLBLL_L_X52Y126_SLICE_X79Y126_BO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C = CLBLL_L_X52Y126_SLICE_X79Y126_CO6;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D = CLBLL_L_X52Y126_SLICE_X79Y126_DO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A = CLBLM_L_X8Y146_SLICE_X10Y146_AO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B = CLBLM_L_X8Y146_SLICE_X10Y146_BO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C = CLBLM_L_X8Y146_SLICE_X10Y146_CO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D = CLBLM_L_X8Y146_SLICE_X10Y146_DO6;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_BMUX = CLBLM_L_X8Y146_SLICE_X10Y146_B5Q;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A = CLBLM_L_X8Y146_SLICE_X11Y146_AO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B = CLBLM_L_X8Y146_SLICE_X11Y146_BO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C = CLBLM_L_X8Y146_SLICE_X11Y146_CO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D = CLBLM_L_X8Y146_SLICE_X11Y146_DO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A = CLBLM_L_X8Y147_SLICE_X10Y147_AO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B = CLBLM_L_X8Y147_SLICE_X10Y147_BO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C = CLBLM_L_X8Y147_SLICE_X10Y147_CO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D = CLBLM_L_X8Y147_SLICE_X10Y147_DO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_AMUX = CLBLM_L_X8Y147_SLICE_X10Y147_AO5;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_DMUX = CLBLM_L_X8Y147_SLICE_X10Y147_DO5;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A = CLBLM_L_X8Y147_SLICE_X11Y147_AO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B = CLBLM_L_X8Y147_SLICE_X11Y147_BO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C = CLBLM_L_X8Y147_SLICE_X11Y147_CO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D = CLBLM_L_X8Y147_SLICE_X11Y147_DO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A = CLBLM_L_X8Y148_SLICE_X10Y148_AO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B = CLBLM_L_X8Y148_SLICE_X10Y148_BO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C = CLBLM_L_X8Y148_SLICE_X10Y148_CO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D = CLBLM_L_X8Y148_SLICE_X10Y148_DO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A = CLBLM_L_X8Y148_SLICE_X11Y148_AO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B = CLBLM_L_X8Y148_SLICE_X11Y148_BO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C = CLBLM_L_X8Y148_SLICE_X11Y148_CO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D = CLBLM_L_X8Y148_SLICE_X11Y148_DO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_AMUX = CLBLM_L_X8Y148_SLICE_X11Y148_A5Q;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_BMUX = CLBLM_L_X8Y148_SLICE_X11Y148_B5Q;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_CMUX = CLBLM_L_X8Y148_SLICE_X11Y148_CO5;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_DMUX = CLBLM_L_X8Y148_SLICE_X11Y148_DO5;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A = CLBLM_L_X8Y149_SLICE_X10Y149_AO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B = CLBLM_L_X8Y149_SLICE_X10Y149_BO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C = CLBLM_L_X8Y149_SLICE_X10Y149_CO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D = CLBLM_L_X8Y149_SLICE_X10Y149_DO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_BMUX = CLBLM_L_X8Y149_SLICE_X10Y149_BO5;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A = CLBLM_L_X8Y149_SLICE_X11Y149_AO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B = CLBLM_L_X8Y149_SLICE_X11Y149_BO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C = CLBLM_L_X8Y149_SLICE_X11Y149_CO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D = CLBLM_L_X8Y149_SLICE_X11Y149_DO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A = CLBLM_L_X8Y150_SLICE_X10Y150_AO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B = CLBLM_L_X8Y150_SLICE_X10Y150_BO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C = CLBLM_L_X8Y150_SLICE_X10Y150_CO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D = CLBLM_L_X8Y150_SLICE_X10Y150_DO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_AMUX = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_CMUX = CLBLM_L_X8Y150_SLICE_X10Y150_CO5;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A = CLBLM_L_X8Y150_SLICE_X11Y150_AO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B = CLBLM_L_X8Y150_SLICE_X11Y150_BO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C = CLBLM_L_X8Y150_SLICE_X11Y150_CO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D = CLBLM_L_X8Y150_SLICE_X11Y150_DO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A = CLBLM_L_X8Y151_SLICE_X10Y151_AO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B = CLBLM_L_X8Y151_SLICE_X10Y151_BO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C = CLBLM_L_X8Y151_SLICE_X10Y151_CO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D = CLBLM_L_X8Y151_SLICE_X10Y151_DO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A = CLBLM_L_X8Y151_SLICE_X11Y151_AO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B = CLBLM_L_X8Y151_SLICE_X11Y151_BO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C = CLBLM_L_X8Y151_SLICE_X11Y151_CO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D = CLBLM_L_X8Y151_SLICE_X11Y151_DO6;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_A = CLBLM_L_X8Y152_SLICE_X10Y152_AO6;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_B = CLBLM_L_X8Y152_SLICE_X10Y152_BO6;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_C = CLBLM_L_X8Y152_SLICE_X10Y152_CO6;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_D = CLBLM_L_X8Y152_SLICE_X10Y152_DO6;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_A = CLBLM_L_X8Y152_SLICE_X11Y152_AO6;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_B = CLBLM_L_X8Y152_SLICE_X11Y152_BO6;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_C = CLBLM_L_X8Y152_SLICE_X11Y152_CO6;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_D = CLBLM_L_X8Y152_SLICE_X11Y152_DO6;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_AMUX = CLBLM_L_X8Y152_SLICE_X11Y152_AO5;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_BMUX = CLBLM_L_X8Y152_SLICE_X11Y152_BO5;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_A = CLBLM_L_X8Y153_SLICE_X10Y153_AO6;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_B = CLBLM_L_X8Y153_SLICE_X10Y153_BO6;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_C = CLBLM_L_X8Y153_SLICE_X10Y153_CO6;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_D = CLBLM_L_X8Y153_SLICE_X10Y153_DO6;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_AMUX = CLBLM_L_X8Y153_SLICE_X10Y153_A5Q;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_A = CLBLM_L_X8Y153_SLICE_X11Y153_AO6;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_B = CLBLM_L_X8Y153_SLICE_X11Y153_BO6;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_C = CLBLM_L_X8Y153_SLICE_X11Y153_CO6;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_D = CLBLM_L_X8Y153_SLICE_X11Y153_DO6;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_CMUX = CLBLM_L_X8Y153_SLICE_X11Y153_C5Q;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_A = CLBLM_L_X8Y154_SLICE_X10Y154_AO6;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_B = CLBLM_L_X8Y154_SLICE_X10Y154_BO6;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_C = CLBLM_L_X8Y154_SLICE_X10Y154_CO6;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_D = CLBLM_L_X8Y154_SLICE_X10Y154_DO6;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_AMUX = CLBLM_L_X8Y154_SLICE_X10Y154_A5Q;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_BMUX = CLBLM_L_X8Y154_SLICE_X10Y154_B5Q;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_CMUX = CLBLM_L_X8Y154_SLICE_X10Y154_C5Q;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_A = CLBLM_L_X8Y154_SLICE_X11Y154_AO6;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_B = CLBLM_L_X8Y154_SLICE_X11Y154_BO6;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_C = CLBLM_L_X8Y154_SLICE_X11Y154_CO6;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_D = CLBLM_L_X8Y154_SLICE_X11Y154_DO6;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_AMUX = CLBLM_L_X8Y154_SLICE_X11Y154_A5Q;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_A = CLBLM_L_X8Y155_SLICE_X10Y155_AO6;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_B = CLBLM_L_X8Y155_SLICE_X10Y155_BO6;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_C = CLBLM_L_X8Y155_SLICE_X10Y155_CO6;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_D = CLBLM_L_X8Y155_SLICE_X10Y155_DO6;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_BMUX = CLBLM_L_X8Y155_SLICE_X10Y155_B5Q;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_A = CLBLM_L_X8Y155_SLICE_X11Y155_AO6;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_B = CLBLM_L_X8Y155_SLICE_X11Y155_BO6;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_C = CLBLM_L_X8Y155_SLICE_X11Y155_CO6;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_D = CLBLM_L_X8Y155_SLICE_X11Y155_DO6;
  assign CLBLM_L_X8Y156_SLICE_X10Y156_A = CLBLM_L_X8Y156_SLICE_X10Y156_AO6;
  assign CLBLM_L_X8Y156_SLICE_X10Y156_B = CLBLM_L_X8Y156_SLICE_X10Y156_BO6;
  assign CLBLM_L_X8Y156_SLICE_X10Y156_C = CLBLM_L_X8Y156_SLICE_X10Y156_CO6;
  assign CLBLM_L_X8Y156_SLICE_X10Y156_D = CLBLM_L_X8Y156_SLICE_X10Y156_DO6;
  assign CLBLM_L_X8Y156_SLICE_X11Y156_A = CLBLM_L_X8Y156_SLICE_X11Y156_AO6;
  assign CLBLM_L_X8Y156_SLICE_X11Y156_B = CLBLM_L_X8Y156_SLICE_X11Y156_BO6;
  assign CLBLM_L_X8Y156_SLICE_X11Y156_C = CLBLM_L_X8Y156_SLICE_X11Y156_CO6;
  assign CLBLM_L_X8Y156_SLICE_X11Y156_D = CLBLM_L_X8Y156_SLICE_X11Y156_DO6;
  assign CLBLM_L_X8Y156_SLICE_X11Y156_BMUX = CLBLM_L_X8Y156_SLICE_X11Y156_B5Q;
  assign CLBLM_L_X8Y157_SLICE_X10Y157_A = CLBLM_L_X8Y157_SLICE_X10Y157_AO6;
  assign CLBLM_L_X8Y157_SLICE_X10Y157_B = CLBLM_L_X8Y157_SLICE_X10Y157_BO6;
  assign CLBLM_L_X8Y157_SLICE_X10Y157_C = CLBLM_L_X8Y157_SLICE_X10Y157_CO6;
  assign CLBLM_L_X8Y157_SLICE_X10Y157_D = CLBLM_L_X8Y157_SLICE_X10Y157_DO6;
  assign CLBLM_L_X8Y157_SLICE_X11Y157_A = CLBLM_L_X8Y157_SLICE_X11Y157_AO6;
  assign CLBLM_L_X8Y157_SLICE_X11Y157_B = CLBLM_L_X8Y157_SLICE_X11Y157_BO6;
  assign CLBLM_L_X8Y157_SLICE_X11Y157_C = CLBLM_L_X8Y157_SLICE_X11Y157_CO6;
  assign CLBLM_L_X8Y157_SLICE_X11Y157_D = CLBLM_L_X8Y157_SLICE_X11Y157_DO6;
  assign CLBLM_L_X8Y158_SLICE_X10Y158_A = CLBLM_L_X8Y158_SLICE_X10Y158_AO6;
  assign CLBLM_L_X8Y158_SLICE_X10Y158_B = CLBLM_L_X8Y158_SLICE_X10Y158_BO6;
  assign CLBLM_L_X8Y158_SLICE_X10Y158_C = CLBLM_L_X8Y158_SLICE_X10Y158_CO6;
  assign CLBLM_L_X8Y158_SLICE_X10Y158_D = CLBLM_L_X8Y158_SLICE_X10Y158_DO6;
  assign CLBLM_L_X8Y158_SLICE_X11Y158_A = CLBLM_L_X8Y158_SLICE_X11Y158_AO6;
  assign CLBLM_L_X8Y158_SLICE_X11Y158_B = CLBLM_L_X8Y158_SLICE_X11Y158_BO6;
  assign CLBLM_L_X8Y158_SLICE_X11Y158_C = CLBLM_L_X8Y158_SLICE_X11Y158_CO6;
  assign CLBLM_L_X8Y158_SLICE_X11Y158_D = CLBLM_L_X8Y158_SLICE_X11Y158_DO6;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_A = CLBLM_L_X8Y159_SLICE_X10Y159_AO6;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_B = CLBLM_L_X8Y159_SLICE_X10Y159_BO6;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_C = CLBLM_L_X8Y159_SLICE_X10Y159_CO6;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_D = CLBLM_L_X8Y159_SLICE_X10Y159_DO6;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_BMUX = CLBLM_L_X8Y159_SLICE_X10Y159_BO5;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_A = CLBLM_L_X8Y159_SLICE_X11Y159_AO6;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_B = CLBLM_L_X8Y159_SLICE_X11Y159_BO6;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_C = CLBLM_L_X8Y159_SLICE_X11Y159_CO6;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_D = CLBLM_L_X8Y159_SLICE_X11Y159_DO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A = CLBLM_L_X10Y144_SLICE_X12Y144_AO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B = CLBLM_L_X10Y144_SLICE_X12Y144_BO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C = CLBLM_L_X10Y144_SLICE_X12Y144_CO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D = CLBLM_L_X10Y144_SLICE_X12Y144_DO6;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_AMUX = CLBLM_L_X10Y144_SLICE_X12Y144_AO5;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A = CLBLM_L_X10Y144_SLICE_X13Y144_AO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B = CLBLM_L_X10Y144_SLICE_X13Y144_BO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C = CLBLM_L_X10Y144_SLICE_X13Y144_CO6;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D = CLBLM_L_X10Y144_SLICE_X13Y144_DO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A = CLBLM_L_X10Y145_SLICE_X12Y145_AO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B = CLBLM_L_X10Y145_SLICE_X12Y145_BO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C = CLBLM_L_X10Y145_SLICE_X12Y145_CO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D = CLBLM_L_X10Y145_SLICE_X12Y145_DO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A = CLBLM_L_X10Y145_SLICE_X13Y145_AO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B = CLBLM_L_X10Y145_SLICE_X13Y145_BO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C = CLBLM_L_X10Y145_SLICE_X13Y145_CO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D = CLBLM_L_X10Y145_SLICE_X13Y145_DO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_DMUX = CLBLM_L_X10Y145_SLICE_X13Y145_DO5;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A = CLBLM_L_X10Y146_SLICE_X12Y146_AO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B = CLBLM_L_X10Y146_SLICE_X12Y146_BO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C = CLBLM_L_X10Y146_SLICE_X12Y146_CO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D = CLBLM_L_X10Y146_SLICE_X12Y146_DO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_CMUX = CLBLM_L_X10Y146_SLICE_X12Y146_C5Q;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A = CLBLM_L_X10Y146_SLICE_X13Y146_AO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B = CLBLM_L_X10Y146_SLICE_X13Y146_BO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C = CLBLM_L_X10Y146_SLICE_X13Y146_CO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_BMUX = CLBLM_L_X10Y146_SLICE_X13Y146_BO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A = CLBLM_L_X10Y147_SLICE_X12Y147_AO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B = CLBLM_L_X10Y147_SLICE_X12Y147_BO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C = CLBLM_L_X10Y147_SLICE_X12Y147_CO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D = CLBLM_L_X10Y147_SLICE_X12Y147_DO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A = CLBLM_L_X10Y147_SLICE_X13Y147_AO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B = CLBLM_L_X10Y147_SLICE_X13Y147_BO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C = CLBLM_L_X10Y147_SLICE_X13Y147_CO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D = CLBLM_L_X10Y147_SLICE_X13Y147_DO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_DMUX = CLBLM_L_X10Y147_SLICE_X13Y147_DO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A = CLBLM_L_X10Y148_SLICE_X12Y148_AO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B = CLBLM_L_X10Y148_SLICE_X12Y148_BO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C = CLBLM_L_X10Y148_SLICE_X12Y148_CO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D = CLBLM_L_X10Y148_SLICE_X12Y148_DO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_BMUX = CLBLM_L_X10Y148_SLICE_X12Y148_BO5;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_CMUX = CLBLM_L_X10Y148_SLICE_X12Y148_CO5;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A = CLBLM_L_X10Y148_SLICE_X13Y148_AO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B = CLBLM_L_X10Y148_SLICE_X13Y148_BO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C = CLBLM_L_X10Y148_SLICE_X13Y148_CO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D = CLBLM_L_X10Y148_SLICE_X13Y148_DO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A = CLBLM_L_X10Y149_SLICE_X12Y149_AO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B = CLBLM_L_X10Y149_SLICE_X12Y149_BO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C = CLBLM_L_X10Y149_SLICE_X12Y149_CO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D = CLBLM_L_X10Y149_SLICE_X12Y149_DO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_CMUX = CLBLM_L_X10Y149_SLICE_X12Y149_C5Q;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_DMUX = CLBLM_L_X10Y149_SLICE_X12Y149_DO5;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A = CLBLM_L_X10Y149_SLICE_X13Y149_AO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B = CLBLM_L_X10Y149_SLICE_X13Y149_BO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C = CLBLM_L_X10Y149_SLICE_X13Y149_CO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D = CLBLM_L_X10Y149_SLICE_X13Y149_DO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_AMUX = CLBLM_L_X10Y149_SLICE_X13Y149_A5Q;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_BMUX = CLBLM_L_X10Y149_SLICE_X13Y149_BO5;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_CMUX = CLBLM_L_X10Y149_SLICE_X13Y149_CO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A = CLBLM_L_X10Y150_SLICE_X12Y150_AO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B = CLBLM_L_X10Y150_SLICE_X12Y150_BO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C = CLBLM_L_X10Y150_SLICE_X12Y150_CO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D = CLBLM_L_X10Y150_SLICE_X12Y150_DO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_AMUX = CLBLM_L_X10Y150_SLICE_X12Y150_A5Q;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_BMUX = CLBLM_L_X10Y150_SLICE_X12Y150_BO5;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A = CLBLM_L_X10Y150_SLICE_X13Y150_AO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B = CLBLM_L_X10Y150_SLICE_X13Y150_BO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C = CLBLM_L_X10Y150_SLICE_X13Y150_CO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D = CLBLM_L_X10Y150_SLICE_X13Y150_DO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_BMUX = CLBLM_L_X10Y150_SLICE_X13Y150_B5Q;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_CMUX = CLBLM_L_X10Y150_SLICE_X13Y150_C5Q;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A = CLBLM_L_X10Y151_SLICE_X12Y151_AO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B = CLBLM_L_X10Y151_SLICE_X12Y151_BO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C = CLBLM_L_X10Y151_SLICE_X12Y151_CO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D = CLBLM_L_X10Y151_SLICE_X12Y151_DO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A = CLBLM_L_X10Y151_SLICE_X13Y151_AO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B = CLBLM_L_X10Y151_SLICE_X13Y151_BO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C = CLBLM_L_X10Y151_SLICE_X13Y151_CO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D = CLBLM_L_X10Y151_SLICE_X13Y151_DO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_BMUX = CLBLM_L_X10Y151_SLICE_X13Y151_B5Q;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A = CLBLM_L_X10Y152_SLICE_X12Y152_AO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B = CLBLM_L_X10Y152_SLICE_X12Y152_BO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C = CLBLM_L_X10Y152_SLICE_X12Y152_CO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D = CLBLM_L_X10Y152_SLICE_X12Y152_DO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_CMUX = CLBLM_L_X10Y152_SLICE_X12Y152_CO5;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A = CLBLM_L_X10Y152_SLICE_X13Y152_AO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B = CLBLM_L_X10Y152_SLICE_X13Y152_BO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C = CLBLM_L_X10Y152_SLICE_X13Y152_CO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D = CLBLM_L_X10Y152_SLICE_X13Y152_DO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_BMUX = CLBLM_L_X10Y152_SLICE_X13Y152_BO5;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_CMUX = CLBLM_L_X10Y152_SLICE_X13Y152_CO5;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A = CLBLM_L_X10Y153_SLICE_X12Y153_AO6;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B = CLBLM_L_X10Y153_SLICE_X12Y153_BO6;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C = CLBLM_L_X10Y153_SLICE_X12Y153_CO6;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D = CLBLM_L_X10Y153_SLICE_X12Y153_DO6;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A = CLBLM_L_X10Y153_SLICE_X13Y153_AO6;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B = CLBLM_L_X10Y153_SLICE_X13Y153_BO6;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C = CLBLM_L_X10Y153_SLICE_X13Y153_CO6;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D = CLBLM_L_X10Y153_SLICE_X13Y153_DO6;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_BMUX = CLBLM_L_X10Y153_SLICE_X13Y153_BO5;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_A = CLBLM_L_X10Y154_SLICE_X12Y154_AO6;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_B = CLBLM_L_X10Y154_SLICE_X12Y154_BO6;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_C = CLBLM_L_X10Y154_SLICE_X12Y154_CO6;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_D = CLBLM_L_X10Y154_SLICE_X12Y154_DO6;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_AMUX = CLBLM_L_X10Y154_SLICE_X12Y154_A5Q;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_BMUX = CLBLM_L_X10Y154_SLICE_X12Y154_BO5;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_A = CLBLM_L_X10Y154_SLICE_X13Y154_AO6;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_B = CLBLM_L_X10Y154_SLICE_X13Y154_BO6;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_C = CLBLM_L_X10Y154_SLICE_X13Y154_CO6;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_D = CLBLM_L_X10Y154_SLICE_X13Y154_DO6;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_AMUX = CLBLM_L_X10Y154_SLICE_X13Y154_AO5;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_CMUX = CLBLM_L_X10Y154_SLICE_X13Y154_C5Q;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_A = CLBLM_L_X10Y155_SLICE_X12Y155_AO6;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_B = CLBLM_L_X10Y155_SLICE_X12Y155_BO6;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_C = CLBLM_L_X10Y155_SLICE_X12Y155_CO6;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_D = CLBLM_L_X10Y155_SLICE_X12Y155_DO6;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_A = CLBLM_L_X10Y155_SLICE_X13Y155_AO6;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_B = CLBLM_L_X10Y155_SLICE_X13Y155_BO6;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_C = CLBLM_L_X10Y155_SLICE_X13Y155_CO6;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_D = CLBLM_L_X10Y155_SLICE_X13Y155_DO6;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_AMUX = CLBLM_L_X10Y155_SLICE_X13Y155_A5Q;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_DMUX = CLBLM_L_X10Y155_SLICE_X13Y155_DO6;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_A = CLBLM_L_X10Y156_SLICE_X12Y156_AO6;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_B = CLBLM_L_X10Y156_SLICE_X12Y156_BO6;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_C = CLBLM_L_X10Y156_SLICE_X12Y156_CO6;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_D = CLBLM_L_X10Y156_SLICE_X12Y156_DO6;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_CMUX = CLBLM_L_X10Y156_SLICE_X12Y156_CO6;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_A = CLBLM_L_X10Y156_SLICE_X13Y156_AO6;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_B = CLBLM_L_X10Y156_SLICE_X13Y156_BO6;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_C = CLBLM_L_X10Y156_SLICE_X13Y156_CO6;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_D = CLBLM_L_X10Y156_SLICE_X13Y156_DO6;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_AMUX = CLBLM_L_X10Y156_SLICE_X13Y156_AO5;
  assign CLBLM_L_X10Y157_SLICE_X12Y157_A = CLBLM_L_X10Y157_SLICE_X12Y157_AO6;
  assign CLBLM_L_X10Y157_SLICE_X12Y157_B = CLBLM_L_X10Y157_SLICE_X12Y157_BO6;
  assign CLBLM_L_X10Y157_SLICE_X12Y157_C = CLBLM_L_X10Y157_SLICE_X12Y157_CO6;
  assign CLBLM_L_X10Y157_SLICE_X12Y157_D = CLBLM_L_X10Y157_SLICE_X12Y157_DO6;
  assign CLBLM_L_X10Y157_SLICE_X12Y157_CMUX = CLBLM_L_X10Y157_SLICE_X12Y157_CO5;
  assign CLBLM_L_X10Y157_SLICE_X13Y157_A = CLBLM_L_X10Y157_SLICE_X13Y157_AO6;
  assign CLBLM_L_X10Y157_SLICE_X13Y157_B = CLBLM_L_X10Y157_SLICE_X13Y157_BO6;
  assign CLBLM_L_X10Y157_SLICE_X13Y157_C = CLBLM_L_X10Y157_SLICE_X13Y157_CO6;
  assign CLBLM_L_X10Y157_SLICE_X13Y157_D = CLBLM_L_X10Y157_SLICE_X13Y157_DO6;
  assign CLBLM_L_X10Y157_SLICE_X13Y157_AMUX = CLBLM_L_X10Y157_SLICE_X13Y157_AO5;
  assign CLBLM_L_X10Y158_SLICE_X12Y158_A = CLBLM_L_X10Y158_SLICE_X12Y158_AO6;
  assign CLBLM_L_X10Y158_SLICE_X12Y158_B = CLBLM_L_X10Y158_SLICE_X12Y158_BO6;
  assign CLBLM_L_X10Y158_SLICE_X12Y158_C = CLBLM_L_X10Y158_SLICE_X12Y158_CO6;
  assign CLBLM_L_X10Y158_SLICE_X12Y158_D = CLBLM_L_X10Y158_SLICE_X12Y158_DO6;
  assign CLBLM_L_X10Y158_SLICE_X13Y158_A = CLBLM_L_X10Y158_SLICE_X13Y158_AO6;
  assign CLBLM_L_X10Y158_SLICE_X13Y158_B = CLBLM_L_X10Y158_SLICE_X13Y158_BO6;
  assign CLBLM_L_X10Y158_SLICE_X13Y158_C = CLBLM_L_X10Y158_SLICE_X13Y158_CO6;
  assign CLBLM_L_X10Y158_SLICE_X13Y158_D = CLBLM_L_X10Y158_SLICE_X13Y158_DO6;
  assign CLBLM_L_X10Y159_SLICE_X12Y159_A = CLBLM_L_X10Y159_SLICE_X12Y159_AO6;
  assign CLBLM_L_X10Y159_SLICE_X12Y159_B = CLBLM_L_X10Y159_SLICE_X12Y159_BO6;
  assign CLBLM_L_X10Y159_SLICE_X12Y159_C = CLBLM_L_X10Y159_SLICE_X12Y159_CO6;
  assign CLBLM_L_X10Y159_SLICE_X12Y159_D = CLBLM_L_X10Y159_SLICE_X12Y159_DO6;
  assign CLBLM_L_X10Y159_SLICE_X13Y159_A = CLBLM_L_X10Y159_SLICE_X13Y159_AO6;
  assign CLBLM_L_X10Y159_SLICE_X13Y159_B = CLBLM_L_X10Y159_SLICE_X13Y159_BO6;
  assign CLBLM_L_X10Y159_SLICE_X13Y159_C = CLBLM_L_X10Y159_SLICE_X13Y159_CO6;
  assign CLBLM_L_X10Y159_SLICE_X13Y159_D = CLBLM_L_X10Y159_SLICE_X13Y159_DO6;
  assign CLBLM_L_X10Y159_SLICE_X13Y159_AMUX = CLBLM_L_X10Y159_SLICE_X13Y159_AO5;
  assign CLBLM_L_X10Y159_SLICE_X13Y159_BMUX = CLBLM_L_X10Y159_SLICE_X13Y159_BO5;
  assign CLBLM_L_X10Y163_SLICE_X12Y163_A = CLBLM_L_X10Y163_SLICE_X12Y163_AO6;
  assign CLBLM_L_X10Y163_SLICE_X12Y163_B = CLBLM_L_X10Y163_SLICE_X12Y163_BO6;
  assign CLBLM_L_X10Y163_SLICE_X12Y163_C = CLBLM_L_X10Y163_SLICE_X12Y163_CO6;
  assign CLBLM_L_X10Y163_SLICE_X12Y163_D = CLBLM_L_X10Y163_SLICE_X12Y163_DO6;
  assign CLBLM_L_X10Y163_SLICE_X13Y163_A = CLBLM_L_X10Y163_SLICE_X13Y163_AO6;
  assign CLBLM_L_X10Y163_SLICE_X13Y163_B = CLBLM_L_X10Y163_SLICE_X13Y163_BO6;
  assign CLBLM_L_X10Y163_SLICE_X13Y163_C = CLBLM_L_X10Y163_SLICE_X13Y163_CO6;
  assign CLBLM_L_X10Y163_SLICE_X13Y163_D = CLBLM_L_X10Y163_SLICE_X13Y163_DO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A = CLBLM_L_X12Y146_SLICE_X16Y146_AO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B = CLBLM_L_X12Y146_SLICE_X16Y146_BO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C = CLBLM_L_X12Y146_SLICE_X16Y146_CO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D = CLBLM_L_X12Y146_SLICE_X16Y146_DO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A = CLBLM_L_X12Y146_SLICE_X17Y146_AO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B = CLBLM_L_X12Y146_SLICE_X17Y146_BO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C = CLBLM_L_X12Y146_SLICE_X17Y146_CO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D = CLBLM_L_X12Y146_SLICE_X17Y146_DO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A = CLBLM_L_X12Y147_SLICE_X16Y147_AO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B = CLBLM_L_X12Y147_SLICE_X16Y147_BO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C = CLBLM_L_X12Y147_SLICE_X16Y147_CO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_BMUX = CLBLM_L_X12Y147_SLICE_X16Y147_BO5;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A = CLBLM_L_X12Y147_SLICE_X17Y147_AO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B = CLBLM_L_X12Y147_SLICE_X17Y147_BO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C = CLBLM_L_X12Y147_SLICE_X17Y147_CO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D = CLBLM_L_X12Y147_SLICE_X17Y147_DO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A = CLBLM_L_X12Y148_SLICE_X16Y148_AO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B = CLBLM_L_X12Y148_SLICE_X16Y148_BO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C = CLBLM_L_X12Y148_SLICE_X16Y148_CO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D = CLBLM_L_X12Y148_SLICE_X16Y148_DO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_AMUX = CLBLM_L_X12Y148_SLICE_X16Y148_AO5;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A = CLBLM_L_X12Y148_SLICE_X17Y148_AO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B = CLBLM_L_X12Y148_SLICE_X17Y148_BO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C = CLBLM_L_X12Y148_SLICE_X17Y148_CO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D = CLBLM_L_X12Y148_SLICE_X17Y148_DO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_DMUX = CLBLM_L_X12Y148_SLICE_X17Y148_DO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A = CLBLM_L_X12Y149_SLICE_X16Y149_AO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B = CLBLM_L_X12Y149_SLICE_X16Y149_BO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C = CLBLM_L_X12Y149_SLICE_X16Y149_CO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D = CLBLM_L_X12Y149_SLICE_X16Y149_DO6;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_BMUX = CLBLM_L_X12Y149_SLICE_X16Y149_B5Q;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A = CLBLM_L_X12Y149_SLICE_X17Y149_AO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B = CLBLM_L_X12Y149_SLICE_X17Y149_BO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C = CLBLM_L_X12Y149_SLICE_X17Y149_CO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D = CLBLM_L_X12Y149_SLICE_X17Y149_DO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_AMUX = CLBLM_L_X12Y149_SLICE_X17Y149_A5Q;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_BMUX = CLBLM_L_X12Y149_SLICE_X17Y149_BO5;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_CMUX = CLBLM_L_X12Y149_SLICE_X17Y149_CO5;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_DMUX = CLBLM_L_X12Y149_SLICE_X17Y149_DO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A = CLBLM_L_X12Y150_SLICE_X16Y150_AO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B = CLBLM_L_X12Y150_SLICE_X16Y150_BO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C = CLBLM_L_X12Y150_SLICE_X16Y150_CO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D = CLBLM_L_X12Y150_SLICE_X16Y150_DO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_AMUX = CLBLM_L_X12Y150_SLICE_X16Y150_A5Q;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A = CLBLM_L_X12Y150_SLICE_X17Y150_AO6;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B = CLBLM_L_X12Y150_SLICE_X17Y150_BO6;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C = CLBLM_L_X12Y150_SLICE_X17Y150_CO6;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D = CLBLM_L_X12Y150_SLICE_X17Y150_DO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A = CLBLM_L_X12Y151_SLICE_X16Y151_AO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B = CLBLM_L_X12Y151_SLICE_X16Y151_BO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C = CLBLM_L_X12Y151_SLICE_X16Y151_CO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_CMUX = CLBLM_L_X12Y151_SLICE_X16Y151_C5Q;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A = CLBLM_L_X12Y151_SLICE_X17Y151_AO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B = CLBLM_L_X12Y151_SLICE_X17Y151_BO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C = CLBLM_L_X12Y151_SLICE_X17Y151_CO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D = CLBLM_L_X12Y151_SLICE_X17Y151_DO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_AMUX = CLBLM_L_X12Y151_SLICE_X17Y151_A5Q;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_A = CLBLM_L_X12Y152_SLICE_X16Y152_AO6;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_B = CLBLM_L_X12Y152_SLICE_X16Y152_BO6;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_C = CLBLM_L_X12Y152_SLICE_X16Y152_CO6;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_D = CLBLM_L_X12Y152_SLICE_X16Y152_DO6;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_AMUX = CLBLM_L_X12Y152_SLICE_X16Y152_AO5;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_BMUX = CLBLM_L_X12Y152_SLICE_X16Y152_B5Q;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_A = CLBLM_L_X12Y152_SLICE_X17Y152_AO6;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_B = CLBLM_L_X12Y152_SLICE_X17Y152_BO6;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_C = CLBLM_L_X12Y152_SLICE_X17Y152_CO6;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_D = CLBLM_L_X12Y152_SLICE_X17Y152_DO6;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_AMUX = CLBLM_L_X12Y152_SLICE_X17Y152_A5Q;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_BMUX = CLBLM_L_X12Y152_SLICE_X17Y152_BO5;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_A = CLBLM_L_X12Y153_SLICE_X16Y153_AO6;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_B = CLBLM_L_X12Y153_SLICE_X16Y153_BO6;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_C = CLBLM_L_X12Y153_SLICE_X16Y153_CO6;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_D = CLBLM_L_X12Y153_SLICE_X16Y153_DO6;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_BMUX = CLBLM_L_X12Y153_SLICE_X16Y153_BO5;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_A = CLBLM_L_X12Y153_SLICE_X17Y153_AO6;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_B = CLBLM_L_X12Y153_SLICE_X17Y153_BO6;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_C = CLBLM_L_X12Y153_SLICE_X17Y153_CO6;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_D = CLBLM_L_X12Y153_SLICE_X17Y153_DO6;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_DMUX = CLBLM_L_X12Y153_SLICE_X17Y153_DO5;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_A = CLBLM_L_X12Y154_SLICE_X16Y154_AO6;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_B = CLBLM_L_X12Y154_SLICE_X16Y154_BO6;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_C = CLBLM_L_X12Y154_SLICE_X16Y154_CO6;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_D = CLBLM_L_X12Y154_SLICE_X16Y154_DO6;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_AMUX = CLBLM_L_X12Y154_SLICE_X16Y154_A5Q;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_CMUX = CLBLM_L_X12Y154_SLICE_X16Y154_CO5;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_DMUX = CLBLM_L_X12Y154_SLICE_X16Y154_DO5;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_A = CLBLM_L_X12Y154_SLICE_X17Y154_AO6;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_B = CLBLM_L_X12Y154_SLICE_X17Y154_BO6;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_C = CLBLM_L_X12Y154_SLICE_X17Y154_CO6;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_D = CLBLM_L_X12Y154_SLICE_X17Y154_DO6;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_AMUX = CLBLM_L_X12Y154_SLICE_X17Y154_A5Q;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_CMUX = CLBLM_L_X12Y154_SLICE_X17Y154_CO5;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_A = CLBLM_L_X12Y155_SLICE_X16Y155_AO6;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_B = CLBLM_L_X12Y155_SLICE_X16Y155_BO6;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_C = CLBLM_L_X12Y155_SLICE_X16Y155_CO6;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_D = CLBLM_L_X12Y155_SLICE_X16Y155_DO6;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_AMUX = CLBLM_L_X12Y155_SLICE_X16Y155_AO5;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_BMUX = CLBLM_L_X12Y155_SLICE_X16Y155_BO5;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_A = CLBLM_L_X12Y155_SLICE_X17Y155_AO6;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_B = CLBLM_L_X12Y155_SLICE_X17Y155_BO6;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_C = CLBLM_L_X12Y155_SLICE_X17Y155_CO6;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_D = CLBLM_L_X12Y155_SLICE_X17Y155_DO6;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_DMUX = CLBLM_L_X12Y155_SLICE_X17Y155_DO5;
  assign CLBLM_L_X12Y156_SLICE_X16Y156_A = CLBLM_L_X12Y156_SLICE_X16Y156_AO6;
  assign CLBLM_L_X12Y156_SLICE_X16Y156_B = CLBLM_L_X12Y156_SLICE_X16Y156_BO6;
  assign CLBLM_L_X12Y156_SLICE_X16Y156_C = CLBLM_L_X12Y156_SLICE_X16Y156_CO6;
  assign CLBLM_L_X12Y156_SLICE_X16Y156_D = CLBLM_L_X12Y156_SLICE_X16Y156_DO6;
  assign CLBLM_L_X12Y156_SLICE_X17Y156_A = CLBLM_L_X12Y156_SLICE_X17Y156_AO6;
  assign CLBLM_L_X12Y156_SLICE_X17Y156_B = CLBLM_L_X12Y156_SLICE_X17Y156_BO6;
  assign CLBLM_L_X12Y156_SLICE_X17Y156_C = CLBLM_L_X12Y156_SLICE_X17Y156_CO6;
  assign CLBLM_L_X12Y156_SLICE_X17Y156_D = CLBLM_L_X12Y156_SLICE_X17Y156_DO6;
  assign CLBLM_L_X12Y157_SLICE_X16Y157_A = CLBLM_L_X12Y157_SLICE_X16Y157_AO6;
  assign CLBLM_L_X12Y157_SLICE_X16Y157_B = CLBLM_L_X12Y157_SLICE_X16Y157_BO6;
  assign CLBLM_L_X12Y157_SLICE_X16Y157_C = CLBLM_L_X12Y157_SLICE_X16Y157_CO6;
  assign CLBLM_L_X12Y157_SLICE_X16Y157_D = CLBLM_L_X12Y157_SLICE_X16Y157_DO6;
  assign CLBLM_L_X12Y157_SLICE_X16Y157_AMUX = CLBLM_L_X12Y157_SLICE_X16Y157_A5Q;
  assign CLBLM_L_X12Y157_SLICE_X16Y157_DMUX = CLBLM_L_X12Y157_SLICE_X16Y157_DO5;
  assign CLBLM_L_X12Y157_SLICE_X17Y157_A = CLBLM_L_X12Y157_SLICE_X17Y157_AO6;
  assign CLBLM_L_X12Y157_SLICE_X17Y157_B = CLBLM_L_X12Y157_SLICE_X17Y157_BO6;
  assign CLBLM_L_X12Y157_SLICE_X17Y157_C = CLBLM_L_X12Y157_SLICE_X17Y157_CO6;
  assign CLBLM_L_X12Y157_SLICE_X17Y157_D = CLBLM_L_X12Y157_SLICE_X17Y157_DO6;
  assign CLBLM_L_X12Y157_SLICE_X17Y157_AMUX = CLBLM_L_X12Y157_SLICE_X17Y157_A5Q;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_A = CLBLM_L_X12Y158_SLICE_X16Y158_AO6;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_B = CLBLM_L_X12Y158_SLICE_X16Y158_BO6;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_C = CLBLM_L_X12Y158_SLICE_X16Y158_CO6;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_D = CLBLM_L_X12Y158_SLICE_X16Y158_DO6;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_AMUX = CLBLM_L_X12Y158_SLICE_X16Y158_A5Q;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_BMUX = CLBLM_L_X12Y158_SLICE_X16Y158_BO5;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_CMUX = CLBLM_L_X12Y158_SLICE_X16Y158_CO5;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_DMUX = CLBLM_L_X12Y158_SLICE_X16Y158_DO6;
  assign CLBLM_L_X12Y158_SLICE_X17Y158_A = CLBLM_L_X12Y158_SLICE_X17Y158_AO6;
  assign CLBLM_L_X12Y158_SLICE_X17Y158_B = CLBLM_L_X12Y158_SLICE_X17Y158_BO6;
  assign CLBLM_L_X12Y158_SLICE_X17Y158_C = CLBLM_L_X12Y158_SLICE_X17Y158_CO6;
  assign CLBLM_L_X12Y158_SLICE_X17Y158_D = CLBLM_L_X12Y158_SLICE_X17Y158_DO6;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_A = CLBLM_L_X12Y159_SLICE_X16Y159_AO6;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_B = CLBLM_L_X12Y159_SLICE_X16Y159_BO6;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_C = CLBLM_L_X12Y159_SLICE_X16Y159_CO6;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_D = CLBLM_L_X12Y159_SLICE_X16Y159_DO6;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_AMUX = CLBLM_L_X12Y159_SLICE_X16Y159_AO5;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_BMUX = CLBLM_L_X12Y159_SLICE_X16Y159_BO5;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_CMUX = CLBLM_L_X12Y159_SLICE_X16Y159_CO5;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_A = CLBLM_L_X12Y159_SLICE_X17Y159_AO6;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_B = CLBLM_L_X12Y159_SLICE_X17Y159_BO6;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_C = CLBLM_L_X12Y159_SLICE_X17Y159_CO6;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_D = CLBLM_L_X12Y159_SLICE_X17Y159_DO6;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_AMUX = CLBLM_L_X12Y159_SLICE_X17Y159_AO5;
  assign CLBLM_L_X16Y156_SLICE_X22Y156_A = CLBLM_L_X16Y156_SLICE_X22Y156_AO6;
  assign CLBLM_L_X16Y156_SLICE_X22Y156_B = CLBLM_L_X16Y156_SLICE_X22Y156_BO6;
  assign CLBLM_L_X16Y156_SLICE_X22Y156_C = CLBLM_L_X16Y156_SLICE_X22Y156_CO6;
  assign CLBLM_L_X16Y156_SLICE_X22Y156_D = CLBLM_L_X16Y156_SLICE_X22Y156_DO6;
  assign CLBLM_L_X16Y156_SLICE_X22Y156_AMUX = CLBLM_L_X16Y156_SLICE_X22Y156_AO5;
  assign CLBLM_L_X16Y156_SLICE_X23Y156_A = CLBLM_L_X16Y156_SLICE_X23Y156_AO6;
  assign CLBLM_L_X16Y156_SLICE_X23Y156_B = CLBLM_L_X16Y156_SLICE_X23Y156_BO6;
  assign CLBLM_L_X16Y156_SLICE_X23Y156_C = CLBLM_L_X16Y156_SLICE_X23Y156_CO6;
  assign CLBLM_L_X16Y156_SLICE_X23Y156_D = CLBLM_L_X16Y156_SLICE_X23Y156_DO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A = CLBLM_R_X3Y142_SLICE_X2Y142_AO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B = CLBLM_R_X3Y142_SLICE_X2Y142_BO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C = CLBLM_R_X3Y142_SLICE_X2Y142_CO6;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D = CLBLM_R_X3Y142_SLICE_X2Y142_DO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A = CLBLM_R_X3Y142_SLICE_X3Y142_AO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B = CLBLM_R_X3Y142_SLICE_X3Y142_BO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C = CLBLM_R_X3Y142_SLICE_X3Y142_CO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D = CLBLM_R_X3Y142_SLICE_X3Y142_DO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A = CLBLM_R_X3Y150_SLICE_X2Y150_AO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B = CLBLM_R_X3Y150_SLICE_X2Y150_BO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C = CLBLM_R_X3Y150_SLICE_X2Y150_CO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D = CLBLM_R_X3Y150_SLICE_X2Y150_DO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_AMUX = CLBLM_R_X3Y150_SLICE_X2Y150_A5Q;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_BMUX = CLBLM_R_X3Y150_SLICE_X2Y150_BO5;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A = CLBLM_R_X3Y150_SLICE_X3Y150_AO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B = CLBLM_R_X3Y150_SLICE_X3Y150_BO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C = CLBLM_R_X3Y150_SLICE_X3Y150_CO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D = CLBLM_R_X3Y150_SLICE_X3Y150_DO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A = CLBLM_R_X3Y151_SLICE_X2Y151_AO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B = CLBLM_R_X3Y151_SLICE_X2Y151_BO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C = CLBLM_R_X3Y151_SLICE_X2Y151_CO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D = CLBLM_R_X3Y151_SLICE_X2Y151_DO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_AMUX = CLBLM_R_X3Y151_SLICE_X2Y151_AO5;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_CMUX = CLBLM_R_X3Y151_SLICE_X2Y151_CO5;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A = CLBLM_R_X3Y151_SLICE_X3Y151_AO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B = CLBLM_R_X3Y151_SLICE_X3Y151_BO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C = CLBLM_R_X3Y151_SLICE_X3Y151_CO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D = CLBLM_R_X3Y151_SLICE_X3Y151_DO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_AMUX = CLBLM_R_X3Y151_SLICE_X3Y151_AO5;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_BMUX = CLBLM_R_X3Y151_SLICE_X3Y151_BO5;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A = CLBLM_R_X3Y152_SLICE_X2Y152_AO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B = CLBLM_R_X3Y152_SLICE_X2Y152_BO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_AMUX = CLBLM_R_X3Y152_SLICE_X2Y152_AO5;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_DMUX = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A = CLBLM_R_X3Y152_SLICE_X3Y152_AO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B = CLBLM_R_X3Y152_SLICE_X3Y152_BO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C = CLBLM_R_X3Y152_SLICE_X3Y152_CO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D = CLBLM_R_X3Y152_SLICE_X3Y152_DO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_AMUX = CLBLM_R_X3Y152_SLICE_X3Y152_AO5;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_BMUX = CLBLM_R_X3Y152_SLICE_X3Y152_BO5;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A = CLBLM_R_X3Y153_SLICE_X2Y153_AO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B = CLBLM_R_X3Y153_SLICE_X2Y153_BO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C = CLBLM_R_X3Y153_SLICE_X2Y153_CO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D = CLBLM_R_X3Y153_SLICE_X2Y153_DO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_AMUX = CLBLM_R_X3Y153_SLICE_X2Y153_AO5;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_BMUX = CLBLM_R_X3Y153_SLICE_X2Y153_BO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A = CLBLM_R_X3Y153_SLICE_X3Y153_AO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B = CLBLM_R_X3Y153_SLICE_X3Y153_BO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C = CLBLM_R_X3Y153_SLICE_X3Y153_CO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D = CLBLM_R_X3Y153_SLICE_X3Y153_DO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_AMUX = CLBLM_R_X3Y153_SLICE_X3Y153_AO5;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_A = CLBLM_R_X3Y154_SLICE_X2Y154_AO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_B = CLBLM_R_X3Y154_SLICE_X2Y154_BO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_C = CLBLM_R_X3Y154_SLICE_X2Y154_CO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_D = CLBLM_R_X3Y154_SLICE_X2Y154_DO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_A = CLBLM_R_X3Y154_SLICE_X3Y154_AO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_B = CLBLM_R_X3Y154_SLICE_X3Y154_BO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_C = CLBLM_R_X3Y154_SLICE_X3Y154_CO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_D = CLBLM_R_X3Y154_SLICE_X3Y154_DO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_AMUX = CLBLM_R_X3Y154_SLICE_X3Y154_AO5;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_A = CLBLM_R_X3Y155_SLICE_X2Y155_AO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_B = CLBLM_R_X3Y155_SLICE_X2Y155_BO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_C = CLBLM_R_X3Y155_SLICE_X2Y155_CO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_D = CLBLM_R_X3Y155_SLICE_X2Y155_DO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_CMUX = CLBLM_R_X3Y155_SLICE_X2Y155_CO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_A = CLBLM_R_X3Y155_SLICE_X3Y155_AO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_B = CLBLM_R_X3Y155_SLICE_X3Y155_BO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_C = CLBLM_R_X3Y155_SLICE_X3Y155_CO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_D = CLBLM_R_X3Y155_SLICE_X3Y155_DO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_CMUX = CLBLM_R_X3Y155_SLICE_X3Y155_CO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_DMUX = CLBLM_R_X3Y155_SLICE_X3Y155_DO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_A = CLBLM_R_X3Y156_SLICE_X2Y156_AO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_B = CLBLM_R_X3Y156_SLICE_X2Y156_BO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_C = CLBLM_R_X3Y156_SLICE_X2Y156_CO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_D = CLBLM_R_X3Y156_SLICE_X2Y156_DO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_BMUX = CLBLM_R_X3Y156_SLICE_X2Y156_BO6;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_A = CLBLM_R_X3Y156_SLICE_X3Y156_AO6;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_B = CLBLM_R_X3Y156_SLICE_X3Y156_BO6;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_C = CLBLM_R_X3Y156_SLICE_X3Y156_CO6;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_D = CLBLM_R_X3Y156_SLICE_X3Y156_DO6;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_AMUX = CLBLM_R_X3Y156_SLICE_X3Y156_AO5;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_CMUX = CLBLM_R_X3Y156_SLICE_X3Y156_CO6;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_A = CLBLM_R_X3Y157_SLICE_X2Y157_AO6;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_B = CLBLM_R_X3Y157_SLICE_X2Y157_BO6;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_C = CLBLM_R_X3Y157_SLICE_X2Y157_CO6;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_D = CLBLM_R_X3Y157_SLICE_X2Y157_DO6;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_AMUX = CLBLM_R_X3Y157_SLICE_X2Y157_AO5;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_A = CLBLM_R_X3Y157_SLICE_X3Y157_AO6;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_B = CLBLM_R_X3Y157_SLICE_X3Y157_BO6;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_C = CLBLM_R_X3Y157_SLICE_X3Y157_CO6;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_D = CLBLM_R_X3Y157_SLICE_X3Y157_DO6;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_DMUX = CLBLM_R_X3Y157_SLICE_X3Y157_DO6;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_A = CLBLM_R_X3Y158_SLICE_X2Y158_AO6;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_B = CLBLM_R_X3Y158_SLICE_X2Y158_BO6;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_C = CLBLM_R_X3Y158_SLICE_X2Y158_CO6;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_D = CLBLM_R_X3Y158_SLICE_X2Y158_DO6;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_AMUX = CLBLM_R_X3Y158_SLICE_X2Y158_AO5;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_A = CLBLM_R_X3Y158_SLICE_X3Y158_AO6;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_B = CLBLM_R_X3Y158_SLICE_X3Y158_BO6;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_C = CLBLM_R_X3Y158_SLICE_X3Y158_CO6;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_D = CLBLM_R_X3Y158_SLICE_X3Y158_DO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A = CLBLM_R_X5Y144_SLICE_X6Y144_AO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B = CLBLM_R_X5Y144_SLICE_X6Y144_BO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C = CLBLM_R_X5Y144_SLICE_X6Y144_CO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D = CLBLM_R_X5Y144_SLICE_X6Y144_DO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_CMUX = CLBLM_R_X5Y144_SLICE_X6Y144_CO5;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A = CLBLM_R_X5Y144_SLICE_X7Y144_AO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B = CLBLM_R_X5Y144_SLICE_X7Y144_BO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C = CLBLM_R_X5Y144_SLICE_X7Y144_CO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D = CLBLM_R_X5Y144_SLICE_X7Y144_DO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A = CLBLM_R_X5Y146_SLICE_X6Y146_AO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B = CLBLM_R_X5Y146_SLICE_X6Y146_BO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D = CLBLM_R_X5Y146_SLICE_X6Y146_DO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_AMUX = CLBLM_R_X5Y146_SLICE_X6Y146_A5Q;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_CMUX = CLBLM_R_X5Y146_SLICE_X6Y146_CO5;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A = CLBLM_R_X5Y146_SLICE_X7Y146_AO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B = CLBLM_R_X5Y146_SLICE_X7Y146_BO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C = CLBLM_R_X5Y146_SLICE_X7Y146_CO6;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D = CLBLM_R_X5Y146_SLICE_X7Y146_DO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A = CLBLM_R_X5Y147_SLICE_X6Y147_AO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B = CLBLM_R_X5Y147_SLICE_X6Y147_BO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C = CLBLM_R_X5Y147_SLICE_X6Y147_CO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D = CLBLM_R_X5Y147_SLICE_X6Y147_DO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A = CLBLM_R_X5Y147_SLICE_X7Y147_AO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B = CLBLM_R_X5Y147_SLICE_X7Y147_BO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C = CLBLM_R_X5Y147_SLICE_X7Y147_CO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D = CLBLM_R_X5Y147_SLICE_X7Y147_DO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_CMUX = CLBLM_R_X5Y147_SLICE_X7Y147_C5Q;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A = CLBLM_R_X5Y148_SLICE_X6Y148_AO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B = CLBLM_R_X5Y148_SLICE_X6Y148_BO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C = CLBLM_R_X5Y148_SLICE_X6Y148_CO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D = CLBLM_R_X5Y148_SLICE_X6Y148_DO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_AMUX = CLBLM_R_X5Y148_SLICE_X6Y148_A5Q;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_CMUX = CLBLM_R_X5Y148_SLICE_X6Y148_CO5;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A = CLBLM_R_X5Y148_SLICE_X7Y148_AO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B = CLBLM_R_X5Y148_SLICE_X7Y148_BO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C = CLBLM_R_X5Y148_SLICE_X7Y148_CO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D = CLBLM_R_X5Y148_SLICE_X7Y148_DO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_AMUX = CLBLM_R_X5Y148_SLICE_X7Y148_A5Q;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_BMUX = CLBLM_R_X5Y148_SLICE_X7Y148_B5Q;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A = CLBLM_R_X5Y149_SLICE_X6Y149_AO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B = CLBLM_R_X5Y149_SLICE_X6Y149_BO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C = CLBLM_R_X5Y149_SLICE_X6Y149_CO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D = CLBLM_R_X5Y149_SLICE_X6Y149_DO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_AMUX = CLBLM_R_X5Y149_SLICE_X6Y149_A5Q;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_BMUX = CLBLM_R_X5Y149_SLICE_X6Y149_B5Q;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_CMUX = CLBLM_R_X5Y149_SLICE_X6Y149_CO5;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A = CLBLM_R_X5Y149_SLICE_X7Y149_AO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B = CLBLM_R_X5Y149_SLICE_X7Y149_BO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C = CLBLM_R_X5Y149_SLICE_X7Y149_CO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D = CLBLM_R_X5Y149_SLICE_X7Y149_DO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_AMUX = CLBLM_R_X5Y149_SLICE_X7Y149_A5Q;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_DMUX = CLBLM_R_X5Y149_SLICE_X7Y149_DO5;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A = CLBLM_R_X5Y150_SLICE_X6Y150_AO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B = CLBLM_R_X5Y150_SLICE_X6Y150_BO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C = CLBLM_R_X5Y150_SLICE_X6Y150_CO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D = CLBLM_R_X5Y150_SLICE_X6Y150_DO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A = CLBLM_R_X5Y150_SLICE_X7Y150_AO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B = CLBLM_R_X5Y150_SLICE_X7Y150_BO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C = CLBLM_R_X5Y150_SLICE_X7Y150_CO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D = CLBLM_R_X5Y150_SLICE_X7Y150_DO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_AMUX = CLBLM_R_X5Y150_SLICE_X7Y150_A5Q;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A = CLBLM_R_X5Y151_SLICE_X6Y151_AO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B = CLBLM_R_X5Y151_SLICE_X6Y151_BO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C = CLBLM_R_X5Y151_SLICE_X6Y151_CO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D = CLBLM_R_X5Y151_SLICE_X6Y151_DO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_CMUX = CLBLM_R_X5Y151_SLICE_X6Y151_C5Q;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A = CLBLM_R_X5Y151_SLICE_X7Y151_AO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B = CLBLM_R_X5Y151_SLICE_X7Y151_BO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C = CLBLM_R_X5Y151_SLICE_X7Y151_CO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D = CLBLM_R_X5Y151_SLICE_X7Y151_DO6;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_A = CLBLM_R_X5Y152_SLICE_X6Y152_AO6;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_B = CLBLM_R_X5Y152_SLICE_X6Y152_BO6;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_C = CLBLM_R_X5Y152_SLICE_X6Y152_CO6;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_D = CLBLM_R_X5Y152_SLICE_X6Y152_DO6;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_CMUX = CLBLM_R_X5Y152_SLICE_X6Y152_CO5;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_DMUX = CLBLM_R_X5Y152_SLICE_X6Y152_DO6;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_A = CLBLM_R_X5Y152_SLICE_X7Y152_AO6;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_B = CLBLM_R_X5Y152_SLICE_X7Y152_BO6;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_C = CLBLM_R_X5Y152_SLICE_X7Y152_CO6;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_D = CLBLM_R_X5Y152_SLICE_X7Y152_DO6;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_A = CLBLM_R_X5Y153_SLICE_X6Y153_AO6;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_B = CLBLM_R_X5Y153_SLICE_X6Y153_BO6;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_C = CLBLM_R_X5Y153_SLICE_X6Y153_CO6;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_D = CLBLM_R_X5Y153_SLICE_X6Y153_DO6;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_BMUX = CLBLM_R_X5Y153_SLICE_X6Y153_BO5;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_DMUX = CLBLM_R_X5Y153_SLICE_X6Y153_DO6;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_A = CLBLM_R_X5Y153_SLICE_X7Y153_AO6;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_B = CLBLM_R_X5Y153_SLICE_X7Y153_BO6;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_C = CLBLM_R_X5Y153_SLICE_X7Y153_CO6;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_D = CLBLM_R_X5Y153_SLICE_X7Y153_DO6;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_CMUX = CLBLM_R_X5Y153_SLICE_X7Y153_CO6;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_A = CLBLM_R_X5Y154_SLICE_X6Y154_AO6;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_B = CLBLM_R_X5Y154_SLICE_X6Y154_BO6;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_C = CLBLM_R_X5Y154_SLICE_X6Y154_CO6;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_D = CLBLM_R_X5Y154_SLICE_X6Y154_DO6;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_A = CLBLM_R_X5Y154_SLICE_X7Y154_AO6;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_B = CLBLM_R_X5Y154_SLICE_X7Y154_BO6;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_C = CLBLM_R_X5Y154_SLICE_X7Y154_CO6;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_D = CLBLM_R_X5Y154_SLICE_X7Y154_DO6;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_A = CLBLM_R_X5Y155_SLICE_X6Y155_AO6;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_B = CLBLM_R_X5Y155_SLICE_X6Y155_BO6;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_C = CLBLM_R_X5Y155_SLICE_X6Y155_CO6;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_D = CLBLM_R_X5Y155_SLICE_X6Y155_DO6;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_A = CLBLM_R_X5Y155_SLICE_X7Y155_AO6;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_B = CLBLM_R_X5Y155_SLICE_X7Y155_BO6;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_C = CLBLM_R_X5Y155_SLICE_X7Y155_CO6;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_D = CLBLM_R_X5Y155_SLICE_X7Y155_DO6;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_DMUX = CLBLM_R_X5Y155_SLICE_X7Y155_DO6;
  assign CLBLM_R_X5Y156_SLICE_X6Y156_A = CLBLM_R_X5Y156_SLICE_X6Y156_AO6;
  assign CLBLM_R_X5Y156_SLICE_X6Y156_B = CLBLM_R_X5Y156_SLICE_X6Y156_BO6;
  assign CLBLM_R_X5Y156_SLICE_X6Y156_C = CLBLM_R_X5Y156_SLICE_X6Y156_CO6;
  assign CLBLM_R_X5Y156_SLICE_X6Y156_D = CLBLM_R_X5Y156_SLICE_X6Y156_DO6;
  assign CLBLM_R_X5Y156_SLICE_X7Y156_A = CLBLM_R_X5Y156_SLICE_X7Y156_AO6;
  assign CLBLM_R_X5Y156_SLICE_X7Y156_B = CLBLM_R_X5Y156_SLICE_X7Y156_BO6;
  assign CLBLM_R_X5Y156_SLICE_X7Y156_C = CLBLM_R_X5Y156_SLICE_X7Y156_CO6;
  assign CLBLM_R_X5Y156_SLICE_X7Y156_D = CLBLM_R_X5Y156_SLICE_X7Y156_DO6;
  assign CLBLM_R_X5Y157_SLICE_X6Y157_A = CLBLM_R_X5Y157_SLICE_X6Y157_AO6;
  assign CLBLM_R_X5Y157_SLICE_X6Y157_B = CLBLM_R_X5Y157_SLICE_X6Y157_BO6;
  assign CLBLM_R_X5Y157_SLICE_X6Y157_C = CLBLM_R_X5Y157_SLICE_X6Y157_CO6;
  assign CLBLM_R_X5Y157_SLICE_X6Y157_D = CLBLM_R_X5Y157_SLICE_X6Y157_DO6;
  assign CLBLM_R_X5Y157_SLICE_X6Y157_BMUX = CLBLM_R_X5Y157_SLICE_X6Y157_BO6;
  assign CLBLM_R_X5Y157_SLICE_X7Y157_A = CLBLM_R_X5Y157_SLICE_X7Y157_AO6;
  assign CLBLM_R_X5Y157_SLICE_X7Y157_B = CLBLM_R_X5Y157_SLICE_X7Y157_BO6;
  assign CLBLM_R_X5Y157_SLICE_X7Y157_C = CLBLM_R_X5Y157_SLICE_X7Y157_CO6;
  assign CLBLM_R_X5Y157_SLICE_X7Y157_D = CLBLM_R_X5Y157_SLICE_X7Y157_DO6;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_A = CLBLM_R_X5Y158_SLICE_X6Y158_AO6;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_B = CLBLM_R_X5Y158_SLICE_X6Y158_BO6;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_C = CLBLM_R_X5Y158_SLICE_X6Y158_CO6;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_D = CLBLM_R_X5Y158_SLICE_X6Y158_DO6;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_A = CLBLM_R_X5Y158_SLICE_X7Y158_AO6;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_B = CLBLM_R_X5Y158_SLICE_X7Y158_BO6;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_C = CLBLM_R_X5Y158_SLICE_X7Y158_CO6;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_D = CLBLM_R_X5Y158_SLICE_X7Y158_DO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A = CLBLM_R_X7Y144_SLICE_X8Y144_AO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B = CLBLM_R_X7Y144_SLICE_X8Y144_BO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C = CLBLM_R_X7Y144_SLICE_X8Y144_CO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D = CLBLM_R_X7Y144_SLICE_X8Y144_DO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A = CLBLM_R_X7Y144_SLICE_X9Y144_AO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B = CLBLM_R_X7Y144_SLICE_X9Y144_BO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C = CLBLM_R_X7Y144_SLICE_X9Y144_CO6;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D = CLBLM_R_X7Y144_SLICE_X9Y144_DO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A = CLBLM_R_X7Y145_SLICE_X8Y145_AO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B = CLBLM_R_X7Y145_SLICE_X8Y145_BO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C = CLBLM_R_X7Y145_SLICE_X8Y145_CO6;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D = CLBLM_R_X7Y145_SLICE_X8Y145_DO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A = CLBLM_R_X7Y145_SLICE_X9Y145_AO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B = CLBLM_R_X7Y145_SLICE_X9Y145_BO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C = CLBLM_R_X7Y145_SLICE_X9Y145_CO6;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D = CLBLM_R_X7Y145_SLICE_X9Y145_DO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A = CLBLM_R_X7Y146_SLICE_X8Y146_AO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B = CLBLM_R_X7Y146_SLICE_X8Y146_BO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D = CLBLM_R_X7Y146_SLICE_X8Y146_DO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_BMUX = CLBLM_R_X7Y146_SLICE_X8Y146_BO5;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_DMUX = CLBLM_R_X7Y146_SLICE_X8Y146_DO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A = CLBLM_R_X7Y146_SLICE_X9Y146_AO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B = CLBLM_R_X7Y146_SLICE_X9Y146_BO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C = CLBLM_R_X7Y146_SLICE_X9Y146_CO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D = CLBLM_R_X7Y146_SLICE_X9Y146_DO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_BMUX = CLBLM_R_X7Y146_SLICE_X9Y146_BO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A = CLBLM_R_X7Y147_SLICE_X8Y147_AO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B = CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C = CLBLM_R_X7Y147_SLICE_X8Y147_CO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D = CLBLM_R_X7Y147_SLICE_X8Y147_DO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_BMUX = CLBLM_R_X7Y147_SLICE_X8Y147_BO5;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_DMUX = CLBLM_R_X7Y147_SLICE_X8Y147_DO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A = CLBLM_R_X7Y147_SLICE_X9Y147_AO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B = CLBLM_R_X7Y147_SLICE_X9Y147_BO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C = CLBLM_R_X7Y147_SLICE_X9Y147_CO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D = CLBLM_R_X7Y147_SLICE_X9Y147_DO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_AMUX = CLBLM_R_X7Y147_SLICE_X9Y147_A5Q;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_DMUX = CLBLM_R_X7Y147_SLICE_X9Y147_DO5;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A = CLBLM_R_X7Y148_SLICE_X8Y148_AO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B = CLBLM_R_X7Y148_SLICE_X8Y148_BO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C = CLBLM_R_X7Y148_SLICE_X8Y148_CO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D = CLBLM_R_X7Y148_SLICE_X8Y148_DO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_AMUX = CLBLM_R_X7Y148_SLICE_X8Y148_A5Q;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_DMUX = CLBLM_R_X7Y148_SLICE_X8Y148_DO5;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A = CLBLM_R_X7Y148_SLICE_X9Y148_AO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B = CLBLM_R_X7Y148_SLICE_X9Y148_BO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C = CLBLM_R_X7Y148_SLICE_X9Y148_CO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D = CLBLM_R_X7Y148_SLICE_X9Y148_DO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_CMUX = CLBLM_R_X7Y148_SLICE_X9Y148_CO5;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A = CLBLM_R_X7Y149_SLICE_X8Y149_AO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B = CLBLM_R_X7Y149_SLICE_X8Y149_BO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C = CLBLM_R_X7Y149_SLICE_X8Y149_CO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D = CLBLM_R_X7Y149_SLICE_X8Y149_DO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_DMUX = CLBLM_R_X7Y149_SLICE_X8Y149_DO5;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A = CLBLM_R_X7Y149_SLICE_X9Y149_AO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B = CLBLM_R_X7Y149_SLICE_X9Y149_BO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C = CLBLM_R_X7Y149_SLICE_X9Y149_CO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D = CLBLM_R_X7Y149_SLICE_X9Y149_DO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_CMUX = CLBLM_R_X7Y149_SLICE_X9Y149_C5Q;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_DMUX = CLBLM_R_X7Y149_SLICE_X9Y149_DO5;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A = CLBLM_R_X7Y150_SLICE_X8Y150_AO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B = CLBLM_R_X7Y150_SLICE_X8Y150_BO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C = CLBLM_R_X7Y150_SLICE_X8Y150_CO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D = CLBLM_R_X7Y150_SLICE_X8Y150_DO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_CMUX = CLBLM_R_X7Y150_SLICE_X8Y150_CO5;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A = CLBLM_R_X7Y150_SLICE_X9Y150_AO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B = CLBLM_R_X7Y150_SLICE_X9Y150_BO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C = CLBLM_R_X7Y150_SLICE_X9Y150_CO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D = CLBLM_R_X7Y150_SLICE_X9Y150_DO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_AMUX = CLBLM_R_X7Y150_SLICE_X9Y150_AO5;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A = CLBLM_R_X7Y151_SLICE_X8Y151_AO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B = CLBLM_R_X7Y151_SLICE_X8Y151_BO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C = CLBLM_R_X7Y151_SLICE_X8Y151_CO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D = CLBLM_R_X7Y151_SLICE_X8Y151_DO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A = CLBLM_R_X7Y151_SLICE_X9Y151_AO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B = CLBLM_R_X7Y151_SLICE_X9Y151_BO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C = CLBLM_R_X7Y151_SLICE_X9Y151_CO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D = CLBLM_R_X7Y151_SLICE_X9Y151_DO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_CMUX = CLBLM_R_X7Y151_SLICE_X9Y151_C5Q;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_DMUX = CLBLM_R_X7Y151_SLICE_X9Y151_DO6;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_A = CLBLM_R_X7Y152_SLICE_X8Y152_AO6;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_B = CLBLM_R_X7Y152_SLICE_X8Y152_BO6;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_C = CLBLM_R_X7Y152_SLICE_X8Y152_CO6;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_D = CLBLM_R_X7Y152_SLICE_X8Y152_DO6;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_AMUX = CLBLM_R_X7Y152_SLICE_X8Y152_A5Q;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_BMUX = CLBLM_R_X7Y152_SLICE_X8Y152_BO5;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_A = CLBLM_R_X7Y152_SLICE_X9Y152_AO6;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_B = CLBLM_R_X7Y152_SLICE_X9Y152_BO6;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_C = CLBLM_R_X7Y152_SLICE_X9Y152_CO6;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_D = CLBLM_R_X7Y152_SLICE_X9Y152_DO6;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_CMUX = CLBLM_R_X7Y152_SLICE_X9Y152_CO5;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_A = CLBLM_R_X7Y153_SLICE_X8Y153_AO6;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_B = CLBLM_R_X7Y153_SLICE_X8Y153_BO6;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_C = CLBLM_R_X7Y153_SLICE_X8Y153_CO6;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_D = CLBLM_R_X7Y153_SLICE_X8Y153_DO6;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_AMUX = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_A = CLBLM_R_X7Y153_SLICE_X9Y153_AO6;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_B = CLBLM_R_X7Y153_SLICE_X9Y153_BO6;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_C = CLBLM_R_X7Y153_SLICE_X9Y153_CO6;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_D = CLBLM_R_X7Y153_SLICE_X9Y153_DO6;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_CMUX = CLBLM_R_X7Y153_SLICE_X9Y153_CO5;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_A = CLBLM_R_X7Y154_SLICE_X8Y154_AO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_B = CLBLM_R_X7Y154_SLICE_X8Y154_BO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_C = CLBLM_R_X7Y154_SLICE_X8Y154_CO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_D = CLBLM_R_X7Y154_SLICE_X8Y154_DO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_AMUX = CLBLM_R_X7Y154_SLICE_X8Y154_AO5;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_A = CLBLM_R_X7Y154_SLICE_X9Y154_AO6;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_B = CLBLM_R_X7Y154_SLICE_X9Y154_BO6;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_C = CLBLM_R_X7Y154_SLICE_X9Y154_CO6;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_D = CLBLM_R_X7Y154_SLICE_X9Y154_DO6;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_A = CLBLM_R_X7Y155_SLICE_X8Y155_AO6;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_B = CLBLM_R_X7Y155_SLICE_X8Y155_BO6;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_C = CLBLM_R_X7Y155_SLICE_X8Y155_CO6;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_D = CLBLM_R_X7Y155_SLICE_X8Y155_DO6;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_AMUX = CLBLM_R_X7Y155_SLICE_X8Y155_A5Q;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_BMUX = CLBLM_R_X7Y155_SLICE_X8Y155_BO5;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_A = CLBLM_R_X7Y155_SLICE_X9Y155_AO6;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_B = CLBLM_R_X7Y155_SLICE_X9Y155_BO6;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_C = CLBLM_R_X7Y155_SLICE_X9Y155_CO6;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_D = CLBLM_R_X7Y155_SLICE_X9Y155_DO6;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_AMUX = CLBLM_R_X7Y155_SLICE_X9Y155_A5Q;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_CMUX = CLBLM_R_X7Y155_SLICE_X9Y155_CO5;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_DMUX = CLBLM_R_X7Y155_SLICE_X9Y155_DO6;
  assign CLBLM_R_X7Y156_SLICE_X8Y156_A = CLBLM_R_X7Y156_SLICE_X8Y156_AO6;
  assign CLBLM_R_X7Y156_SLICE_X8Y156_B = CLBLM_R_X7Y156_SLICE_X8Y156_BO6;
  assign CLBLM_R_X7Y156_SLICE_X8Y156_C = CLBLM_R_X7Y156_SLICE_X8Y156_CO6;
  assign CLBLM_R_X7Y156_SLICE_X8Y156_D = CLBLM_R_X7Y156_SLICE_X8Y156_DO6;
  assign CLBLM_R_X7Y156_SLICE_X9Y156_A = CLBLM_R_X7Y156_SLICE_X9Y156_AO6;
  assign CLBLM_R_X7Y156_SLICE_X9Y156_B = CLBLM_R_X7Y156_SLICE_X9Y156_BO6;
  assign CLBLM_R_X7Y156_SLICE_X9Y156_C = CLBLM_R_X7Y156_SLICE_X9Y156_CO6;
  assign CLBLM_R_X7Y156_SLICE_X9Y156_D = CLBLM_R_X7Y156_SLICE_X9Y156_DO6;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_A = CLBLM_R_X7Y157_SLICE_X8Y157_AO6;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_B = CLBLM_R_X7Y157_SLICE_X8Y157_BO6;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_C = CLBLM_R_X7Y157_SLICE_X8Y157_CO6;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_D = CLBLM_R_X7Y157_SLICE_X8Y157_DO6;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_A = CLBLM_R_X7Y157_SLICE_X9Y157_AO6;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_B = CLBLM_R_X7Y157_SLICE_X9Y157_BO6;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_C = CLBLM_R_X7Y157_SLICE_X9Y157_CO6;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_D = CLBLM_R_X7Y157_SLICE_X9Y157_DO6;
  assign CLBLM_R_X7Y158_SLICE_X8Y158_A = CLBLM_R_X7Y158_SLICE_X8Y158_AO6;
  assign CLBLM_R_X7Y158_SLICE_X8Y158_B = CLBLM_R_X7Y158_SLICE_X8Y158_BO6;
  assign CLBLM_R_X7Y158_SLICE_X8Y158_C = CLBLM_R_X7Y158_SLICE_X8Y158_CO6;
  assign CLBLM_R_X7Y158_SLICE_X8Y158_D = CLBLM_R_X7Y158_SLICE_X8Y158_DO6;
  assign CLBLM_R_X7Y158_SLICE_X8Y158_CMUX = CLBLM_R_X7Y158_SLICE_X8Y158_CO5;
  assign CLBLM_R_X7Y158_SLICE_X9Y158_A = CLBLM_R_X7Y158_SLICE_X9Y158_AO6;
  assign CLBLM_R_X7Y158_SLICE_X9Y158_B = CLBLM_R_X7Y158_SLICE_X9Y158_BO6;
  assign CLBLM_R_X7Y158_SLICE_X9Y158_C = CLBLM_R_X7Y158_SLICE_X9Y158_CO6;
  assign CLBLM_R_X7Y158_SLICE_X9Y158_D = CLBLM_R_X7Y158_SLICE_X9Y158_DO6;
  assign CLBLM_R_X7Y159_SLICE_X8Y159_A = CLBLM_R_X7Y159_SLICE_X8Y159_AO6;
  assign CLBLM_R_X7Y159_SLICE_X8Y159_B = CLBLM_R_X7Y159_SLICE_X8Y159_BO6;
  assign CLBLM_R_X7Y159_SLICE_X8Y159_C = CLBLM_R_X7Y159_SLICE_X8Y159_CO6;
  assign CLBLM_R_X7Y159_SLICE_X8Y159_D = CLBLM_R_X7Y159_SLICE_X8Y159_DO6;
  assign CLBLM_R_X7Y159_SLICE_X8Y159_BMUX = CLBLM_R_X7Y159_SLICE_X8Y159_BO5;
  assign CLBLM_R_X7Y159_SLICE_X9Y159_A = CLBLM_R_X7Y159_SLICE_X9Y159_AO6;
  assign CLBLM_R_X7Y159_SLICE_X9Y159_B = CLBLM_R_X7Y159_SLICE_X9Y159_BO6;
  assign CLBLM_R_X7Y159_SLICE_X9Y159_C = CLBLM_R_X7Y159_SLICE_X9Y159_CO6;
  assign CLBLM_R_X7Y159_SLICE_X9Y159_D = CLBLM_R_X7Y159_SLICE_X9Y159_DO6;
  assign CLBLM_R_X7Y159_SLICE_X9Y159_BMUX = CLBLM_R_X7Y159_SLICE_X9Y159_BO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A = CLBLM_R_X11Y144_SLICE_X14Y144_AO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B = CLBLM_R_X11Y144_SLICE_X14Y144_BO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C = CLBLM_R_X11Y144_SLICE_X14Y144_CO6;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D = CLBLM_R_X11Y144_SLICE_X14Y144_DO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A = CLBLM_R_X11Y144_SLICE_X15Y144_AO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B = CLBLM_R_X11Y144_SLICE_X15Y144_BO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C = CLBLM_R_X11Y144_SLICE_X15Y144_CO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D = CLBLM_R_X11Y144_SLICE_X15Y144_DO6;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_AMUX = CLBLM_R_X11Y144_SLICE_X15Y144_A5Q;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A = CLBLM_R_X11Y146_SLICE_X14Y146_AO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B = CLBLM_R_X11Y146_SLICE_X14Y146_BO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C = CLBLM_R_X11Y146_SLICE_X14Y146_CO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D = CLBLM_R_X11Y146_SLICE_X14Y146_DO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A = CLBLM_R_X11Y146_SLICE_X15Y146_AO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B = CLBLM_R_X11Y146_SLICE_X15Y146_BO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C = CLBLM_R_X11Y146_SLICE_X15Y146_CO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D = CLBLM_R_X11Y146_SLICE_X15Y146_DO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_DMUX = CLBLM_R_X11Y146_SLICE_X15Y146_DO5;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A = CLBLM_R_X11Y147_SLICE_X14Y147_AO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B = CLBLM_R_X11Y147_SLICE_X14Y147_BO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D = CLBLM_R_X11Y147_SLICE_X14Y147_DO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_AMUX = CLBLM_R_X11Y147_SLICE_X14Y147_AO5;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A = CLBLM_R_X11Y147_SLICE_X15Y147_AO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B = CLBLM_R_X11Y147_SLICE_X15Y147_BO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C = CLBLM_R_X11Y147_SLICE_X15Y147_CO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D = CLBLM_R_X11Y147_SLICE_X15Y147_DO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_BMUX = CLBLM_R_X11Y147_SLICE_X15Y147_BO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A = CLBLM_R_X11Y148_SLICE_X14Y148_AO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B = CLBLM_R_X11Y148_SLICE_X14Y148_BO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C = CLBLM_R_X11Y148_SLICE_X14Y148_CO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D = CLBLM_R_X11Y148_SLICE_X14Y148_DO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A = CLBLM_R_X11Y148_SLICE_X15Y148_AO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B = CLBLM_R_X11Y148_SLICE_X15Y148_BO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C = CLBLM_R_X11Y148_SLICE_X15Y148_CO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D = CLBLM_R_X11Y148_SLICE_X15Y148_DO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A = CLBLM_R_X11Y149_SLICE_X14Y149_AO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B = CLBLM_R_X11Y149_SLICE_X14Y149_BO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C = CLBLM_R_X11Y149_SLICE_X14Y149_CO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D = CLBLM_R_X11Y149_SLICE_X14Y149_DO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A = CLBLM_R_X11Y149_SLICE_X15Y149_AO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B = CLBLM_R_X11Y149_SLICE_X15Y149_BO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C = CLBLM_R_X11Y149_SLICE_X15Y149_CO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D = CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_AMUX = CLBLM_R_X11Y149_SLICE_X15Y149_A5Q;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_DMUX = CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A = CLBLM_R_X11Y150_SLICE_X14Y150_AO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B = CLBLM_R_X11Y150_SLICE_X14Y150_BO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C = CLBLM_R_X11Y150_SLICE_X14Y150_CO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D = CLBLM_R_X11Y150_SLICE_X14Y150_DO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_BMUX = CLBLM_R_X11Y150_SLICE_X14Y150_BO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A = CLBLM_R_X11Y150_SLICE_X15Y150_AO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B = CLBLM_R_X11Y150_SLICE_X15Y150_BO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C = CLBLM_R_X11Y150_SLICE_X15Y150_CO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D = CLBLM_R_X11Y150_SLICE_X15Y150_DO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_AMUX = CLBLM_R_X11Y150_SLICE_X15Y150_AO5;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A = CLBLM_R_X11Y151_SLICE_X14Y151_AO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B = CLBLM_R_X11Y151_SLICE_X14Y151_BO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C = CLBLM_R_X11Y151_SLICE_X14Y151_CO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D = CLBLM_R_X11Y151_SLICE_X14Y151_DO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A = CLBLM_R_X11Y151_SLICE_X15Y151_AO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B = CLBLM_R_X11Y151_SLICE_X15Y151_BO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C = CLBLM_R_X11Y151_SLICE_X15Y151_CO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D = CLBLM_R_X11Y151_SLICE_X15Y151_DO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_AMUX = CLBLM_R_X11Y151_SLICE_X15Y151_A5Q;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_DMUX = CLBLM_R_X11Y151_SLICE_X15Y151_DO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A = CLBLM_R_X11Y152_SLICE_X14Y152_AO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B = CLBLM_R_X11Y152_SLICE_X14Y152_BO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C = CLBLM_R_X11Y152_SLICE_X14Y152_CO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D = CLBLM_R_X11Y152_SLICE_X14Y152_DO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_BMUX = CLBLM_R_X11Y152_SLICE_X14Y152_B5Q;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_DMUX = CLBLM_R_X11Y152_SLICE_X14Y152_DO5;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A = CLBLM_R_X11Y152_SLICE_X15Y152_AO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B = CLBLM_R_X11Y152_SLICE_X15Y152_BO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C = CLBLM_R_X11Y152_SLICE_X15Y152_CO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D = CLBLM_R_X11Y152_SLICE_X15Y152_DO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A = CLBLM_R_X11Y153_SLICE_X14Y153_AO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B = CLBLM_R_X11Y153_SLICE_X14Y153_BO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C = CLBLM_R_X11Y153_SLICE_X14Y153_CO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D = CLBLM_R_X11Y153_SLICE_X14Y153_DO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A = CLBLM_R_X11Y153_SLICE_X15Y153_AO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B = CLBLM_R_X11Y153_SLICE_X15Y153_BO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C = CLBLM_R_X11Y153_SLICE_X15Y153_CO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D = CLBLM_R_X11Y153_SLICE_X15Y153_DO6;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_A = CLBLM_R_X11Y154_SLICE_X14Y154_AO6;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_B = CLBLM_R_X11Y154_SLICE_X14Y154_BO6;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_C = CLBLM_R_X11Y154_SLICE_X14Y154_CO6;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_D = CLBLM_R_X11Y154_SLICE_X14Y154_DO6;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_BMUX = CLBLM_R_X11Y154_SLICE_X14Y154_BO5;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_DMUX = CLBLM_R_X11Y154_SLICE_X14Y154_D5Q;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_A = CLBLM_R_X11Y154_SLICE_X15Y154_AO6;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_B = CLBLM_R_X11Y154_SLICE_X15Y154_BO6;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_C = CLBLM_R_X11Y154_SLICE_X15Y154_CO6;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_D = CLBLM_R_X11Y154_SLICE_X15Y154_DO6;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_CMUX = CLBLM_R_X11Y154_SLICE_X15Y154_CO5;
  assign CLBLM_R_X11Y155_SLICE_X14Y155_A = CLBLM_R_X11Y155_SLICE_X14Y155_AO6;
  assign CLBLM_R_X11Y155_SLICE_X14Y155_B = CLBLM_R_X11Y155_SLICE_X14Y155_BO6;
  assign CLBLM_R_X11Y155_SLICE_X14Y155_C = CLBLM_R_X11Y155_SLICE_X14Y155_CO6;
  assign CLBLM_R_X11Y155_SLICE_X14Y155_D = CLBLM_R_X11Y155_SLICE_X14Y155_DO6;
  assign CLBLM_R_X11Y155_SLICE_X15Y155_A = CLBLM_R_X11Y155_SLICE_X15Y155_AO6;
  assign CLBLM_R_X11Y155_SLICE_X15Y155_B = CLBLM_R_X11Y155_SLICE_X15Y155_BO6;
  assign CLBLM_R_X11Y155_SLICE_X15Y155_C = CLBLM_R_X11Y155_SLICE_X15Y155_CO6;
  assign CLBLM_R_X11Y155_SLICE_X15Y155_D = CLBLM_R_X11Y155_SLICE_X15Y155_DO6;
  assign CLBLM_R_X11Y155_SLICE_X15Y155_DMUX = CLBLM_R_X11Y155_SLICE_X15Y155_DO6;
  assign CLBLM_R_X11Y156_SLICE_X14Y156_A = CLBLM_R_X11Y156_SLICE_X14Y156_AO6;
  assign CLBLM_R_X11Y156_SLICE_X14Y156_B = CLBLM_R_X11Y156_SLICE_X14Y156_BO6;
  assign CLBLM_R_X11Y156_SLICE_X14Y156_C = CLBLM_R_X11Y156_SLICE_X14Y156_CO6;
  assign CLBLM_R_X11Y156_SLICE_X14Y156_D = CLBLM_R_X11Y156_SLICE_X14Y156_DO6;
  assign CLBLM_R_X11Y156_SLICE_X15Y156_A = CLBLM_R_X11Y156_SLICE_X15Y156_AO6;
  assign CLBLM_R_X11Y156_SLICE_X15Y156_B = CLBLM_R_X11Y156_SLICE_X15Y156_BO6;
  assign CLBLM_R_X11Y156_SLICE_X15Y156_C = CLBLM_R_X11Y156_SLICE_X15Y156_CO6;
  assign CLBLM_R_X11Y156_SLICE_X15Y156_D = CLBLM_R_X11Y156_SLICE_X15Y156_DO6;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_A = CLBLM_R_X11Y157_SLICE_X14Y157_AO6;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_B = CLBLM_R_X11Y157_SLICE_X14Y157_BO6;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_C = CLBLM_R_X11Y157_SLICE_X14Y157_CO6;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_D = CLBLM_R_X11Y157_SLICE_X14Y157_DO6;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_A = CLBLM_R_X11Y157_SLICE_X15Y157_AO6;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_B = CLBLM_R_X11Y157_SLICE_X15Y157_BO6;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_C = CLBLM_R_X11Y157_SLICE_X15Y157_CO6;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_D = CLBLM_R_X11Y157_SLICE_X15Y157_DO6;
  assign CLBLM_R_X11Y158_SLICE_X14Y158_A = CLBLM_R_X11Y158_SLICE_X14Y158_AO6;
  assign CLBLM_R_X11Y158_SLICE_X14Y158_B = CLBLM_R_X11Y158_SLICE_X14Y158_BO6;
  assign CLBLM_R_X11Y158_SLICE_X14Y158_C = CLBLM_R_X11Y158_SLICE_X14Y158_CO6;
  assign CLBLM_R_X11Y158_SLICE_X14Y158_D = CLBLM_R_X11Y158_SLICE_X14Y158_DO6;
  assign CLBLM_R_X11Y158_SLICE_X14Y158_DMUX = CLBLM_R_X11Y158_SLICE_X14Y158_DO5;
  assign CLBLM_R_X11Y158_SLICE_X15Y158_A = CLBLM_R_X11Y158_SLICE_X15Y158_AO6;
  assign CLBLM_R_X11Y158_SLICE_X15Y158_B = CLBLM_R_X11Y158_SLICE_X15Y158_BO6;
  assign CLBLM_R_X11Y158_SLICE_X15Y158_C = CLBLM_R_X11Y158_SLICE_X15Y158_CO6;
  assign CLBLM_R_X11Y158_SLICE_X15Y158_D = CLBLM_R_X11Y158_SLICE_X15Y158_DO6;
  assign CLBLM_R_X11Y158_SLICE_X15Y158_BMUX = CLBLM_R_X11Y158_SLICE_X15Y158_BO5;
  assign CLBLM_R_X11Y159_SLICE_X14Y159_A = CLBLM_R_X11Y159_SLICE_X14Y159_AO6;
  assign CLBLM_R_X11Y159_SLICE_X14Y159_B = CLBLM_R_X11Y159_SLICE_X14Y159_BO6;
  assign CLBLM_R_X11Y159_SLICE_X14Y159_C = CLBLM_R_X11Y159_SLICE_X14Y159_CO6;
  assign CLBLM_R_X11Y159_SLICE_X14Y159_D = CLBLM_R_X11Y159_SLICE_X14Y159_DO6;
  assign CLBLM_R_X11Y159_SLICE_X15Y159_A = CLBLM_R_X11Y159_SLICE_X15Y159_AO6;
  assign CLBLM_R_X11Y159_SLICE_X15Y159_B = CLBLM_R_X11Y159_SLICE_X15Y159_BO6;
  assign CLBLM_R_X11Y159_SLICE_X15Y159_C = CLBLM_R_X11Y159_SLICE_X15Y159_CO6;
  assign CLBLM_R_X11Y159_SLICE_X15Y159_D = CLBLM_R_X11Y159_SLICE_X15Y159_DO6;
  assign CLBLM_R_X11Y159_SLICE_X15Y159_CMUX = CLBLM_R_X11Y159_SLICE_X15Y159_CO5;
  assign CLBLM_R_X11Y159_SLICE_X15Y159_DMUX = CLBLM_R_X11Y159_SLICE_X15Y159_DO5;
  assign CLBLM_R_X11Y160_SLICE_X14Y160_A = CLBLM_R_X11Y160_SLICE_X14Y160_AO6;
  assign CLBLM_R_X11Y160_SLICE_X14Y160_B = CLBLM_R_X11Y160_SLICE_X14Y160_BO6;
  assign CLBLM_R_X11Y160_SLICE_X14Y160_C = CLBLM_R_X11Y160_SLICE_X14Y160_CO6;
  assign CLBLM_R_X11Y160_SLICE_X14Y160_D = CLBLM_R_X11Y160_SLICE_X14Y160_DO6;
  assign CLBLM_R_X11Y160_SLICE_X15Y160_A = CLBLM_R_X11Y160_SLICE_X15Y160_AO6;
  assign CLBLM_R_X11Y160_SLICE_X15Y160_B = CLBLM_R_X11Y160_SLICE_X15Y160_BO6;
  assign CLBLM_R_X11Y160_SLICE_X15Y160_C = CLBLM_R_X11Y160_SLICE_X15Y160_CO6;
  assign CLBLM_R_X11Y160_SLICE_X15Y160_D = CLBLM_R_X11Y160_SLICE_X15Y160_DO6;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_A = CLBLM_R_X13Y147_SLICE_X18Y147_AO6;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_B = CLBLM_R_X13Y147_SLICE_X18Y147_BO6;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_C = CLBLM_R_X13Y147_SLICE_X18Y147_CO6;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_D = CLBLM_R_X13Y147_SLICE_X18Y147_DO6;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_AMUX = CLBLM_R_X13Y147_SLICE_X18Y147_AO5;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_BMUX = CLBLM_R_X13Y147_SLICE_X18Y147_BO5;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_A = CLBLM_R_X13Y147_SLICE_X19Y147_AO6;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_B = CLBLM_R_X13Y147_SLICE_X19Y147_BO6;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_C = CLBLM_R_X13Y147_SLICE_X19Y147_CO6;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_D = CLBLM_R_X13Y147_SLICE_X19Y147_DO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_A = CLBLM_R_X13Y148_SLICE_X18Y148_AO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_B = CLBLM_R_X13Y148_SLICE_X18Y148_BO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_C = CLBLM_R_X13Y148_SLICE_X18Y148_CO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_D = CLBLM_R_X13Y148_SLICE_X18Y148_DO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_AMUX = CLBLM_R_X13Y148_SLICE_X18Y148_AO5;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_BMUX = CLBLM_R_X13Y148_SLICE_X18Y148_BO5;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_CMUX = CLBLM_R_X13Y148_SLICE_X18Y148_CO6;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_A = CLBLM_R_X13Y148_SLICE_X19Y148_AO6;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_B = CLBLM_R_X13Y148_SLICE_X19Y148_BO6;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_C = CLBLM_R_X13Y148_SLICE_X19Y148_CO6;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_D = CLBLM_R_X13Y148_SLICE_X19Y148_DO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_A = CLBLM_R_X13Y149_SLICE_X18Y149_AO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_B = CLBLM_R_X13Y149_SLICE_X18Y149_BO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_C = CLBLM_R_X13Y149_SLICE_X18Y149_CO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_D = CLBLM_R_X13Y149_SLICE_X18Y149_DO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_AMUX = CLBLM_R_X13Y149_SLICE_X18Y149_A5Q;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_A = CLBLM_R_X13Y149_SLICE_X19Y149_AO6;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_B = CLBLM_R_X13Y149_SLICE_X19Y149_BO6;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_C = CLBLM_R_X13Y149_SLICE_X19Y149_CO6;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_D = CLBLM_R_X13Y149_SLICE_X19Y149_DO6;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_AMUX = CLBLM_R_X13Y149_SLICE_X19Y149_A5Q;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_BMUX = CLBLM_R_X13Y149_SLICE_X19Y149_BO5;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_A = CLBLM_R_X13Y150_SLICE_X18Y150_AO6;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_B = CLBLM_R_X13Y150_SLICE_X18Y150_BO6;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_C = CLBLM_R_X13Y150_SLICE_X18Y150_CO6;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_D = CLBLM_R_X13Y150_SLICE_X18Y150_DO6;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_DMUX = CLBLM_R_X13Y150_SLICE_X18Y150_DO5;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_A = CLBLM_R_X13Y150_SLICE_X19Y150_AO6;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_B = CLBLM_R_X13Y150_SLICE_X19Y150_BO6;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_C = CLBLM_R_X13Y150_SLICE_X19Y150_CO6;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_D = CLBLM_R_X13Y150_SLICE_X19Y150_DO6;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_A = CLBLM_R_X13Y151_SLICE_X18Y151_AO6;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_B = CLBLM_R_X13Y151_SLICE_X18Y151_BO6;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_C = CLBLM_R_X13Y151_SLICE_X18Y151_CO6;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_D = CLBLM_R_X13Y151_SLICE_X18Y151_DO6;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_A = CLBLM_R_X13Y151_SLICE_X19Y151_AO6;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_B = CLBLM_R_X13Y151_SLICE_X19Y151_BO6;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_C = CLBLM_R_X13Y151_SLICE_X19Y151_CO6;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_D = CLBLM_R_X13Y151_SLICE_X19Y151_DO6;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_A = CLBLM_R_X13Y152_SLICE_X18Y152_AO6;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_B = CLBLM_R_X13Y152_SLICE_X18Y152_BO6;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_C = CLBLM_R_X13Y152_SLICE_X18Y152_CO6;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_D = CLBLM_R_X13Y152_SLICE_X18Y152_DO6;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_AMUX = CLBLM_R_X13Y152_SLICE_X18Y152_A5Q;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_BMUX = CLBLM_R_X13Y152_SLICE_X18Y152_BO5;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_A = CLBLM_R_X13Y152_SLICE_X19Y152_AO6;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_B = CLBLM_R_X13Y152_SLICE_X19Y152_BO6;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_C = CLBLM_R_X13Y152_SLICE_X19Y152_CO6;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_D = CLBLM_R_X13Y152_SLICE_X19Y152_DO6;
  assign CLBLM_R_X13Y153_SLICE_X18Y153_A = CLBLM_R_X13Y153_SLICE_X18Y153_AO6;
  assign CLBLM_R_X13Y153_SLICE_X18Y153_B = CLBLM_R_X13Y153_SLICE_X18Y153_BO6;
  assign CLBLM_R_X13Y153_SLICE_X18Y153_C = CLBLM_R_X13Y153_SLICE_X18Y153_CO6;
  assign CLBLM_R_X13Y153_SLICE_X18Y153_D = CLBLM_R_X13Y153_SLICE_X18Y153_DO6;
  assign CLBLM_R_X13Y153_SLICE_X18Y153_CMUX = CLBLM_R_X13Y153_SLICE_X18Y153_C5Q;
  assign CLBLM_R_X13Y153_SLICE_X19Y153_A = CLBLM_R_X13Y153_SLICE_X19Y153_AO6;
  assign CLBLM_R_X13Y153_SLICE_X19Y153_B = CLBLM_R_X13Y153_SLICE_X19Y153_BO6;
  assign CLBLM_R_X13Y153_SLICE_X19Y153_C = CLBLM_R_X13Y153_SLICE_X19Y153_CO6;
  assign CLBLM_R_X13Y153_SLICE_X19Y153_D = CLBLM_R_X13Y153_SLICE_X19Y153_DO6;
  assign CLBLM_R_X13Y154_SLICE_X18Y154_A = CLBLM_R_X13Y154_SLICE_X18Y154_AO6;
  assign CLBLM_R_X13Y154_SLICE_X18Y154_B = CLBLM_R_X13Y154_SLICE_X18Y154_BO6;
  assign CLBLM_R_X13Y154_SLICE_X18Y154_C = CLBLM_R_X13Y154_SLICE_X18Y154_CO6;
  assign CLBLM_R_X13Y154_SLICE_X18Y154_D = CLBLM_R_X13Y154_SLICE_X18Y154_DO6;
  assign CLBLM_R_X13Y154_SLICE_X19Y154_A = CLBLM_R_X13Y154_SLICE_X19Y154_AO6;
  assign CLBLM_R_X13Y154_SLICE_X19Y154_B = CLBLM_R_X13Y154_SLICE_X19Y154_BO6;
  assign CLBLM_R_X13Y154_SLICE_X19Y154_C = CLBLM_R_X13Y154_SLICE_X19Y154_CO6;
  assign CLBLM_R_X13Y154_SLICE_X19Y154_D = CLBLM_R_X13Y154_SLICE_X19Y154_DO6;
  assign CLBLM_R_X13Y155_SLICE_X18Y155_A = CLBLM_R_X13Y155_SLICE_X18Y155_AO6;
  assign CLBLM_R_X13Y155_SLICE_X18Y155_B = CLBLM_R_X13Y155_SLICE_X18Y155_BO6;
  assign CLBLM_R_X13Y155_SLICE_X18Y155_C = CLBLM_R_X13Y155_SLICE_X18Y155_CO6;
  assign CLBLM_R_X13Y155_SLICE_X18Y155_D = CLBLM_R_X13Y155_SLICE_X18Y155_DO6;
  assign CLBLM_R_X13Y155_SLICE_X18Y155_CMUX = CLBLM_R_X13Y155_SLICE_X18Y155_CO5;
  assign CLBLM_R_X13Y155_SLICE_X18Y155_DMUX = CLBLM_R_X13Y155_SLICE_X18Y155_DO6;
  assign CLBLM_R_X13Y155_SLICE_X19Y155_A = CLBLM_R_X13Y155_SLICE_X19Y155_AO6;
  assign CLBLM_R_X13Y155_SLICE_X19Y155_B = CLBLM_R_X13Y155_SLICE_X19Y155_BO6;
  assign CLBLM_R_X13Y155_SLICE_X19Y155_C = CLBLM_R_X13Y155_SLICE_X19Y155_CO6;
  assign CLBLM_R_X13Y155_SLICE_X19Y155_D = CLBLM_R_X13Y155_SLICE_X19Y155_DO6;
  assign CLBLM_R_X13Y156_SLICE_X18Y156_A = CLBLM_R_X13Y156_SLICE_X18Y156_AO6;
  assign CLBLM_R_X13Y156_SLICE_X18Y156_B = CLBLM_R_X13Y156_SLICE_X18Y156_BO6;
  assign CLBLM_R_X13Y156_SLICE_X18Y156_C = CLBLM_R_X13Y156_SLICE_X18Y156_CO6;
  assign CLBLM_R_X13Y156_SLICE_X18Y156_D = CLBLM_R_X13Y156_SLICE_X18Y156_DO6;
  assign CLBLM_R_X13Y156_SLICE_X19Y156_A = CLBLM_R_X13Y156_SLICE_X19Y156_AO6;
  assign CLBLM_R_X13Y156_SLICE_X19Y156_B = CLBLM_R_X13Y156_SLICE_X19Y156_BO6;
  assign CLBLM_R_X13Y156_SLICE_X19Y156_C = CLBLM_R_X13Y156_SLICE_X19Y156_CO6;
  assign CLBLM_R_X13Y156_SLICE_X19Y156_D = CLBLM_R_X13Y156_SLICE_X19Y156_DO6;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_A = CLBLM_R_X13Y157_SLICE_X18Y157_AO6;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_B = CLBLM_R_X13Y157_SLICE_X18Y157_BO6;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_C = CLBLM_R_X13Y157_SLICE_X18Y157_CO6;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_D = CLBLM_R_X13Y157_SLICE_X18Y157_DO6;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_AMUX = CLBLM_R_X13Y157_SLICE_X18Y157_AO5;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_BMUX = CLBLM_R_X13Y157_SLICE_X18Y157_BO6;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_CMUX = CLBLM_R_X13Y157_SLICE_X18Y157_CO6;
  assign CLBLM_R_X13Y157_SLICE_X19Y157_A = CLBLM_R_X13Y157_SLICE_X19Y157_AO6;
  assign CLBLM_R_X13Y157_SLICE_X19Y157_B = CLBLM_R_X13Y157_SLICE_X19Y157_BO6;
  assign CLBLM_R_X13Y157_SLICE_X19Y157_C = CLBLM_R_X13Y157_SLICE_X19Y157_CO6;
  assign CLBLM_R_X13Y157_SLICE_X19Y157_D = CLBLM_R_X13Y157_SLICE_X19Y157_DO6;
  assign CLBLM_R_X13Y157_SLICE_X19Y157_BMUX = CLBLM_R_X13Y157_SLICE_X19Y157_BO6;
  assign CLBLM_R_X13Y158_SLICE_X18Y158_A = CLBLM_R_X13Y158_SLICE_X18Y158_AO6;
  assign CLBLM_R_X13Y158_SLICE_X18Y158_B = CLBLM_R_X13Y158_SLICE_X18Y158_BO6;
  assign CLBLM_R_X13Y158_SLICE_X18Y158_C = CLBLM_R_X13Y158_SLICE_X18Y158_CO6;
  assign CLBLM_R_X13Y158_SLICE_X18Y158_D = CLBLM_R_X13Y158_SLICE_X18Y158_DO6;
  assign CLBLM_R_X13Y158_SLICE_X19Y158_A = CLBLM_R_X13Y158_SLICE_X19Y158_AO6;
  assign CLBLM_R_X13Y158_SLICE_X19Y158_B = CLBLM_R_X13Y158_SLICE_X19Y158_BO6;
  assign CLBLM_R_X13Y158_SLICE_X19Y158_C = CLBLM_R_X13Y158_SLICE_X19Y158_CO6;
  assign CLBLM_R_X13Y158_SLICE_X19Y158_D = CLBLM_R_X13Y158_SLICE_X19Y158_DO6;
  assign CLBLM_R_X13Y158_SLICE_X19Y158_AMUX = CLBLM_R_X13Y158_SLICE_X19Y158_AO6;
  assign CLBLM_R_X13Y158_SLICE_X19Y158_BMUX = CLBLM_R_X13Y158_SLICE_X19Y158_BO6;
  assign CLBLM_R_X13Y159_SLICE_X18Y159_A = CLBLM_R_X13Y159_SLICE_X18Y159_AO6;
  assign CLBLM_R_X13Y159_SLICE_X18Y159_B = CLBLM_R_X13Y159_SLICE_X18Y159_BO6;
  assign CLBLM_R_X13Y159_SLICE_X18Y159_C = CLBLM_R_X13Y159_SLICE_X18Y159_CO6;
  assign CLBLM_R_X13Y159_SLICE_X18Y159_D = CLBLM_R_X13Y159_SLICE_X18Y159_DO6;
  assign CLBLM_R_X13Y159_SLICE_X19Y159_A = CLBLM_R_X13Y159_SLICE_X19Y159_AO6;
  assign CLBLM_R_X13Y159_SLICE_X19Y159_B = CLBLM_R_X13Y159_SLICE_X19Y159_BO6;
  assign CLBLM_R_X13Y159_SLICE_X19Y159_C = CLBLM_R_X13Y159_SLICE_X19Y159_CO6;
  assign CLBLM_R_X13Y159_SLICE_X19Y159_D = CLBLM_R_X13Y159_SLICE_X19Y159_DO6;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_A = CLBLM_R_X103Y141_SLICE_X162Y141_AO6;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_B = CLBLM_R_X103Y141_SLICE_X162Y141_BO6;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_C = CLBLM_R_X103Y141_SLICE_X162Y141_CO6;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_D = CLBLM_R_X103Y141_SLICE_X162Y141_DO6;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_A = CLBLM_R_X103Y141_SLICE_X163Y141_AO6;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_B = CLBLM_R_X103Y141_SLICE_X163Y141_BO6;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_C = CLBLM_R_X103Y141_SLICE_X163Y141_CO6;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_D = CLBLM_R_X103Y141_SLICE_X163Y141_DO6;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_AMUX = CLBLM_R_X103Y141_SLICE_X163Y141_AO5;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A = CLBLM_R_X103Y169_SLICE_X162Y169_AO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B = CLBLM_R_X103Y169_SLICE_X162Y169_BO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C = CLBLM_R_X103Y169_SLICE_X162Y169_CO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D = CLBLM_R_X103Y169_SLICE_X162Y169_DO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B = CLBLM_R_X103Y169_SLICE_X163Y169_BO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C = CLBLM_R_X103Y169_SLICE_X163Y169_CO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D = CLBLM_R_X103Y169_SLICE_X163Y169_DO6;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_AMUX = CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A = CLBLM_R_X103Y172_SLICE_X162Y172_AO6;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B = CLBLM_R_X103Y172_SLICE_X162Y172_BO6;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C = CLBLM_R_X103Y172_SLICE_X162Y172_CO6;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D = CLBLM_R_X103Y172_SLICE_X162Y172_DO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A = CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B = CLBLM_R_X103Y172_SLICE_X163Y172_BO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C = CLBLM_R_X103Y172_SLICE_X163Y172_CO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D = CLBLM_R_X103Y172_SLICE_X163Y172_DO6;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_AMUX = CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A = CLBLM_R_X103Y174_SLICE_X162Y174_AO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B = CLBLM_R_X103Y174_SLICE_X162Y174_BO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C = CLBLM_R_X103Y174_SLICE_X162Y174_CO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D = CLBLM_R_X103Y174_SLICE_X162Y174_DO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B = CLBLM_R_X103Y174_SLICE_X163Y174_BO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C = CLBLM_R_X103Y174_SLICE_X163Y174_CO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D = CLBLM_R_X103Y174_SLICE_X163Y174_DO6;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_AMUX = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A = CLBLM_R_X103Y177_SLICE_X162Y177_AO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B = CLBLM_R_X103Y177_SLICE_X162Y177_BO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C = CLBLM_R_X103Y177_SLICE_X162Y177_CO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D = CLBLM_R_X103Y177_SLICE_X162Y177_DO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B = CLBLM_R_X103Y177_SLICE_X163Y177_BO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C = CLBLM_R_X103Y177_SLICE_X163Y177_CO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D = CLBLM_R_X103Y177_SLICE_X163Y177_DO6;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_AMUX = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_O = LIOB33_X0Y51_IOB_X0Y51_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_O = LIOB33_X0Y53_IOB_X0Y53_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_O = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_O = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_O = LIOB33_X0Y65_IOB_X0Y65_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_O = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_O = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_O = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_O = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_O = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_X0Y73_ILOGIC_X0Y73_O = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_O = LIOB33_X0Y75_IOB_X0Y76_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_O = LIOB33_X0Y75_IOB_X0Y75_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_O = LIOB33_X0Y77_IOB_X0Y78_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_O = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_O = LIOB33_X0Y79_IOB_X0Y79_I;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_OQ = CLBLL_L_X2Y140_SLICE_X0Y140_AO6;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_OQ = CLBLL_L_X2Y139_SLICE_X0Y139_AO5;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_TQ = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_OQ = CLBLL_L_X2Y139_SLICE_X0Y139_AO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_OQ = CLBLL_L_X2Y139_SLICE_X0Y139_BO5;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_TQ = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_OQ = CLBLL_L_X2Y139_SLICE_X0Y139_BO6;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_OQ = CLBLL_L_X2Y140_SLICE_X0Y140_BO5;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_TQ = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_OQ = CLBLL_L_X2Y140_SLICE_X0Y140_BO6;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_OQ = CLBLM_R_X3Y142_SLICE_X3Y142_BO6;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_TQ = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_OQ = CLBLM_R_X3Y142_SLICE_X3Y142_DO6;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_OQ = CLBLM_L_X12Y151_SLICE_X16Y151_C5Q;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_TQ = 1'b1;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_OQ = 1'b0;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_OQ = CLBLM_R_X11Y144_SLICE_X15Y144_AQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_TQ = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_OQ = CLBLM_L_X12Y151_SLICE_X16Y151_CQ;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_OQ = CLBLM_R_X5Y148_SLICE_X7Y148_BQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_TQ = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_OQ = CLBLM_R_X5Y147_SLICE_X7Y147_CQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = CLBLL_L_X4Y149_SLICE_X5Y149_A5Q;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = CLBLM_R_X11Y144_SLICE_X15Y144_A5Q;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = CLBLM_R_X5Y148_SLICE_X7Y148_B5Q;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = CLBLM_L_X8Y146_SLICE_X10Y146_B5Q;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_OQ = CLBLL_L_X4Y147_SLICE_X5Y147_AQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_OQ = CLBLM_L_X8Y154_SLICE_X10Y154_C5Q;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_OQ = CLBLM_R_X3Y151_SLICE_X2Y151_AQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_OQ = CLBLL_L_X4Y152_SLICE_X4Y152_AQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_OQ = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_OQ = CLBLL_L_X4Y151_SLICE_X5Y151_CQ;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_OQ = CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_OQ = CLBLM_R_X5Y146_SLICE_X6Y146_A5Q;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_OQ = CLBLM_R_X5Y146_SLICE_X6Y146_AQ;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = CLBLM_R_X5Y144_SLICE_X6Y144_AQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_OQ = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_OQ = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_OQ = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_OQ = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_OQ = LIOB33_X0Y61_IOB_X0Y61_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_OQ = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_OQ = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_TQ = 1'b1;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_OQ = LIOB33_X0Y65_IOB_X0Y65_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_OQ = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_TQ = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_OQ = LIOB33_X0Y67_IOB_X0Y67_I;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_OQ = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_TQ = 1'b1;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_OQ = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_OQ = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_TQ = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_OQ = RIOB33_X105Y117_IOB_X1Y117_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_OQ = RIOB33_X105Y109_IOB_X1Y109_I;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_TQ = 1'b1;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_OQ = RIOB33_X105Y107_IOB_X1Y108_I;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_OQ = RIOB33_X105Y113_IOB_X1Y113_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_TQ = 1'b1;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_OQ = RIOB33_X105Y111_IOB_X1Y112_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_OQ = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_TQ = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_OQ = RIOB33_X105Y113_IOB_X1Y114_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_OQ = CLBLM_R_X103Y141_SLICE_X163Y141_AO6;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_TQ = 1'b1;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_OQ = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_OQ = CLBLM_L_X10Y163_SLICE_X13Y163_AO6;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_TQ = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_OQ = CLBLM_R_X103Y141_SLICE_X163Y141_AO5;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_OQ = RIOB33_X105Y127_IOB_X1Y128_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_TQ = 1'b1;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_OQ = RIOB33_X105Y127_IOB_X1Y127_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_OQ = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_TQ = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_OQ = RIOB33_X105Y129_IOB_X1Y129_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_OQ = RIOB33_X105Y131_IOB_X1Y132_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_TQ = 1'b1;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_OQ = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_OQ = RIOB33_X105Y135_IOB_X1Y136_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_TQ = 1'b1;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_OQ = RIOB33_X105Y135_IOB_X1Y135_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_OQ = RIOB33_X105Y143_IOB_X1Y143_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_TQ = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_OQ = RIOB33_X105Y137_IOB_X1Y137_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_OQ = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_TQ = 1'b1;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_OQ = RIOB33_X105Y145_IOB_X1Y146_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_OQ = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_TQ = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_OQ = RIOB33_X105Y147_IOB_X1Y148_I;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_OQ = LIOB33_X0Y69_IOB_X0Y69_I;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_TQ = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_OQ = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_OQ = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_TQ = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_OQ = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_TQ = 1'b1;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_OQ = CLBLL_L_X2Y140_SLICE_X0Y140_AO5;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_TQ = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ = 1'b1;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_OQ = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_TQ = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_OQ = LIOB33_X0Y73_IOB_X0Y74_I;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_O = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_O = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_O = LIOB33_X0Y69_IOB_X0Y69_I;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_OQ = CLBLM_R_X3Y151_SLICE_X3Y151_BO6;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_OQ = CLBLM_R_X3Y142_SLICE_X3Y142_CO6;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = CLBLM_L_X12Y149_SLICE_X16Y149_BQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = CLBLM_R_X11Y149_SLICE_X15Y149_AQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ = CLBLM_L_X10Y144_SLICE_X12Y144_AO5;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ = LIOB33_X0Y57_IOB_X0Y57_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ = LIOB33_X0Y55_IOB_X0Y55_I;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_OQ = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_OQ = RIOB33_X105Y115_IOB_X1Y115_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_OQ = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_OQ = RIOB33_X105Y121_IOB_X1Y122_I;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_OQ = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_OQ = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_OQ = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_OQ = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_O = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_OQ = CLBLM_L_X8Y146_SLICE_X10Y146_BQ;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_OQ = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = CLBLM_R_X5Y146_SLICE_X6Y146_BQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = CLBLM_R_X5Y144_SLICE_X6Y144_BQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_OQ = RIOB33_X105Y111_IOB_X1Y111_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_OQ = RIOB33_X105Y109_IOB_X1Y110_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_OQ = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_OQ = RIOB33_X105Y143_IOB_X1Y144_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_TQ = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_O = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_O = RIOB33_X105Y123_IOB_X1Y124_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_O = RIOB33_X105Y135_IOB_X1Y136_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_O = RIOB33_X105Y135_IOB_X1Y135_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_O = RIOB33_X105Y139_IOB_X1Y140_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_O = RIOB33_X105Y139_IOB_X1Y139_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_O = RIOB33_X105Y141_IOB_X1Y142_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_O = RIOB33_X105Y141_IOB_X1Y141_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_O = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_O = RIOB33_X105Y145_IOB_X1Y145_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_O = RIOB33_X105Y147_IOB_X1Y148_I;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_O = RIOB33_X105Y147_IOB_X1Y147_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_OQ = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_TQ = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_OQ = LIOB33_X0Y75_IOB_X0Y76_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_OQ = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_TQ = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_OQ = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_OQ = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_TQ = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_OQ = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_OQ = CLBLM_R_X13Y155_SLICE_X18Y155_CO6;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_TQ = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_OQ = CLBLM_R_X13Y154_SLICE_X18Y154_DO6;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_OQ = CLBLM_L_X12Y155_SLICE_X17Y155_DO6;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_TQ = 1'b1;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_OQ = CLBLM_R_X13Y155_SLICE_X18Y155_CO5;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_OQ = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_TQ = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_OQ = RIOB33_X105Y125_IOB_X1Y125_I;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_OQ = CLBLM_L_X10Y163_SLICE_X13Y163_AO6;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_TQ = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_OQ = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_OQ = CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_TQ = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_OQ = CLBLM_L_X12Y159_SLICE_X16Y159_CO6;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_OQ = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_TQ = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_OQ = CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_OQ = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_TQ = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_OQ = CLBLM_R_X13Y157_SLICE_X18Y157_AO5;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_TQ = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_OQ = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_OQ = CLBLM_R_X13Y154_SLICE_X18Y154_DO6;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_TQ = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_OQ = CLBLM_L_X12Y159_SLICE_X16Y159_AO5;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_OQ = CLBLM_L_X12Y155_SLICE_X17Y155_DO5;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_TQ = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_OQ = CLBLM_L_X12Y155_SLICE_X17Y155_DO6;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_OQ = CLBLM_R_X13Y154_SLICE_X18Y154_AQ;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_TQ = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_OQ = CLBLM_R_X7Y149_SLICE_X9Y149_DO5;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_OQ = CLBLM_R_X13Y156_SLICE_X18Y156_AQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_TQ = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_OQ = CLBLM_L_X12Y159_SLICE_X16Y159_BQ;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_OQ = CLBLM_R_X13Y153_SLICE_X19Y153_BQ;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_TQ = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_OQ = CLBLM_L_X12Y156_SLICE_X16Y156_BQ;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_OQ = CLBLM_L_X12Y159_SLICE_X16Y159_AQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_TQ = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_OQ = CLBLM_R_X13Y157_SLICE_X18Y157_AQ;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_OQ = CLBLM_L_X16Y156_SLICE_X22Y156_AO5;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_TQ = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_OQ = CLBLM_L_X16Y156_SLICE_X22Y156_AO5;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_TQ = 1'b1;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_OQ = LIOB33_X0Y75_IOB_X0Y75_I;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_TQ = 1'b1;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_OQ = CLBLM_R_X13Y156_SLICE_X19Y156_AQ;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_O = RIOB33_X105Y119_IOB_X1Y119_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_O = RIOB33_X105Y131_IOB_X1Y131_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_O = RIOB33_X105Y143_IOB_X1Y144_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_O = RIOB33_X105Y143_IOB_X1Y143_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_OQ = CLBLL_L_X36Y150_SLICE_X54Y150_AO6;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_OQ = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_OQ = CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_OQ = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_OQ = CLBLM_R_X13Y155_SLICE_X18Y155_CO5;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_OQ = CLBLM_R_X13Y155_SLICE_X18Y155_CO6;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_OQ = CLBLM_R_X13Y156_SLICE_X19Y156_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_OQ = CLBLM_L_X12Y156_SLICE_X16Y156_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_O = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_O = RIOB33_X105Y137_IOB_X1Y137_I;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_OQ = CLBLM_R_X7Y149_SLICE_X9Y149_DO5;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_OQ = CLBLM_L_X12Y155_SLICE_X17Y155_DO5;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_OQ = CLBLM_R_X11Y156_SLICE_X15Y156_BQ;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_OQ = CLBLM_L_X12Y155_SLICE_X16Y155_AQ;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_TQ = 1'b1;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_T1 = 1'b1;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_D1 = CLBLM_L_X10Y154_SLICE_X12Y154_A5Q;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_D2 = CLBLM_L_X10Y155_SLICE_X13Y155_AQ;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_D3 = 1'b1;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_D4 = CLBLM_L_X8Y158_SLICE_X10Y158_BQ;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_D5 = 1'b1;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_D6 = CLBLM_L_X10Y154_SLICE_X13Y154_C5Q;
  assign LIOB33_X0Y147_IOB_X0Y147_O = LIOB33_X0Y71_IOB_X0Y71_I;
  assign LIOB33_X0Y147_IOB_X0Y148_O = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLM_R_X13Y159_SLICE_X19Y159_A1 = 1'b1;
  assign CLBLM_R_X13Y159_SLICE_X19Y159_A2 = 1'b1;
  assign CLBLM_R_X13Y159_SLICE_X19Y159_A3 = 1'b1;
  assign CLBLM_R_X13Y159_SLICE_X19Y159_A4 = 1'b1;
  assign CLBLM_R_X13Y159_SLICE_X19Y159_A5 = 1'b1;
  assign CLBLM_R_X13Y159_SLICE_X19Y159_A6 = 1'b1;
  assign CLBLM_R_X13Y159_SLICE_X19Y159_B1 = 1'b1;
  assign CLBLM_R_X13Y159_SLICE_X19Y159_B2 = 1'b1;
  assign CLBLM_R_X13Y159_SLICE_X19Y159_B3 = 1'b1;
  assign CLBLM_R_X13Y159_SLICE_X19Y159_B4 = 1'b1;
  assign CLBLM_R_X13Y159_SLICE_X19Y159_B5 = 1'b1;
  assign CLBLM_R_X13Y159_SLICE_X19Y159_B6 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A1 = CLBLM_R_X13Y149_SLICE_X18Y149_CQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A3 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_A6 = 1'b1;
  assign CLBLM_R_X13Y159_SLICE_X19Y159_C1 = 1'b1;
  assign CLBLM_R_X13Y159_SLICE_X19Y159_C2 = 1'b1;
  assign CLBLM_R_X13Y159_SLICE_X19Y159_C3 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B1 = CLBLM_L_X10Y149_SLICE_X13Y149_A5Q;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B2 = CLBLM_R_X13Y155_SLICE_X19Y155_AO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B3 = CLBLM_R_X5Y155_SLICE_X6Y155_DO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B4 = CLBLM_R_X13Y153_SLICE_X18Y153_AQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B5 = CLBLM_L_X10Y153_SLICE_X13Y153_AQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_B6 = CLBLM_R_X11Y149_SLICE_X15Y149_CO6;
  assign CLBLM_R_X13Y159_SLICE_X19Y159_D1 = 1'b1;
  assign CLBLM_R_X13Y159_SLICE_X19Y159_D2 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C1 = CLBLM_L_X10Y151_SLICE_X12Y151_AQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C2 = CLBLM_R_X11Y150_SLICE_X15Y150_CO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C3 = CLBLM_R_X7Y148_SLICE_X9Y148_BQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C4 = CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C5 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A1 = CLBLM_R_X7Y155_SLICE_X9Y155_A5Q;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A2 = CLBLM_L_X12Y149_SLICE_X16Y149_AQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A3 = CLBLL_L_X4Y155_SLICE_X4Y155_AQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A4 = CLBLL_L_X4Y155_SLICE_X4Y155_BQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_A6 = CLBLL_L_X4Y149_SLICE_X4Y149_AQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_C6 = CLBLM_R_X11Y149_SLICE_X14Y149_BQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B1 = CLBLL_L_X4Y152_SLICE_X4Y152_DO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B2 = CLBLL_L_X4Y152_SLICE_X5Y152_DO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B3 = CLBLM_R_X3Y151_SLICE_X2Y151_CO5;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B4 = CLBLM_R_X5Y152_SLICE_X6Y152_DO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B5 = CLBLM_R_X7Y153_SLICE_X9Y153_BQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_B6 = CLBLL_L_X4Y152_SLICE_X4Y152_CO6;
  assign CLBLM_L_X10Y163_SLICE_X13Y163_C3 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D1 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D2 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C1 = CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C2 = CLBLL_L_X2Y155_SLICE_X1Y155_CO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C3 = CLBLM_R_X3Y158_SLICE_X2Y158_AO5;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_C6 = CLBLL_L_X2Y155_SLICE_X1Y155_CO5;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A1 = CLBLM_R_X13Y151_SLICE_X18Y151_AQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A3 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A5 = CLBLM_L_X10Y147_SLICE_X12Y147_BQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_A6 = CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D1 = CLBLL_L_X4Y157_SLICE_X4Y157_CO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D3 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D4 = CLBLL_L_X2Y155_SLICE_X1Y155_CO6;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D5 = CLBLM_R_X5Y149_SLICE_X6Y149_BQ;
  assign CLBLL_L_X4Y152_SLICE_X4Y152_D6 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B3 = CLBLM_R_X11Y148_SLICE_X14Y148_AQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B4 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C1 = CLBLM_L_X12Y150_SLICE_X17Y150_AQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C2 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C3 = CLBLM_R_X11Y149_SLICE_X14Y149_DQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C4 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C5 = CLBLM_L_X10Y148_SLICE_X13Y148_DO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y159_SLICE_X18Y159_D4 = CLBLM_L_X12Y158_SLICE_X16Y158_AQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y159_SLICE_X18Y159_D6 = CLBLM_L_X8Y154_SLICE_X10Y154_AQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D1 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D2 = CLBLM_L_X10Y148_SLICE_X13Y148_DO6;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D3 = CLBLM_R_X11Y149_SLICE_X14Y149_DQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D4 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_D6 = CLBLM_R_X13Y152_SLICE_X19Y152_AQ;
  assign RIOB33_SING_X105Y150_IOB_X1Y150_O = LIOB33_X0Y75_IOB_X0Y75_I;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_D1 = CLBLM_R_X13Y155_SLICE_X18Y155_CO5;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A1 = CLBLL_L_X4Y151_SLICE_X4Y151_BQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A2 = CLBLL_L_X4Y148_SLICE_X5Y148_CQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A3 = CLBLL_L_X4Y152_SLICE_X5Y152_AQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A5 = CLBLM_L_X10Y151_SLICE_X12Y151_CQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_A6 = CLBLM_L_X10Y148_SLICE_X13Y148_BQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B1 = CLBLM_R_X5Y152_SLICE_X6Y152_CO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B2 = CLBLL_L_X4Y152_SLICE_X5Y152_BQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B3 = CLBLM_R_X5Y150_SLICE_X6Y150_AQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B4 = CLBLM_R_X7Y152_SLICE_X9Y152_AQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_B6 = 1'b1;
  assign CLBLM_L_X10Y163_SLICE_X13Y163_D2 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y182_T1 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C2 = CLBLL_L_X4Y152_SLICE_X5Y152_CQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C3 = 1'b1;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C4 = CLBLL_L_X4Y151_SLICE_X5Y151_BQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C5 = CLBLL_L_X4Y147_SLICE_X4Y147_BO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_C6 = CLBLM_L_X8Y153_SLICE_X11Y153_C5Q;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_D1 = CLBLM_R_X13Y155_SLICE_X18Y155_CO6;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D1 = CLBLM_R_X5Y149_SLICE_X7Y149_BQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D2 = CLBLM_R_X3Y156_SLICE_X3Y156_AO5;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D3 = CLBLL_L_X4Y148_SLICE_X5Y148_CQ;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D5 = CLBLL_L_X4Y157_SLICE_X4Y157_CO5;
  assign CLBLL_L_X4Y152_SLICE_X5Y152_D6 = CLBLL_L_X4Y157_SLICE_X5Y157_AO6;
  assign RIOI3_TBYTESRC_X105Y181_OLOGIC_X1Y181_T1 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_A1 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_A2 = CLBLM_R_X7Y148_SLICE_X8Y148_BQ;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_A3 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_A4 = CLBLM_R_X7Y148_SLICE_X8Y148_AQ;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_A5 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_A6 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_B2 = CLBLM_L_X8Y158_SLICE_X11Y158_AQ;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_B4 = CLBLM_L_X10Y153_SLICE_X13Y153_CQ;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_B5 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_B6 = CLBLM_L_X12Y152_SLICE_X16Y152_AO5;
  assign CLBLM_L_X10Y163_SLICE_X12Y163_A5 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A2 = CLBLM_L_X8Y154_SLICE_X11Y154_BQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A3 = CLBLM_L_X8Y146_SLICE_X11Y146_AQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A4 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A5 = CLBLM_L_X10Y146_SLICE_X12Y146_AQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_A6 = CLBLM_R_X7Y146_SLICE_X9Y146_DO6;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_C1 = CLBLM_L_X10Y157_SLICE_X12Y157_BQ;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_C2 = CLBLM_L_X12Y157_SLICE_X16Y157_CQ;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_C3 = CLBLM_R_X11Y156_SLICE_X15Y156_AQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B2 = CLBLM_L_X8Y146_SLICE_X11Y146_BQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B3 = CLBLM_L_X8Y148_SLICE_X11Y148_AQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B4 = CLBLM_R_X7Y146_SLICE_X9Y146_AQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B5 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_B6 = CLBLM_R_X7Y146_SLICE_X8Y146_DO6;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_D1 = CLBLM_L_X10Y156_SLICE_X13Y156_BQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C1 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C2 = CLBLM_L_X8Y146_SLICE_X11Y146_CQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C3 = CLBLM_L_X8Y146_SLICE_X11Y146_BQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C4 = CLBLM_R_X7Y146_SLICE_X8Y146_DO6;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_C6 = CLBLM_L_X8Y146_SLICE_X10Y146_BQ;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_D3 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_D4 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_A1 = CLBLM_R_X11Y154_SLICE_X15Y154_CO5;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_A2 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_A5 = CLBLM_R_X7Y159_SLICE_X8Y159_AQ;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D1 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D2 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D3 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D4 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D5 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X11Y146_D6 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_A6 = CLBLM_L_X10Y155_SLICE_X12Y155_CQ;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_B1 = CLBLM_L_X10Y156_SLICE_X12Y156_DO6;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_B2 = CLBLM_L_X10Y156_SLICE_X13Y156_DO6;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_B3 = CLBLM_L_X10Y156_SLICE_X12Y156_AQ;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_B4 = CLBLM_L_X10Y153_SLICE_X13Y153_CQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A1 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A3 = CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A5 = CLBLM_L_X8Y150_SLICE_X11Y150_BQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_A6 = CLBLM_R_X11Y146_SLICE_X14Y146_CQ;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_C1 = CLBLM_L_X8Y155_SLICE_X11Y155_CQ;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_C2 = CLBLM_L_X8Y156_SLICE_X10Y156_CQ;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_C3 = CLBLM_L_X10Y154_SLICE_X12Y154_DQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B1 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B2 = CLBLM_R_X7Y154_SLICE_X9Y154_BQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B3 = CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_B6 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_D1 = CLBLM_L_X8Y153_SLICE_X11Y153_CQ;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_D2 = CLBLM_L_X12Y149_SLICE_X16Y149_CQ;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C1 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C2 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C3 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C4 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C5 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_C6 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_D3 = CLBLM_R_X13Y150_SLICE_X18Y150_AQ;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_D6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X13Y157_SLICE_X19Y157_D5 = 1'b1;
  assign CLBLM_R_X13Y157_SLICE_X19Y157_D6 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D1 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D2 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D3 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D4 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D5 = 1'b1;
  assign CLBLM_L_X8Y146_SLICE_X10Y146_D6 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A1 = CLBLM_R_X11Y149_SLICE_X15Y149_A5Q;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A4 = CLBLM_L_X12Y150_SLICE_X16Y150_AQ;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A5 = CLBLM_R_X11Y150_SLICE_X14Y150_AQ;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_A6 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B1 = CLBLM_R_X11Y150_SLICE_X14Y150_CO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B2 = CLBLM_L_X10Y149_SLICE_X12Y149_DO5;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B3 = CLBLM_R_X13Y148_SLICE_X18Y148_AQ;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B4 = CLBLM_R_X13Y149_SLICE_X19Y149_AQ;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B5 = CLBLM_R_X13Y150_SLICE_X18Y150_CQ;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_B6 = CLBLL_L_X4Y157_SLICE_X4Y157_BO6;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_A5 = CLBLM_L_X12Y156_SLICE_X16Y156_AQ;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_A1 = CLBLL_L_X4Y153_SLICE_X4Y153_DO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_A2 = CLBLL_L_X4Y154_SLICE_X4Y154_DO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_A3 = CLBLM_R_X5Y156_SLICE_X7Y156_DO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_A4 = CLBLM_R_X3Y151_SLICE_X2Y151_DO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_A5 = CLBLM_R_X3Y155_SLICE_X3Y155_DO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_A6 = CLBLM_R_X5Y153_SLICE_X6Y153_CO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C1 = CLBLM_R_X13Y150_SLICE_X19Y150_AQ;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C2 = CLBLM_R_X11Y155_SLICE_X14Y155_BQ;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C3 = CLBLM_R_X7Y149_SLICE_X8Y149_BQ;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_B1 = CLBLM_R_X3Y154_SLICE_X3Y154_DO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_B2 = CLBLM_R_X3Y155_SLICE_X2Y155_DO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_B3 = CLBLM_R_X5Y153_SLICE_X6Y153_DO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_B4 = CLBLM_R_X5Y154_SLICE_X7Y154_CO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_B5 = CLBLL_L_X4Y152_SLICE_X5Y152_DO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_B6 = CLBLL_L_X4Y153_SLICE_X4Y153_CO6;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D1 = CLBLM_L_X8Y147_SLICE_X11Y147_BQ;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D2 = 1'b1;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_C1 = CLBLM_R_X5Y149_SLICE_X6Y149_BQ;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_C2 = CLBLM_R_X3Y152_SLICE_X3Y152_AO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_C3 = CLBLL_L_X2Y153_SLICE_X1Y153_AO5;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_C4 = CLBLM_R_X3Y151_SLICE_X2Y151_CO5;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_C5 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_C6 = CLBLM_R_X7Y153_SLICE_X9Y153_BQ;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D3 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D4 = CLBLM_R_X13Y152_SLICE_X19Y152_AQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A2 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A3 = CLBLM_R_X11Y150_SLICE_X14Y150_AQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A4 = CLBLM_L_X12Y149_SLICE_X17Y149_A5Q;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A5 = CLBLM_L_X10Y150_SLICE_X12Y150_BQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_A6 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_D1 = CLBLL_L_X4Y153_SLICE_X5Y153_BO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_D2 = 1'b1;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_D3 = CLBLM_R_X3Y153_SLICE_X2Y153_CO6;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_D4 = CLBLM_R_X7Y155_SLICE_X9Y155_A5Q;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_D5 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign CLBLL_L_X4Y153_SLICE_X4Y153_D6 = CLBLM_R_X3Y153_SLICE_X2Y153_AO6;
  assign CLBLM_L_X10Y163_SLICE_X12Y163_D4 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B1 = CLBLM_R_X11Y150_SLICE_X14Y150_DO6;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B2 = CLBLM_R_X11Y149_SLICE_X15Y149_A5Q;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B3 = CLBLM_R_X5Y152_SLICE_X6Y152_BQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B4 = CLBLM_L_X10Y150_SLICE_X13Y150_AQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B5 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_B6 = CLBLM_L_X10Y152_SLICE_X12Y152_BQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C1 = CLBLM_R_X11Y146_SLICE_X15Y146_BQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C2 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C3 = CLBLM_R_X11Y146_SLICE_X14Y146_DQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C4 = CLBLL_L_X4Y148_SLICE_X5Y148_DQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C5 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_C6 = 1'b1;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_B4 = CLBLM_L_X12Y158_SLICE_X16Y158_BO5;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_B5 = CLBLM_L_X12Y156_SLICE_X17Y156_BQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_B6 = CLBLM_L_X8Y154_SLICE_X10Y154_AQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D1 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D2 = CLBLM_R_X7Y151_SLICE_X8Y151_DQ;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D3 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D4 = CLBLM_R_X11Y151_SLICE_X15Y151_AQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_A2 = 1'b1;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_A3 = CLBLL_L_X4Y150_SLICE_X4Y150_AQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_A5 = CLBLM_R_X5Y152_SLICE_X7Y152_DQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_A6 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D5 = 1'b1;
  assign CLBLM_R_X11Y150_SLICE_X14Y150_D6 = CLBLM_R_X5Y151_SLICE_X6Y151_CQ;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_A1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_A2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_B3 = CLBLL_L_X4Y157_SLICE_X4Y157_CO6;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_A3 = CLBLM_R_X3Y156_SLICE_X2Y156_DO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_B4 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_B5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_B6 = CLBLM_R_X7Y147_SLICE_X8Y147_AQ;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_A4 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_A5 = CLBLL_L_X4Y154_SLICE_X4Y154_BO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_C1 = CLBLM_R_X3Y154_SLICE_X3Y154_AO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_C2 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_A6 = 1'b1;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_C3 = CLBLM_R_X3Y157_SLICE_X2Y157_AO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_C4 = CLBLL_L_X4Y156_SLICE_X4Y156_CO6;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_C5 = CLBLM_R_X5Y150_SLICE_X6Y150_DQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_C6 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_B1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_B2 = CLBLL_L_X4Y154_SLICE_X5Y154_BO6;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_B3 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_B4 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_B5 = CLBLL_L_X4Y153_SLICE_X4Y153_AO6;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_B6 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_C1 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_C2 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_C3 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_C4 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_C5 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_C6 = 1'b1;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_D1 = CLBLL_L_X4Y150_SLICE_X4Y150_AQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_D2 = CLBLM_R_X5Y153_SLICE_X6Y153_BO5;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_D6 = CLBLM_R_X13Y153_SLICE_X18Y153_C5Q;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_D3 = CLBLL_L_X2Y155_SLICE_X1Y155_BO5;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_D4 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_D1 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_D2 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_D3 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_D4 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_D5 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X0Y139_D6 = 1'b1;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y157_SLICE_X13Y157_A1 = CLBLM_L_X8Y158_SLICE_X10Y158_AQ;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_A1 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_A2 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_A3 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_A4 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_A5 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_A6 = 1'b1;
  assign CLBLM_L_X10Y157_SLICE_X13Y157_A2 = CLBLM_R_X7Y148_SLICE_X8Y148_BQ;
  assign CLBLM_L_X10Y157_SLICE_X13Y157_A3 = CLBLM_R_X11Y156_SLICE_X15Y156_AQ;
  assign CLBLM_L_X10Y157_SLICE_X13Y157_A4 = CLBLM_R_X7Y148_SLICE_X8Y148_AQ;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_B1 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_B2 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_B3 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_B4 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_B5 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_B6 = 1'b1;
  assign CLBLM_L_X10Y157_SLICE_X13Y157_B1 = CLBLM_L_X8Y157_SLICE_X11Y157_DO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A1 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_C1 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_C2 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_C3 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_C4 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_C5 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_C6 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A2 = CLBLM_R_X5Y148_SLICE_X6Y148_BQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A3 = CLBLM_L_X8Y147_SLICE_X11Y147_AQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A5 = CLBLM_R_X11Y146_SLICE_X15Y146_AQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_A6 = CLBLM_R_X7Y146_SLICE_X9Y146_DO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B3 = CLBLM_L_X8Y148_SLICE_X11Y148_AQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B1 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B2 = CLBLM_L_X8Y147_SLICE_X11Y147_BQ;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_D1 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_D2 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_D3 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_D4 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_D5 = 1'b1;
  assign CLBLL_L_X2Y139_SLICE_X1Y139_D6 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C1 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C2 = CLBLM_R_X11Y147_SLICE_X14Y147_CO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C3 = CLBLM_R_X7Y147_SLICE_X9Y147_CQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C4 = CLBLM_R_X7Y147_SLICE_X9Y147_BQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C5 = CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_C6 = CLBLM_L_X8Y147_SLICE_X10Y147_BQ;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y157_SLICE_X12Y157_A1 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D1 = CLBLL_L_X4Y154_SLICE_X5Y154_BO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D2 = CLBLM_R_X3Y156_SLICE_X2Y156_DO6;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D3 = CLBLM_R_X3Y152_SLICE_X3Y152_BO5;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D4 = CLBLM_R_X7Y148_SLICE_X9Y148_CO5;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D5 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_D6 = CLBLM_R_X13Y155_SLICE_X19Y155_AO6;
  assign CLBLM_L_X10Y157_SLICE_X12Y157_A5 = CLBLM_L_X10Y155_SLICE_X12Y155_AQ;
  assign CLBLM_L_X10Y157_SLICE_X12Y157_A6 = CLBLM_L_X10Y150_SLICE_X12Y150_CQ;
  assign CLBLM_L_X10Y157_SLICE_X12Y157_B1 = CLBLM_L_X10Y159_SLICE_X12Y159_CO6;
  assign CLBLM_L_X10Y157_SLICE_X12Y157_B2 = CLBLM_L_X10Y157_SLICE_X13Y157_BO6;
  assign CLBLM_L_X10Y157_SLICE_X12Y157_B3 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A1 = CLBLM_L_X8Y147_SLICE_X10Y147_DO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A3 = CLBLM_L_X10Y154_SLICE_X13Y154_CQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A4 = CLBLM_L_X10Y148_SLICE_X13Y148_CQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_A6 = 1'b1;
  assign CLBLM_L_X10Y157_SLICE_X12Y157_C1 = 1'b1;
  assign CLBLM_L_X10Y157_SLICE_X12Y157_C2 = CLBLM_L_X10Y156_SLICE_X13Y156_CO6;
  assign CLBLM_L_X10Y157_SLICE_X12Y157_C3 = CLBLM_L_X10Y157_SLICE_X13Y157_DO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B1 = CLBLM_R_X7Y156_SLICE_X8Y156_BQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B2 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B4 = CLBLM_L_X8Y147_SLICE_X10Y147_DO5;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B5 = CLBLM_L_X8Y147_SLICE_X10Y147_BQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_B6 = CLBLM_L_X8Y147_SLICE_X10Y147_AO5;
  assign CLBLM_L_X10Y157_SLICE_X12Y157_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y157_SLICE_X12Y157_D1 = CLBLM_L_X10Y157_SLICE_X12Y157_CO5;
  assign CLBLM_L_X10Y157_SLICE_X12Y157_D4 = CLBLM_L_X10Y157_SLICE_X12Y157_CO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C1 = CLBLM_R_X5Y144_SLICE_X6Y144_BQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C2 = CLBLM_L_X8Y147_SLICE_X10Y147_CQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C3 = 1'b1;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C4 = CLBLM_R_X7Y151_SLICE_X9Y151_CQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y157_SLICE_X12Y157_D5 = CLBLM_L_X8Y157_SLICE_X11Y157_DO6;
  assign CLBLM_L_X10Y157_SLICE_X12Y157_D6 = CLBLM_L_X8Y156_SLICE_X11Y156_DO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D1 = CLBLM_L_X8Y147_SLICE_X10Y147_BQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D2 = CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D3 = CLBLM_R_X7Y147_SLICE_X9Y147_BQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D4 = CLBLM_R_X7Y146_SLICE_X9Y146_DO6;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D5 = CLBLM_R_X7Y147_SLICE_X9Y147_CQ;
  assign CLBLM_L_X8Y147_SLICE_X10Y147_D6 = 1'b1;
  assign CLBLM_R_X11Y159_SLICE_X14Y159_C4 = CLBLM_R_X11Y159_SLICE_X14Y159_BQ;
  assign LIOB33_X0Y155_IOB_X0Y156_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X11Y159_SLICE_X14Y159_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y159_SLICE_X14Y159_C6 = CLBLM_L_X12Y158_SLICE_X17Y158_AQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A1 = CLBLM_L_X12Y151_SLICE_X17Y151_A5Q;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A2 = CLBLM_L_X10Y147_SLICE_X12Y147_AQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A5 = CLBLM_L_X8Y154_SLICE_X10Y154_BQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_A6 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B1 = CLBLM_R_X11Y152_SLICE_X15Y152_DQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B2 = CLBLM_R_X11Y151_SLICE_X15Y151_BQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B3 = CLBLM_R_X13Y149_SLICE_X19Y149_CQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B4 = CLBLM_L_X12Y155_SLICE_X16Y155_CO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_A1 = CLBLM_R_X3Y155_SLICE_X3Y155_AO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_A2 = CLBLM_R_X7Y155_SLICE_X9Y155_DO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_A3 = CLBLM_R_X5Y156_SLICE_X6Y156_AO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_A4 = CLBLL_L_X4Y152_SLICE_X4Y152_BO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_A5 = CLBLM_R_X3Y154_SLICE_X3Y154_BO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_A6 = CLBLM_R_X5Y154_SLICE_X7Y154_CO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_B6 = CLBLM_L_X10Y150_SLICE_X12Y150_A5Q;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C1 = CLBLM_L_X12Y152_SLICE_X16Y152_BQ;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_B1 = CLBLM_R_X3Y153_SLICE_X3Y153_DO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_B2 = CLBLM_R_X3Y155_SLICE_X3Y155_DO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_B3 = CLBLL_L_X4Y156_SLICE_X5Y156_CO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_B4 = CLBLM_R_X3Y153_SLICE_X3Y153_CO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_B5 = CLBLM_R_X5Y154_SLICE_X6Y154_BO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_B6 = CLBLL_L_X4Y154_SLICE_X4Y154_CO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C3 = CLBLM_L_X10Y158_SLICE_X13Y158_BQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C4 = CLBLM_R_X7Y149_SLICE_X8Y149_CQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C6 = CLBLM_R_X11Y151_SLICE_X15Y151_DO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_C1 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_C2 = CLBLL_L_X4Y156_SLICE_X4Y156_CO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_C3 = CLBLL_L_X4Y155_SLICE_X4Y155_DO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_C4 = CLBLL_L_X4Y157_SLICE_X4Y157_BO5;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_C5 = CLBLM_R_X11Y151_SLICE_X15Y151_BQ;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_C6 = CLBLM_R_X7Y154_SLICE_X9Y154_BQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D1 = CLBLM_R_X7Y153_SLICE_X8Y153_BQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D2 = CLBLM_R_X11Y151_SLICE_X14Y151_CO6;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D3 = CLBLM_L_X10Y154_SLICE_X13Y154_BQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D4 = CLBLM_R_X13Y149_SLICE_X18Y149_CQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D5 = CLBLM_L_X12Y151_SLICE_X17Y151_BQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_D6 = CLBLM_R_X11Y151_SLICE_X14Y151_BQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A1 = CLBLM_R_X5Y151_SLICE_X7Y151_AQ;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_D1 = CLBLM_R_X3Y153_SLICE_X3Y153_AO6;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_D2 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_D3 = CLBLM_R_X3Y154_SLICE_X3Y154_AO5;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_D4 = CLBLM_L_X8Y154_SLICE_X11Y154_BQ;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_D5 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X4Y154_D6 = CLBLM_R_X11Y154_SLICE_X15Y154_AQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A3 = CLBLM_R_X11Y151_SLICE_X14Y151_AQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A4 = CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_A6 = CLBLM_R_X13Y152_SLICE_X19Y152_AQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B1 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B3 = CLBLM_L_X10Y153_SLICE_X13Y153_AQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B4 = CLBLM_L_X10Y149_SLICE_X12Y149_C5Q;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B5 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C1 = CLBLM_R_X7Y151_SLICE_X9Y151_C5Q;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C2 = CLBLM_L_X12Y152_SLICE_X17Y152_AQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C3 = CLBLM_L_X10Y151_SLICE_X13Y151_BQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C4 = CLBLM_L_X10Y151_SLICE_X13Y151_CQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C5 = CLBLM_L_X12Y151_SLICE_X17Y151_AQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_C6 = CLBLM_L_X10Y149_SLICE_X12Y149_C5Q;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_A2 = CLBLM_R_X5Y152_SLICE_X6Y152_CO5;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_A3 = CLBLL_L_X4Y154_SLICE_X5Y154_AQ;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_A4 = CLBLM_R_X7Y154_SLICE_X8Y154_AQ;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_A5 = CLBLM_R_X5Y152_SLICE_X7Y152_DQ;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_A6 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D1 = CLBLM_R_X7Y149_SLICE_X8Y149_BQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D2 = CLBLM_R_X11Y151_SLICE_X14Y151_AQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D3 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_A1 = CLBLM_R_X5Y155_SLICE_X6Y155_DO6;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_A2 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_A3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_A4 = CLBLM_R_X3Y155_SLICE_X2Y155_BO6;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_A5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_A6 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_B1 = CLBLM_R_X5Y154_SLICE_X6Y154_CO6;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_B2 = CLBLM_R_X3Y155_SLICE_X3Y155_DO6;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_B3 = CLBLL_L_X4Y153_SLICE_X5Y153_DO6;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_B1 = CLBLL_L_X4Y154_SLICE_X5Y154_CO6;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_B2 = CLBLL_L_X4Y153_SLICE_X4Y153_BO6;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_B3 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_B4 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_B6 = CLBLM_R_X3Y151_SLICE_X3Y151_CO6;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_B6 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_C1 = CLBLM_R_X3Y154_SLICE_X3Y154_CO6;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_C2 = CLBLL_L_X4Y153_SLICE_X5Y153_CO6;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_C3 = CLBLM_R_X5Y154_SLICE_X7Y154_DO6;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_C4 = CLBLM_R_X5Y154_SLICE_X6Y154_DO6;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_C5 = CLBLL_L_X4Y154_SLICE_X5Y154_DO6;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_C3 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_C4 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_D1 = CLBLM_R_X3Y153_SLICE_X3Y153_AO5;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_D2 = CLBLL_L_X4Y155_SLICE_X5Y155_A5Q;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_D3 = CLBLM_R_X3Y152_SLICE_X3Y152_AO6;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_D4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_D5 = CLBLM_R_X7Y154_SLICE_X8Y154_CQ;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_D6 = CLBLM_R_X11Y154_SLICE_X14Y154_D5Q;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_C6 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_C5 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_D1 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_D2 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_D3 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_D4 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_D5 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_D6 = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_D1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOI3_X0Y159_OLOGIC_X0Y160_T1 = 1'b1;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_D1 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_A1 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_A2 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_A3 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_A4 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_A5 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_A6 = 1'b1;
  assign CLBLM_L_X10Y158_SLICE_X13Y158_A1 = CLBLM_L_X8Y157_SLICE_X10Y157_CQ;
  assign CLBLM_L_X10Y158_SLICE_X13Y158_A2 = CLBLM_R_X11Y159_SLICE_X15Y159_DO5;
  assign CLBLM_L_X10Y158_SLICE_X13Y158_A3 = CLBLM_L_X10Y158_SLICE_X13Y158_AQ;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_B1 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_B2 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_B3 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_B4 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_B5 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_B6 = 1'b1;
  assign CLBLM_L_X10Y158_SLICE_X13Y158_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y158_SLICE_X13Y158_A5 = CLBLM_R_X11Y158_SLICE_X15Y158_BO6;
  assign CLBLM_L_X10Y158_SLICE_X13Y158_B5 = CLBLM_L_X10Y158_SLICE_X12Y158_AQ;
  assign CLBLM_L_X10Y158_SLICE_X13Y158_B6 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_C1 = 1'b1;
  assign CLBLM_L_X10Y158_SLICE_X13Y158_C1 = CLBLM_L_X10Y159_SLICE_X13Y159_AO6;
  assign CLBLM_L_X10Y158_SLICE_X13Y158_C2 = CLBLM_R_X11Y160_SLICE_X14Y160_AQ;
  assign CLBLM_L_X10Y158_SLICE_X13Y158_C3 = CLBLM_L_X10Y159_SLICE_X12Y159_DO6;
  assign CLBLM_L_X10Y158_SLICE_X13Y158_C4 = CLBLM_L_X8Y157_SLICE_X10Y157_BQ;
  assign CLBLM_L_X10Y158_SLICE_X13Y158_C5 = CLBLM_L_X8Y157_SLICE_X11Y157_DO6;
  assign CLBLM_L_X10Y158_SLICE_X13Y158_C6 = CLBLM_L_X8Y156_SLICE_X11Y156_DO6;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_C2 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_C3 = 1'b1;
  assign CLBLM_L_X10Y158_SLICE_X13Y158_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_C5 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_C6 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A3 = CLBLM_L_X8Y148_SLICE_X11Y148_AQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A4 = CLBLM_L_X10Y147_SLICE_X12Y147_BQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A6 = CLBLL_L_X4Y150_SLICE_X5Y150_DQ;
  assign CLBLM_L_X10Y158_SLICE_X13Y158_D1 = 1'b1;
  assign CLBLM_L_X10Y158_SLICE_X13Y158_D2 = 1'b1;
  assign CLBLM_L_X10Y158_SLICE_X13Y158_D3 = 1'b1;
  assign CLBLM_L_X10Y158_SLICE_X13Y158_D4 = 1'b1;
  assign CLBLM_L_X10Y158_SLICE_X13Y158_D5 = 1'b1;
  assign CLBLM_L_X10Y158_SLICE_X13Y158_D6 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_D2 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_D3 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_D5 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_D6 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C1 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C2 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C3 = CLBLM_L_X10Y148_SLICE_X13Y148_DO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C4 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C5 = CLBLM_R_X11Y149_SLICE_X14Y149_DQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_C6 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y158_SLICE_X12Y158_A1 = CLBLM_L_X10Y146_SLICE_X12Y146_BQ;
  assign CLBLM_L_X10Y158_SLICE_X12Y158_A2 = CLBLM_L_X10Y156_SLICE_X12Y156_BO6;
  assign CLBLM_L_X10Y158_SLICE_X12Y158_A3 = CLBLM_L_X10Y158_SLICE_X12Y158_AQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D3 = CLBLM_R_X7Y151_SLICE_X8Y151_BQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D4 = CLBLM_R_X11Y154_SLICE_X14Y154_DQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D5 = CLBLM_L_X8Y149_SLICE_X11Y149_BQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_D6 = 1'b1;
  assign CLBLM_L_X10Y158_SLICE_X12Y158_B1 = CLBLM_L_X10Y159_SLICE_X12Y159_CO6;
  assign CLBLM_L_X10Y158_SLICE_X12Y158_B2 = CLBLM_L_X10Y158_SLICE_X12Y158_BQ;
  assign CLBLM_L_X10Y158_SLICE_X12Y158_B3 = CLBLM_L_X10Y159_SLICE_X12Y159_DO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A1 = CLBLM_R_X11Y149_SLICE_X14Y149_DQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A2 = CLBLL_L_X4Y151_SLICE_X4Y151_BQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A3 = CLBLM_L_X8Y148_SLICE_X10Y148_AQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A4 = CLBLM_L_X12Y152_SLICE_X16Y152_B5Q;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_A6 = CLBLM_L_X10Y151_SLICE_X12Y151_CQ;
  assign CLBLM_L_X10Y158_SLICE_X12Y158_C1 = CLBLM_R_X11Y156_SLICE_X14Y156_BQ;
  assign CLBLM_L_X10Y158_SLICE_X12Y158_C2 = CLBLM_L_X8Y156_SLICE_X11Y156_DO6;
  assign CLBLM_L_X10Y158_SLICE_X12Y158_C3 = CLBLM_L_X8Y157_SLICE_X11Y157_DO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B1 = CLBLM_L_X8Y149_SLICE_X10Y149_BO5;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B2 = CLBLM_L_X8Y148_SLICE_X10Y148_BQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B3 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B5 = CLBLM_L_X8Y148_SLICE_X11Y148_CO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_B6 = CLBLM_L_X10Y151_SLICE_X12Y151_CQ;
  assign CLBLM_L_X10Y158_SLICE_X12Y158_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y158_SLICE_X12Y158_D1 = 1'b1;
  assign CLBLM_L_X10Y158_SLICE_X12Y158_D2 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C2 = CLBLM_L_X8Y148_SLICE_X10Y148_CQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C3 = CLBLM_L_X8Y146_SLICE_X10Y146_B5Q;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C4 = CLBLM_L_X8Y152_SLICE_X11Y152_CO6;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_C6 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X10Y158_SLICE_X12Y158_D4 = 1'b1;
  assign CLBLM_L_X10Y158_SLICE_X12Y158_D5 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D1 = CLBLM_L_X8Y148_SLICE_X11Y148_AQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D2 = CLBLM_L_X8Y147_SLICE_X10Y147_CQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D4 = CLBLM_R_X7Y151_SLICE_X9Y151_CQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D5 = CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  assign CLBLM_L_X8Y148_SLICE_X10Y148_D6 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_T1 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A1 = CLBLM_L_X10Y145_SLICE_X13Y145_AQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A2 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A3 = CLBLM_R_X11Y152_SLICE_X15Y152_AQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A4 = CLBLM_R_X11Y153_SLICE_X14Y153_BO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_A1 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_A3 = CLBLL_L_X4Y155_SLICE_X4Y155_AQ;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_A4 = CLBLM_R_X7Y155_SLICE_X8Y155_A5Q;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_A5 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_A6 = CLBLL_L_X4Y149_SLICE_X4Y149_CO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B4 = CLBLM_L_X8Y152_SLICE_X10Y152_AQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B5 = CLBLM_R_X13Y153_SLICE_X18Y153_BQ;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_B1 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_B2 = CLBLL_L_X4Y155_SLICE_X4Y155_BQ;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_B3 = CLBLM_R_X5Y153_SLICE_X6Y153_AQ;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_B4 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_B6 = CLBLL_L_X4Y149_SLICE_X4Y149_CO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D3 = 1'b1;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_C1 = CLBLM_R_X3Y151_SLICE_X3Y151_AQ;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_C2 = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_C3 = CLBLM_R_X3Y150_SLICE_X3Y150_AQ;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_C4 = CLBLL_L_X4Y156_SLICE_X4Y156_AQ;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_C5 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_C6 = CLBLM_L_X12Y155_SLICE_X16Y155_CO6;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D5 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y149_SLICE_X15Y149_D6 = CLBLL_L_X4Y149_SLICE_X5Y149_AQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D1 = CLBLM_L_X10Y152_SLICE_X13Y152_CO6;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D2 = CLBLM_L_X10Y148_SLICE_X13Y148_AQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D3 = CLBLM_R_X11Y152_SLICE_X15Y152_DQ;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_D1 = CLBLL_L_X4Y154_SLICE_X5Y154_AQ;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_D2 = CLBLM_R_X3Y158_SLICE_X2Y158_AO5;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_D3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_D4 = CLBLL_L_X2Y155_SLICE_X1Y155_CO6;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_D5 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X4Y155_D6 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A1 = CLBLM_R_X7Y153_SLICE_X9Y153_CO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A2 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A3 = CLBLM_R_X11Y152_SLICE_X14Y152_AQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A5 = CLBLM_L_X10Y150_SLICE_X13Y150_AQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_A6 = CLBLM_L_X8Y153_SLICE_X11Y153_CQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B1 = CLBLM_L_X12Y152_SLICE_X17Y152_A5Q;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B2 = CLBLM_L_X12Y152_SLICE_X16Y152_B5Q;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B3 = CLBLM_R_X11Y156_SLICE_X15Y156_AQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B5 = CLBLM_R_X5Y151_SLICE_X6Y151_AQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_B6 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C2 = CLBLM_R_X11Y152_SLICE_X14Y152_CQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C4 = CLBLM_L_X8Y152_SLICE_X10Y152_BQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C5 = CLBLM_L_X10Y152_SLICE_X12Y152_CO6;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_C6 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_A1 = CLBLM_R_X3Y156_SLICE_X2Y156_DO6;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_A3 = CLBLM_R_X11Y155_SLICE_X14Y155_BQ;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_A4 = CLBLM_R_X7Y155_SLICE_X9Y155_BQ;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_A5 = CLBLL_L_X4Y154_SLICE_X5Y154_CO6;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_A6 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D2 = CLBLM_L_X10Y158_SLICE_X13Y158_BQ;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_B1 = 1'b1;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_B2 = CLBLL_L_X4Y155_SLICE_X5Y155_BQ;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_B4 = CLBLL_L_X4Y146_SLICE_X5Y146_AQ;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_B5 = CLBLL_L_X4Y147_SLICE_X4Y147_BO6;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_B6 = CLBLL_L_X4Y155_SLICE_X5Y155_A5Q;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D3 = CLBLM_L_X8Y154_SLICE_X11Y154_CQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D4 = CLBLM_L_X10Y151_SLICE_X13Y151_BQ;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D5 = CLBLM_L_X12Y150_SLICE_X17Y150_AQ;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_C1 = CLBLL_L_X4Y155_SLICE_X5Y155_BQ;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_C2 = CLBLM_R_X3Y156_SLICE_X3Y156_AO5;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_C3 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_C4 = CLBLL_L_X4Y150_SLICE_X5Y150_CQ;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_C5 = CLBLL_L_X4Y157_SLICE_X4Y157_CO6;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_C6 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_D1 = CLBLM_R_X3Y158_SLICE_X2Y158_AO5;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_D2 = CLBLL_L_X2Y155_SLICE_X1Y155_CO6;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_D3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_D4 = CLBLL_L_X2Y155_SLICE_X1Y155_AO5;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_D5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X4Y155_SLICE_X5Y155_D6 = CLBLL_L_X4Y151_SLICE_X5Y151_BQ;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B1 = CLBLM_R_X7Y157_SLICE_X9Y157_BQ;
  assign LIOB33_X0Y157_IOB_X0Y158_O = RIOB33_X105Y115_IOB_X1Y116_I;
  assign LIOB33_X0Y157_IOB_X0Y157_O = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X11Y149_SLICE_X14Y149_B2 = CLBLM_R_X11Y149_SLICE_X14Y149_BQ;
  assign CLBLM_L_X10Y159_SLICE_X13Y159_A1 = CLBLM_L_X10Y158_SLICE_X12Y158_BQ;
  assign CLBLM_L_X10Y159_SLICE_X13Y159_A2 = CLBLM_R_X11Y155_SLICE_X14Y155_CQ;
  assign CLBLM_L_X10Y159_SLICE_X13Y159_A3 = CLBLM_L_X10Y157_SLICE_X12Y157_CO5;
  assign CLBLM_L_X10Y159_SLICE_X13Y159_A4 = CLBLM_L_X10Y156_SLICE_X13Y156_CO6;
  assign CLBLM_L_X10Y159_SLICE_X13Y159_A5 = CLBLM_R_X11Y156_SLICE_X14Y156_BQ;
  assign CLBLM_L_X10Y159_SLICE_X13Y159_A6 = 1'b1;
  assign CLBLM_L_X10Y159_SLICE_X13Y159_B1 = CLBLM_L_X10Y158_SLICE_X12Y158_BQ;
  assign CLBLM_L_X10Y159_SLICE_X13Y159_B2 = CLBLM_R_X11Y155_SLICE_X14Y155_CQ;
  assign CLBLM_L_X10Y159_SLICE_X13Y159_B3 = CLBLM_L_X10Y157_SLICE_X12Y157_CO5;
  assign CLBLM_L_X10Y159_SLICE_X13Y159_B4 = CLBLM_R_X11Y159_SLICE_X15Y159_BQ;
  assign CLBLM_L_X10Y159_SLICE_X13Y159_B5 = CLBLM_R_X11Y160_SLICE_X14Y160_AQ;
  assign CLBLM_L_X10Y159_SLICE_X13Y159_B6 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A1 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A2 = CLBLM_R_X5Y151_SLICE_X6Y151_CQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A3 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_A6 = CLBLM_R_X7Y150_SLICE_X9Y150_CO6;
  assign CLBLM_L_X10Y159_SLICE_X13Y159_C1 = CLBLM_L_X10Y159_SLICE_X13Y159_AO5;
  assign CLBLM_L_X10Y159_SLICE_X13Y159_C2 = CLBLM_L_X8Y157_SLICE_X10Y157_BQ;
  assign CLBLM_L_X10Y159_SLICE_X13Y159_C3 = CLBLM_R_X11Y160_SLICE_X14Y160_AQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B1 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B2 = CLBLM_L_X8Y149_SLICE_X11Y149_BQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B4 = CLBLL_L_X4Y150_SLICE_X5Y150_CQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_B6 = 1'b1;
  assign CLBLM_L_X10Y159_SLICE_X13Y159_D1 = CLBLM_L_X8Y158_SLICE_X11Y158_AQ;
  assign CLBLM_L_X10Y159_SLICE_X13Y159_D2 = CLBLM_L_X8Y156_SLICE_X11Y156_DO6;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C2 = CLBLM_L_X8Y149_SLICE_X11Y149_CQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C4 = CLBLM_R_X7Y147_SLICE_X9Y147_A5Q;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C5 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_C6 = CLBLM_L_X10Y147_SLICE_X13Y147_AQ;
  assign CLBLM_L_X10Y159_SLICE_X13Y159_D3 = CLBLM_R_X11Y160_SLICE_X14Y160_AQ;
  assign CLBLM_L_X10Y159_SLICE_X13Y159_D4 = CLBLM_L_X10Y159_SLICE_X13Y159_AO5;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y159_SLICE_X12Y159_A1 = CLBLM_R_X11Y159_SLICE_X14Y159_DQ;
  assign CLBLM_L_X10Y159_SLICE_X12Y159_A2 = CLBLM_L_X10Y159_SLICE_X13Y159_BO5;
  assign CLBLM_L_X10Y159_SLICE_X12Y159_A3 = CLBLM_R_X11Y160_SLICE_X14Y160_AQ;
  assign CLBLM_L_X10Y159_SLICE_X12Y159_A4 = CLBLM_L_X10Y159_SLICE_X13Y159_AO5;
  assign CLBLM_L_X10Y159_SLICE_X12Y159_A5 = CLBLM_R_X11Y159_SLICE_X15Y159_BQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D1 = CLBLM_L_X10Y148_SLICE_X13Y148_BQ;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D2 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D3 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D4 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D5 = 1'b1;
  assign CLBLM_L_X8Y149_SLICE_X11Y149_D6 = CLBLM_L_X10Y155_SLICE_X12Y155_BQ;
  assign CLBLM_L_X10Y159_SLICE_X12Y159_A6 = CLBLM_L_X8Y156_SLICE_X11Y156_DO6;
  assign CLBLM_L_X10Y159_SLICE_X12Y159_B1 = CLBLM_R_X11Y160_SLICE_X14Y160_AQ;
  assign CLBLM_L_X10Y159_SLICE_X12Y159_B2 = CLBLM_L_X10Y156_SLICE_X13Y156_CO6;
  assign CLBLM_L_X10Y159_SLICE_X12Y159_B3 = CLBLM_R_X11Y156_SLICE_X14Y156_BQ;
  assign CLBLM_L_X10Y159_SLICE_X12Y159_B4 = CLBLM_R_X11Y155_SLICE_X14Y155_CQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A1 = CLBLM_L_X8Y149_SLICE_X10Y149_BO5;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A3 = CLBLM_L_X8Y149_SLICE_X10Y149_AQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A4 = CLBLM_L_X8Y149_SLICE_X10Y149_BO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A5 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_A6 = CLBLM_L_X10Y155_SLICE_X12Y155_BQ;
  assign CLBLM_L_X10Y159_SLICE_X12Y159_C1 = 1'b1;
  assign CLBLM_L_X10Y159_SLICE_X12Y159_C2 = CLBLM_R_X11Y159_SLICE_X14Y159_DQ;
  assign CLBLM_L_X10Y159_SLICE_X12Y159_C3 = CLBLM_L_X10Y159_SLICE_X13Y159_BO5;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B1 = CLBLM_R_X11Y149_SLICE_X14Y149_DQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B2 = CLBLM_L_X8Y148_SLICE_X10Y148_BQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B3 = CLBLM_L_X8Y149_SLICE_X10Y149_AQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B4 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B5 = CLBLM_L_X10Y148_SLICE_X13Y148_DO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_B6 = 1'b1;
  assign CLBLM_L_X10Y159_SLICE_X12Y159_D1 = 1'b1;
  assign CLBLM_L_X10Y159_SLICE_X12Y159_D2 = CLBLM_R_X11Y159_SLICE_X14Y159_DQ;
  assign CLBLM_L_X10Y159_SLICE_X12Y159_D3 = CLBLM_L_X10Y159_SLICE_X13Y159_BO5;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C1 = CLBLM_L_X10Y150_SLICE_X13Y150_BQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C2 = CLBLM_L_X10Y148_SLICE_X13Y148_BQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C3 = CLBLM_L_X8Y155_SLICE_X10Y155_B5Q;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C4 = CLBLM_R_X7Y149_SLICE_X9Y149_C5Q;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C5 = CLBLM_L_X10Y148_SLICE_X13Y148_AQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_C6 = CLBLM_L_X10Y155_SLICE_X12Y155_BQ;
  assign CLBLM_L_X10Y159_SLICE_X12Y159_D4 = CLBLM_L_X8Y156_SLICE_X11Y156_DO6;
  assign CLBLM_L_X10Y159_SLICE_X12Y159_D5 = CLBLM_R_X7Y158_SLICE_X8Y158_CO5;
  assign CLBLM_L_X10Y159_SLICE_X12Y159_D6 = CLBLM_L_X10Y159_SLICE_X12Y159_BO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D1 = CLBLM_L_X10Y148_SLICE_X13Y148_DO6;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D2 = CLBLM_R_X11Y149_SLICE_X14Y149_DQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D3 = CLBLM_L_X8Y149_SLICE_X10Y149_AQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D4 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D5 = CLBLM_L_X8Y155_SLICE_X10Y155_B5Q;
  assign CLBLM_L_X8Y149_SLICE_X10Y149_D6 = CLBLM_L_X8Y148_SLICE_X10Y148_BQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A2 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A3 = CLBLM_R_X11Y153_SLICE_X15Y153_AQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A4 = CLBLM_L_X10Y152_SLICE_X12Y152_DO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_A1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_A3 = CLBLL_L_X4Y155_SLICE_X4Y155_CO6;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_A4 = CLBLL_L_X4Y154_SLICE_X5Y154_AQ;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_A5 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_A6 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_A6 = CLBLM_R_X11Y153_SLICE_X15Y153_DQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B1 = CLBLM_L_X8Y155_SLICE_X11Y155_CQ;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_B1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_B2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_B3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_B4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_B5 = CLBLL_L_X4Y157_SLICE_X4Y157_CO5;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_B6 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B4 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B6 = CLBLM_R_X7Y153_SLICE_X9Y153_CO6;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_C1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_C2 = CLBLM_R_X3Y158_SLICE_X2Y158_AO6;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_C3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_C4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_C6 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C3 = CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C6 = CLBLM_R_X13Y153_SLICE_X19Y153_AQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D2 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_D1 = CLBLM_L_X8Y154_SLICE_X11Y154_AQ;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_D2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_D3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_D4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_D5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y156_SLICE_X4Y156_D6 = CLBLL_L_X4Y157_SLICE_X4Y157_CO5;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D5 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D4 = CLBLM_R_X13Y153_SLICE_X19Y153_CQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A3 = CLBLM_R_X11Y153_SLICE_X14Y153_AQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A4 = CLBLM_R_X11Y153_SLICE_X14Y153_BO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A5 = CLBLM_L_X10Y148_SLICE_X13Y148_AQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_A6 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B2 = CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B3 = CLBLM_L_X8Y154_SLICE_X11Y154_CQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B4 = CLBLM_R_X13Y152_SLICE_X18Y152_BO5;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B5 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_B6 = CLBLM_L_X10Y151_SLICE_X13Y151_BQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_D6 = CLBLM_R_X7Y151_SLICE_X8Y151_DQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C1 = CLBLM_R_X13Y149_SLICE_X19Y149_AQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C2 = CLBLM_L_X8Y153_SLICE_X11Y153_BQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C3 = CLBLM_L_X12Y154_SLICE_X17Y154_A5Q;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C4 = CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C5 = CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_A1 = CLBLL_L_X4Y156_SLICE_X4Y156_CO5;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_A2 = CLBLL_L_X4Y155_SLICE_X5Y155_DO6;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_A3 = CLBLM_R_X3Y151_SLICE_X3Y151_AQ;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_A4 = CLBLM_R_X3Y156_SLICE_X2Y156_CO6;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_A5 = CLBLM_R_X5Y158_SLICE_X6Y158_CO6;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_A6 = CLBLM_R_X5Y157_SLICE_X6Y157_CO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_C6 = CLBLM_L_X8Y158_SLICE_X10Y158_BQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_B2 = CLBLL_L_X4Y157_SLICE_X4Y157_CO5;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_B3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_B4 = CLBLM_R_X7Y152_SLICE_X9Y152_AQ;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_B5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_B6 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D1 = CLBLM_L_X10Y152_SLICE_X13Y152_AQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D2 = CLBLM_L_X10Y150_SLICE_X13Y150_BQ;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D3 = CLBLM_L_X12Y152_SLICE_X17Y152_BO5;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_C1 = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_C2 = CLBLM_R_X3Y154_SLICE_X3Y154_AO6;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_C3 = CLBLL_L_X4Y157_SLICE_X5Y157_CO6;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_C4 = CLBLM_R_X7Y157_SLICE_X8Y157_DQ;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_C5 = CLBLL_L_X4Y156_SLICE_X4Y156_CO5;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_C6 = CLBLL_L_X4Y156_SLICE_X5Y156_BO6;
  assign LIOB33_X0Y159_IOB_X0Y160_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOB33_X0Y159_IOB_X0Y159_O = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_D1 = 1'b1;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_D2 = CLBLL_L_X2Y155_SLICE_X1Y155_CO6;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_D3 = CLBLL_L_X2Y155_SLICE_X1Y155_CO5;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_D4 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_D5 = CLBLL_L_X4Y157_SLICE_X4Y157_CO6;
  assign CLBLL_L_X4Y156_SLICE_X5Y156_D6 = CLBLM_R_X7Y156_SLICE_X8Y156_DQ;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A2 = CLBLM_L_X8Y146_SLICE_X11Y146_BQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A4 = CLBLM_R_X5Y152_SLICE_X7Y152_CQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A5 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_A6 = CLBLM_R_X11Y152_SLICE_X14Y152_DO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B1 = CLBLM_L_X8Y157_SLICE_X10Y157_BQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B2 = CLBLM_L_X8Y150_SLICE_X11Y150_BQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B3 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B4 = CLBLM_L_X8Y151_SLICE_X11Y151_BO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C1 = CLBLM_R_X7Y148_SLICE_X9Y148_CO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C2 = CLBLM_R_X7Y158_SLICE_X8Y158_CO5;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C3 = CLBLM_L_X8Y146_SLICE_X11Y146_AQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C5 = CLBLM_L_X8Y150_SLICE_X11Y150_DO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_C6 = CLBLM_L_X8Y156_SLICE_X11Y156_CO6;
  assign LIOB33_X0Y129_IOB_X0Y129_O = CLBLL_L_X4Y151_SLICE_X5Y151_CQ;
  assign LIOB33_X0Y129_IOB_X0Y130_O = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D1 = CLBLM_L_X10Y148_SLICE_X13Y148_AQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D2 = CLBLM_L_X10Y150_SLICE_X13Y150_BQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D3 = CLBLM_R_X11Y152_SLICE_X15Y152_DQ;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D4 = CLBLM_L_X8Y148_SLICE_X11Y148_CO5;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D5 = CLBLM_L_X8Y150_SLICE_X10Y150_CO5;
  assign CLBLM_L_X8Y150_SLICE_X11Y150_D6 = CLBLM_L_X8Y149_SLICE_X11Y149_DO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A1 = CLBLM_L_X8Y148_SLICE_X11Y148_CO5;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A2 = CLBLM_R_X11Y152_SLICE_X15Y152_DQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A4 = CLBLM_L_X8Y149_SLICE_X10Y149_CO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A5 = CLBLM_L_X8Y150_SLICE_X10Y150_CO5;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_A6 = CLBLM_R_X7Y156_SLICE_X9Y156_CQ;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_D1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_AX = CLBLM_L_X8Y150_SLICE_X10Y150_CO6;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B2 = CLBLM_L_X8Y150_SLICE_X10Y150_BQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B4 = CLBLM_L_X8Y151_SLICE_X10Y151_BQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B5 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_B6 = CLBLM_R_X7Y151_SLICE_X9Y151_CQ;
  assign LIOI3_X0Y161_OLOGIC_X0Y162_T1 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C2 = CLBLM_L_X10Y151_SLICE_X13Y151_CQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C4 = CLBLM_L_X8Y148_SLICE_X10Y148_BQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C5 = CLBLM_L_X8Y149_SLICE_X10Y149_AQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_C6 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_D1 = CLBLL_L_X2Y139_SLICE_X0Y139_AO5;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_D1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOI3_X0Y101_OLOGIC_X0Y102_T1 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D1 = CLBLM_L_X10Y148_SLICE_X12Y148_AQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D2 = CLBLM_R_X5Y151_SLICE_X6Y151_CQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D3 = 1'b1;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D4 = CLBLM_L_X8Y147_SLICE_X10Y147_CQ;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y150_SLICE_X10Y150_D6 = CLBLM_L_X10Y150_SLICE_X12Y150_BO5;
  assign LIOI3_X0Y161_OLOGIC_X0Y161_T1 = 1'b1;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_D1 = CLBLL_L_X2Y139_SLICE_X0Y139_AO6;
  assign LIOI3_X0Y101_OLOGIC_X0Y101_T1 = 1'b1;
  assign CLBLL_L_X4Y157_SLICE_X4Y157_A1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y157_SLICE_X4Y157_A2 = 1'b1;
  assign CLBLL_L_X4Y157_SLICE_X4Y157_A3 = 1'b1;
  assign CLBLL_L_X4Y157_SLICE_X4Y157_A4 = 1'b1;
  assign CLBLL_L_X4Y157_SLICE_X4Y157_A5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y157_SLICE_X4Y157_A6 = 1'b1;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_A1 = CLBLM_R_X7Y153_SLICE_X9Y153_CO6;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_A2 = CLBLM_R_X11Y155_SLICE_X15Y155_AQ;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_A3 = CLBLM_R_X11Y154_SLICE_X15Y154_AQ;
  assign CLBLL_L_X4Y157_SLICE_X4Y157_B1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y157_SLICE_X4Y157_B2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y157_SLICE_X4Y157_B3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y157_SLICE_X4Y157_B4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y157_SLICE_X4Y157_B5 = CLBLL_L_X4Y157_SLICE_X4Y157_CO5;
  assign CLBLL_L_X4Y157_SLICE_X4Y157_B6 = 1'b1;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_B1 = CLBLM_L_X12Y154_SLICE_X16Y154_DO6;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_B2 = CLBLM_R_X11Y154_SLICE_X15Y154_BQ;
  assign CLBLL_L_X4Y157_SLICE_X4Y157_C1 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLL_L_X4Y157_SLICE_X4Y157_C2 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y157_SLICE_X4Y157_C3 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X4Y157_SLICE_X4Y157_C4 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLL_L_X4Y157_SLICE_X4Y157_C5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X4Y157_SLICE_X4Y157_C6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A3 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A4 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A5 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B1 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B2 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B3 = 1'b1;
  assign CLBLL_L_X4Y157_SLICE_X4Y157_D1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y157_SLICE_X4Y157_D2 = CLBLM_R_X3Y158_SLICE_X2Y158_AO6;
  assign CLBLL_L_X4Y157_SLICE_X4Y157_D3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y157_SLICE_X4Y157_D4 = CLBLM_L_X8Y152_SLICE_X10Y152_CQ;
  assign CLBLL_L_X4Y157_SLICE_X4Y157_D5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y157_SLICE_X4Y157_D6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B4 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B5 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_B6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C1 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C2 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C3 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C4 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C5 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_C6 = 1'b1;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_A2 = CLBLM_R_X11Y160_SLICE_X14Y160_AQ;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D1 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D2 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D3 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D4 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D5 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_D6 = 1'b1;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_A5 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_B1 = CLBLM_R_X13Y153_SLICE_X19Y153_CQ;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_B2 = CLBLM_L_X10Y149_SLICE_X12Y149_C5Q;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A1 = CLBLM_R_X7Y157_SLICE_X8Y157_CQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y157_SLICE_X5Y157_A1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X4Y157_SLICE_X5Y157_A2 = 1'b1;
  assign CLBLL_L_X4Y157_SLICE_X5Y157_A3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X4Y157_SLICE_X5Y157_A4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y157_SLICE_X5Y157_A5 = 1'b1;
  assign CLBLL_L_X4Y157_SLICE_X5Y157_A6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A3 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A4 = CLBLM_R_X7Y144_SLICE_X8Y144_BO6;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A5 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLL_L_X4Y157_SLICE_X5Y157_B1 = CLBLL_L_X4Y157_SLICE_X4Y157_AO5;
  assign CLBLL_L_X4Y157_SLICE_X5Y157_B2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X4Y157_SLICE_X5Y157_B3 = CLBLL_L_X4Y157_SLICE_X4Y157_CO5;
  assign CLBLL_L_X4Y157_SLICE_X5Y157_B4 = CLBLM_R_X5Y157_SLICE_X6Y157_AQ;
  assign CLBLL_L_X4Y157_SLICE_X5Y157_B5 = CLBLM_R_X5Y157_SLICE_X7Y157_AQ;
  assign CLBLL_L_X4Y157_SLICE_X5Y157_B6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B1 = CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B2 = 1'b1;
  assign CLBLL_L_X4Y157_SLICE_X5Y157_C1 = CLBLL_L_X4Y157_SLICE_X4Y157_CO6;
  assign CLBLL_L_X4Y157_SLICE_X5Y157_C2 = CLBLM_R_X7Y156_SLICE_X9Y156_CQ;
  assign CLBLL_L_X4Y157_SLICE_X5Y157_C3 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X4Y157_SLICE_X5Y157_C4 = CLBLM_R_X3Y156_SLICE_X3Y156_AO5;
  assign CLBLL_L_X4Y157_SLICE_X5Y157_C5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y157_SLICE_X5Y157_C6 = CLBLM_L_X8Y156_SLICE_X11Y156_B5Q;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C1 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C2 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C3 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C4 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C5 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_C6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y157_SLICE_X5Y157_D1 = 1'b1;
  assign CLBLL_L_X4Y157_SLICE_X5Y157_D2 = 1'b1;
  assign CLBLL_L_X4Y157_SLICE_X5Y157_D3 = 1'b1;
  assign CLBLL_L_X4Y157_SLICE_X5Y157_D4 = 1'b1;
  assign CLBLL_L_X4Y157_SLICE_X5Y157_D5 = 1'b1;
  assign CLBLL_L_X4Y157_SLICE_X5Y157_D6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D1 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D2 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D3 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D4 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D5 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_D6 = 1'b1;
  assign RIOI3_X105Y145_ILOGIC_X1Y146_D = RIOB33_X105Y145_IOB_X1Y146_I;
  assign RIOI3_X105Y145_ILOGIC_X1Y145_D = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y64_D = LIOB33_X0Y63_IOB_X0Y64_I;
  assign LIOI3_TBYTETERM_X0Y63_ILOGIC_X0Y63_D = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A2 = CLBLM_R_X7Y152_SLICE_X9Y152_BQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A4 = CLBLM_L_X8Y151_SLICE_X11Y151_BO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A5 = CLBLM_R_X13Y150_SLICE_X19Y150_AQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_A6 = 1'b1;
  assign CLBLM_R_X13Y158_SLICE_X19Y158_C4 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B1 = CLBLM_L_X8Y152_SLICE_X11Y152_BO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B2 = CLBLM_L_X8Y150_SLICE_X10Y150_BQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B3 = CLBLM_R_X5Y150_SLICE_X7Y150_AQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B5 = CLBLM_L_X8Y152_SLICE_X10Y152_BQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_B6 = CLBLM_R_X7Y151_SLICE_X8Y151_DQ;
  assign CLBLM_R_X13Y158_SLICE_X19Y158_C5 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_T1 = 1'b1;
  assign CLBLM_R_X13Y158_SLICE_X19Y158_C6 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C1 = CLBLM_R_X7Y151_SLICE_X8Y151_CQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C2 = CLBLM_L_X10Y151_SLICE_X13Y151_BQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C4 = CLBLM_L_X8Y147_SLICE_X10Y147_CQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C5 = CLBLM_L_X8Y151_SLICE_X11Y151_DO6;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_C6 = CLBLM_L_X8Y151_SLICE_X10Y151_BQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D1 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D2 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D3 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D4 = CLBLM_L_X8Y152_SLICE_X10Y152_BQ;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D5 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X11Y151_D6 = CLBLM_L_X8Y150_SLICE_X10Y150_BQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A1 = CLBLM_L_X8Y151_SLICE_X11Y151_CO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A2 = CLBLM_L_X12Y154_SLICE_X17Y154_BQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A3 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A5 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B2 = CLBLM_L_X8Y151_SLICE_X10Y151_BQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B3 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B5 = CLBLM_L_X8Y151_SLICE_X11Y151_AQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_B6 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C1 = CLBLM_R_X7Y153_SLICE_X8Y153_BQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C2 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C4 = CLBLM_L_X10Y149_SLICE_X13Y149_CO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C5 = CLBLM_L_X8Y151_SLICE_X10Y151_DO6;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_T1 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D1 = CLBLM_L_X10Y157_SLICE_X12Y157_AQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D2 = CLBLM_L_X8Y151_SLICE_X10Y151_CQ;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D3 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D4 = CLBLM_R_X7Y152_SLICE_X8Y152_A5Q;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D5 = 1'b1;
  assign CLBLM_L_X8Y151_SLICE_X10Y151_D6 = CLBLM_L_X10Y150_SLICE_X12Y150_CQ;
  assign CLBLM_R_X13Y158_SLICE_X19Y158_D5 = 1'b1;
  assign CLBLM_R_X13Y158_SLICE_X19Y158_D6 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X4Y158_A1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLL_L_X4Y158_SLICE_X4Y158_A2 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLL_L_X4Y158_SLICE_X4Y158_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X4Y158_SLICE_X4Y158_A4 = CLBLL_L_X4Y157_SLICE_X4Y157_AO6;
  assign CLBLL_L_X4Y158_SLICE_X4Y158_A5 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X4Y158_A6 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X11Y155_SLICE_X15Y155_A1 = CLBLM_R_X11Y158_SLICE_X15Y158_BO6;
  assign CLBLM_R_X11Y155_SLICE_X15Y155_A2 = CLBLM_R_X5Y150_SLICE_X6Y150_DQ;
  assign CLBLM_R_X11Y155_SLICE_X15Y155_A3 = CLBLM_R_X11Y155_SLICE_X15Y155_AQ;
  assign CLBLL_L_X4Y158_SLICE_X4Y158_B1 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X4Y158_B2 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X4Y158_B3 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X4Y158_B4 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X4Y158_B5 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X4Y158_B6 = 1'b1;
  assign CLBLM_R_X11Y155_SLICE_X15Y155_A4 = 1'b1;
  assign CLBLM_R_X11Y155_SLICE_X15Y155_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y155_SLICE_X15Y155_A6 = CLBLM_L_X12Y155_SLICE_X16Y155_BO6;
  assign CLBLL_L_X4Y158_SLICE_X4Y158_C1 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X4Y158_C2 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X4Y158_C3 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X4Y158_C4 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X4Y158_C5 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X4Y158_C6 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A1 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A2 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A3 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A4 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A5 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_A6 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X4Y158_D1 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X4Y158_D2 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X4Y158_D3 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X4Y158_D4 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X4Y158_D5 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X4Y158_D6 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B1 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B2 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B3 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B4 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B5 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_B6 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C1 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C2 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C3 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C4 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C5 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_C6 = 1'b1;
  assign CLBLM_R_X11Y155_SLICE_X14Y155_A1 = CLBLM_R_X7Y153_SLICE_X9Y153_CO6;
  assign CLBLM_R_X11Y155_SLICE_X14Y155_A2 = CLBLM_R_X11Y154_SLICE_X14Y154_CQ;
  assign CLBLM_R_X11Y155_SLICE_X14Y155_A3 = CLBLM_R_X11Y155_SLICE_X14Y155_AQ;
  assign CLBLM_R_X11Y155_SLICE_X14Y155_A4 = CLBLM_R_X11Y152_SLICE_X15Y152_BQ;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D1 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D2 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D3 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D4 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D5 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X9Y145_D6 = 1'b1;
  assign CLBLM_R_X11Y155_SLICE_X14Y155_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y155_SLICE_X14Y155_A6 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X5Y158_A1 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X5Y158_A2 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X5Y158_A3 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X5Y158_A4 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X5Y158_A5 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X5Y158_A6 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A1 = CLBLM_R_X5Y146_SLICE_X6Y146_A5Q;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A2 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLL_L_X4Y158_SLICE_X5Y158_AX = CLBLM_L_X12Y159_SLICE_X16Y159_CO5;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A3 = CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  assign CLBLL_L_X4Y158_SLICE_X5Y158_B1 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X5Y158_B2 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X5Y158_B3 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X5Y158_B4 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X5Y158_B5 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X5Y158_B6 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A6 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLL_L_X4Y158_SLICE_X5Y158_C1 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X5Y158_C2 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X5Y158_C3 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X5Y158_C4 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X5Y158_C5 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X5Y158_C6 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C2 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C3 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X5Y158_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C4 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C5 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C6 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y158_SLICE_X5Y158_D1 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X5Y158_D2 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X5Y158_D3 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X5Y158_D4 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X5Y158_D5 = 1'b1;
  assign CLBLL_L_X4Y158_SLICE_X5Y158_D6 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D1 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D2 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D3 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D4 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D5 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_D6 = 1'b1;
  assign CLBLM_R_X13Y158_SLICE_X18Y158_C1 = CLBLM_R_X11Y157_SLICE_X14Y157_CQ;
  assign CLBLM_R_X11Y160_SLICE_X15Y160_D2 = 1'b1;
  assign CLBLM_R_X13Y158_SLICE_X18Y158_C2 = CLBLM_R_X13Y158_SLICE_X18Y158_AQ;
  assign CLBLM_R_X11Y160_SLICE_X15Y160_D3 = 1'b1;
  assign CLBLM_R_X13Y158_SLICE_X18Y158_C3 = CLBLM_R_X13Y159_SLICE_X18Y159_BO6;
  assign CLBLM_R_X11Y160_SLICE_X15Y160_D4 = 1'b1;
  assign CLBLM_R_X13Y158_SLICE_X18Y158_C4 = CLBLM_R_X13Y159_SLICE_X18Y159_AO6;
  assign CLBLM_R_X11Y160_SLICE_X15Y160_D5 = 1'b1;
  assign CLBLM_R_X13Y158_SLICE_X18Y158_C5 = CLBLM_R_X11Y158_SLICE_X15Y158_DO6;
  assign CLBLM_R_X11Y160_SLICE_X15Y160_D6 = 1'b1;
  assign CLBLM_R_X13Y158_SLICE_X18Y158_C6 = CLBLM_L_X12Y158_SLICE_X16Y158_BO5;
  assign CLBLM_R_X13Y158_SLICE_X18Y158_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_A1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_A2 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_A3 = CLBLM_L_X8Y150_SLICE_X11Y150_AQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_A4 = CLBLM_R_X5Y151_SLICE_X6Y151_CQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_A5 = CLBLM_L_X8Y152_SLICE_X10Y152_AQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_A6 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_B1 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_B2 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_B3 = CLBLM_R_X7Y151_SLICE_X8Y151_CQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_B4 = CLBLM_L_X8Y147_SLICE_X10Y147_CQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_B5 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_B6 = 1'b1;
  assign CLBLM_R_X13Y158_SLICE_X18Y158_D1 = CLBLM_R_X11Y157_SLICE_X15Y157_BQ;
  assign CLBLM_R_X13Y158_SLICE_X18Y158_D2 = CLBLM_R_X13Y158_SLICE_X19Y158_AO6;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_C1 = CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_C2 = CLBLL_L_X4Y153_SLICE_X4Y153_BO6;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_C4 = CLBLM_L_X8Y152_SLICE_X11Y152_AO5;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_C5 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_C6 = CLBLM_L_X10Y149_SLICE_X13Y149_BO5;
  assign CLBLM_R_X13Y158_SLICE_X18Y158_D3 = CLBLM_R_X13Y158_SLICE_X19Y158_BO6;
  assign CLBLM_R_X13Y158_SLICE_X18Y158_D4 = CLBLM_R_X11Y158_SLICE_X14Y158_BQ;
  assign CLBLM_R_X13Y158_SLICE_X18Y158_D5 = CLBLM_R_X11Y158_SLICE_X15Y158_DO6;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_D1 = CLBLM_L_X8Y147_SLICE_X10Y147_CQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_D2 = CLBLM_L_X10Y151_SLICE_X12Y151_CQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_D3 = CLBLM_L_X8Y152_SLICE_X10Y152_BQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_D4 = CLBLM_L_X8Y155_SLICE_X11Y155_DO6;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_D5 = CLBLM_R_X7Y151_SLICE_X8Y151_CQ;
  assign CLBLM_L_X8Y152_SLICE_X11Y152_D6 = CLBLM_L_X8Y150_SLICE_X10Y150_BQ;
  assign CLBLM_R_X13Y158_SLICE_X18Y158_D6 = CLBLM_L_X12Y158_SLICE_X16Y158_BO5;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_A1 = CLBLM_L_X8Y152_SLICE_X10Y152_DO6;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_A2 = CLBLL_L_X4Y146_SLICE_X5Y146_AQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_A3 = CLBLM_L_X8Y152_SLICE_X10Y152_AQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_A6 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_T1 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_B2 = CLBLM_L_X8Y152_SLICE_X10Y152_BQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_B3 = CLBLM_L_X8Y153_SLICE_X10Y153_AQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_B5 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_B6 = CLBLM_R_X7Y151_SLICE_X9Y151_CQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_C1 = CLBLM_L_X10Y148_SLICE_X13Y148_BQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_C2 = CLBLM_L_X8Y152_SLICE_X10Y152_CQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_C3 = CLBLM_R_X13Y153_SLICE_X19Y153_AQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_C4 = CLBLM_L_X10Y150_SLICE_X12Y150_A5Q;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_C5 = CLBLM_L_X12Y155_SLICE_X16Y155_CO6;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y160_SLICE_X14Y160_B6 = 1'b1;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_D1 = CLBLM_R_X5Y151_SLICE_X7Y151_CQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_D2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_D3 = CLBLM_L_X8Y152_SLICE_X11Y152_BO5;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_D4 = CLBLM_L_X8Y152_SLICE_X10Y152_BQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_D5 = CLBLM_R_X11Y151_SLICE_X15Y151_AQ;
  assign CLBLM_L_X8Y152_SLICE_X10Y152_D6 = CLBLM_L_X8Y150_SLICE_X10Y150_BQ;
  assign CLBLM_R_X11Y160_SLICE_X14Y160_C4 = 1'b1;
  assign CLBLM_R_X11Y160_SLICE_X14Y160_C5 = 1'b1;
  assign CLBLM_R_X11Y156_SLICE_X15Y156_A1 = CLBLM_L_X10Y159_SLICE_X12Y159_DO6;
  assign CLBLM_R_X11Y156_SLICE_X15Y156_A2 = CLBLM_R_X11Y157_SLICE_X15Y157_CO6;
  assign CLBLM_R_X11Y156_SLICE_X15Y156_A3 = CLBLM_R_X11Y156_SLICE_X15Y156_AQ;
  assign CLBLM_R_X11Y156_SLICE_X15Y156_A4 = CLBLM_L_X10Y159_SLICE_X12Y159_CO6;
  assign CLBLM_R_X11Y156_SLICE_X15Y156_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y156_SLICE_X15Y156_A6 = CLBLL_L_X4Y149_SLICE_X5Y149_AQ;
  assign CLBLM_R_X11Y160_SLICE_X14Y160_C6 = 1'b1;
  assign CLBLM_R_X11Y156_SLICE_X15Y156_B1 = 1'b1;
  assign CLBLM_R_X11Y156_SLICE_X15Y156_B2 = CLBLM_R_X11Y156_SLICE_X15Y156_BQ;
  assign CLBLM_R_X11Y156_SLICE_X15Y156_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y156_SLICE_X15Y156_B4 = CLBLM_R_X11Y159_SLICE_X15Y159_BQ;
  assign CLBLM_R_X11Y156_SLICE_X15Y156_B5 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_R_X11Y156_SLICE_X15Y156_B6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign LIOB33_X0Y165_IOB_X0Y165_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign LIOB33_X0Y165_IOB_X0Y166_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A1 = CLBLM_R_X5Y150_SLICE_X7Y150_A5Q;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A2 = CLBLM_R_X7Y146_SLICE_X8Y146_DO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A3 = CLBLM_R_X7Y146_SLICE_X9Y146_AQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A5 = CLBLM_L_X10Y146_SLICE_X12Y146_BQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_A6 = 1'b1;
  assign CLBLM_R_X11Y156_SLICE_X15Y156_C1 = CLBLM_R_X11Y158_SLICE_X15Y158_DO6;
  assign CLBLM_R_X11Y156_SLICE_X15Y156_C2 = CLBLM_R_X11Y156_SLICE_X14Y156_CO6;
  assign CLBLM_R_X11Y156_SLICE_X15Y156_C3 = CLBLM_R_X11Y150_SLICE_X15Y150_BO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B1 = CLBLM_R_X3Y156_SLICE_X2Y156_DO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B2 = CLBLM_R_X3Y155_SLICE_X2Y155_BO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B3 = CLBLL_L_X4Y154_SLICE_X5Y154_CO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B4 = CLBLL_L_X4Y153_SLICE_X4Y153_BO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B5 = CLBLL_L_X4Y154_SLICE_X5Y154_BO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_B6 = CLBLM_R_X5Y155_SLICE_X6Y155_DO6;
  assign CLBLM_R_X11Y156_SLICE_X15Y156_D1 = CLBLM_L_X10Y158_SLICE_X13Y158_AQ;
  assign CLBLM_R_X11Y156_SLICE_X15Y156_D2 = CLBLM_R_X11Y157_SLICE_X14Y157_CQ;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C1 = CLBLM_R_X7Y148_SLICE_X9Y148_CO5;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C2 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C3 = CLBLM_L_X8Y153_SLICE_X11Y153_C5Q;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C4 = CLBLM_R_X7Y147_SLICE_X8Y147_BO5;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_C6 = CLBLM_R_X7Y146_SLICE_X9Y146_BO6;
  assign CLBLM_R_X11Y156_SLICE_X15Y156_D3 = 1'b1;
  assign CLBLM_R_X11Y156_SLICE_X15Y156_D4 = CLBLM_R_X11Y159_SLICE_X15Y159_DO5;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y156_SLICE_X14Y156_A1 = CLBLM_R_X11Y159_SLICE_X15Y159_DO5;
  assign CLBLM_R_X11Y156_SLICE_X14Y156_A2 = CLBLM_R_X11Y158_SLICE_X15Y158_BO6;
  assign CLBLM_R_X11Y156_SLICE_X14Y156_A3 = CLBLM_R_X11Y156_SLICE_X14Y156_AQ;
  assign CLBLM_R_X11Y156_SLICE_X14Y156_A4 = CLBLM_R_X3Y150_SLICE_X3Y150_CQ;
  assign CLBLM_R_X11Y156_SLICE_X14Y156_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D2 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D3 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D4 = CLBLM_R_X7Y146_SLICE_X9Y146_CO6;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D5 = CLBLM_R_X5Y150_SLICE_X7Y150_A5Q;
  assign CLBLM_R_X7Y146_SLICE_X9Y146_D6 = CLBLM_R_X7Y147_SLICE_X9Y147_A5Q;
  assign CLBLM_R_X11Y156_SLICE_X14Y156_A6 = CLBLM_L_X12Y157_SLICE_X16Y157_BQ;
  assign CLBLM_R_X11Y156_SLICE_X14Y156_B1 = CLBLM_L_X10Y157_SLICE_X13Y157_CO6;
  assign CLBLM_R_X11Y156_SLICE_X14Y156_B2 = CLBLM_L_X10Y159_SLICE_X12Y159_CO6;
  assign CLBLM_R_X11Y156_SLICE_X14Y156_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y156_SLICE_X14Y156_B4 = CLBLM_L_X10Y159_SLICE_X12Y159_DO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A3 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A4 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A5 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_A6 = CLBLM_R_X5Y146_SLICE_X6Y146_A5Q;
  assign CLBLM_R_X11Y156_SLICE_X14Y156_C1 = CLBLM_R_X11Y156_SLICE_X15Y156_AQ;
  assign CLBLM_R_X11Y156_SLICE_X14Y156_C2 = CLBLM_L_X8Y156_SLICE_X11Y156_DO6;
  assign CLBLM_R_X11Y156_SLICE_X14Y156_C3 = CLBLM_L_X10Y157_SLICE_X13Y157_AO5;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B1 = CLBLM_R_X5Y150_SLICE_X7Y150_A5Q;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B2 = CLBLM_R_X5Y147_SLICE_X7Y147_C5Q;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B3 = CLBLM_R_X7Y147_SLICE_X8Y147_DO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B4 = CLBLL_L_X4Y146_SLICE_X5Y146_AQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_B6 = 1'b1;
  assign CLBLM_R_X11Y156_SLICE_X14Y156_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y156_SLICE_X14Y156_D1 = 1'b1;
  assign CLBLM_R_X11Y156_SLICE_X14Y156_D2 = CLBLM_R_X11Y155_SLICE_X14Y155_CQ;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C1 = CLBLM_R_X7Y148_SLICE_X9Y148_CO5;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C2 = CLBLM_R_X7Y147_SLICE_X8Y147_DO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C3 = CLBLM_R_X7Y146_SLICE_X9Y146_BO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C4 = CLBLM_R_X5Y147_SLICE_X7Y147_C5Q;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C5 = CLBLM_R_X7Y146_SLICE_X8Y146_BO5;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_C6 = CLBLL_L_X4Y146_SLICE_X5Y146_AQ;
  assign CLBLM_R_X11Y156_SLICE_X14Y156_D3 = CLBLM_L_X10Y157_SLICE_X12Y157_DO6;
  assign CLBLM_R_X11Y156_SLICE_X14Y156_D4 = CLBLM_L_X10Y159_SLICE_X12Y159_DO6;
  assign CLBLM_R_X11Y156_SLICE_X14Y156_D5 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y156_SLICE_X14Y156_D6 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_T1 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D1 = CLBLM_R_X7Y148_SLICE_X9Y148_CO5;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D2 = 1'b1;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D3 = CLBLM_R_X7Y146_SLICE_X9Y146_BO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D4 = CLBLM_R_X7Y147_SLICE_X8Y147_CO6;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D5 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_R_X7Y146_SLICE_X8Y146_D6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_T1 = 1'b1;
  assign CLBLM_L_X10Y163_SLICE_X13Y163_A1 = 1'b1;
  assign CLBLM_L_X10Y163_SLICE_X13Y163_A2 = 1'b1;
  assign CLBLM_L_X10Y163_SLICE_X13Y163_A3 = 1'b1;
  assign CLBLM_L_X10Y163_SLICE_X13Y163_A4 = 1'b1;
  assign CLBLM_L_X10Y163_SLICE_X13Y163_A5 = 1'b1;
  assign CLBLM_L_X10Y163_SLICE_X13Y163_A6 = CLBLM_L_X10Y155_SLICE_X13Y155_A5Q;
  assign CLBLM_L_X10Y163_SLICE_X13Y163_B1 = 1'b1;
  assign CLBLM_L_X10Y163_SLICE_X13Y163_B2 = 1'b1;
  assign CLBLM_L_X10Y163_SLICE_X13Y163_B3 = 1'b1;
  assign CLBLM_L_X10Y163_SLICE_X13Y163_B4 = 1'b1;
  assign CLBLM_L_X10Y163_SLICE_X13Y163_B5 = 1'b1;
  assign CLBLM_L_X10Y163_SLICE_X13Y163_B6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_D1 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_A1 = CLBLM_L_X10Y153_SLICE_X13Y153_DQ;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_A3 = CLBLM_L_X8Y153_SLICE_X11Y153_AQ;
  assign CLBLM_L_X10Y163_SLICE_X13Y163_C4 = 1'b1;
  assign CLBLM_L_X10Y163_SLICE_X13Y163_C5 = 1'b1;
  assign CLBLM_L_X10Y163_SLICE_X13Y163_C6 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_A4 = CLBLL_L_X4Y148_SLICE_X5Y148_DQ;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_A5 = CLBLM_R_X13Y150_SLICE_X18Y150_BQ;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_A6 = CLBLM_R_X7Y153_SLICE_X9Y153_CO6;
  assign CLBLM_L_X10Y163_SLICE_X13Y163_C1 = 1'b1;
  assign CLBLM_L_X10Y163_SLICE_X13Y163_C2 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_B1 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_B3 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_B4 = CLBLM_R_X11Y159_SLICE_X15Y159_CO6;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_B5 = CLBLM_L_X8Y153_SLICE_X10Y153_AQ;
  assign CLBLM_L_X10Y163_SLICE_X13Y163_D3 = 1'b1;
  assign CLBLM_L_X10Y163_SLICE_X13Y163_D4 = 1'b1;
  assign CLBLM_L_X10Y163_SLICE_X13Y163_D5 = 1'b1;
  assign CLBLM_L_X10Y163_SLICE_X13Y163_D6 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_B6 = CLBLM_L_X10Y153_SLICE_X13Y153_DQ;
  assign CLBLM_L_X10Y163_SLICE_X13Y163_D1 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_C2 = CLBLM_L_X10Y154_SLICE_X12Y154_DQ;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_C3 = CLBLM_L_X8Y153_SLICE_X11Y153_DQ;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_C5 = CLBLM_R_X7Y148_SLICE_X8Y148_A5Q;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_C6 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y163_SLICE_X12Y163_A1 = 1'b1;
  assign CLBLM_L_X10Y163_SLICE_X12Y163_A2 = 1'b1;
  assign CLBLM_L_X10Y163_SLICE_X12Y163_A3 = 1'b1;
  assign CLBLM_L_X10Y163_SLICE_X12Y163_A4 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_D1 = CLBLM_L_X10Y152_SLICE_X13Y152_BO5;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_D2 = CLBLM_L_X8Y153_SLICE_X10Y153_A5Q;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_D3 = CLBLM_R_X5Y152_SLICE_X6Y152_AQ;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_D5 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X11Y153_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y163_SLICE_X12Y163_B1 = 1'b1;
  assign CLBLM_L_X10Y163_SLICE_X12Y163_B2 = 1'b1;
  assign CLBLM_L_X10Y163_SLICE_X12Y163_B3 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_A1 = CLBLM_L_X8Y154_SLICE_X10Y154_CQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_A2 = CLBLM_L_X8Y157_SLICE_X10Y157_DQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_A3 = CLBLM_L_X10Y151_SLICE_X13Y151_BQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_A4 = CLBLM_R_X11Y159_SLICE_X15Y159_CO6;
  assign CLBLM_L_X10Y163_SLICE_X12Y163_C4 = 1'b1;
  assign CLBLM_L_X10Y163_SLICE_X12Y163_C5 = 1'b1;
  assign CLBLM_L_X10Y163_SLICE_X12Y163_C6 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_A6 = 1'b1;
  assign CLBLM_L_X10Y163_SLICE_X12Y163_C1 = 1'b1;
  assign CLBLM_L_X10Y163_SLICE_X12Y163_C2 = 1'b1;
  assign CLBLM_L_X10Y163_SLICE_X12Y163_C3 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_B1 = CLBLM_L_X8Y152_SLICE_X11Y152_BO5;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_B2 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_B3 = CLBLM_L_X8Y152_SLICE_X10Y152_BQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_B4 = CLBLM_L_X8Y158_SLICE_X10Y158_BQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_B5 = CLBLM_L_X8Y150_SLICE_X10Y150_BQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_B6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y163_SLICE_X12Y163_D1 = 1'b1;
  assign CLBLM_L_X10Y163_SLICE_X12Y163_D2 = 1'b1;
  assign CLBLM_L_X10Y163_SLICE_X12Y163_D3 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_C1 = CLBLM_L_X8Y152_SLICE_X10Y152_BQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_C2 = CLBLM_L_X8Y150_SLICE_X10Y150_BQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_C3 = CLBLM_R_X5Y152_SLICE_X6Y152_BQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_C4 = CLBLM_R_X7Y157_SLICE_X9Y157_DQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_C5 = CLBLM_L_X8Y152_SLICE_X11Y152_BO5;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_C6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y163_SLICE_X12Y163_D5 = 1'b1;
  assign CLBLM_L_X10Y163_SLICE_X12Y163_D6 = 1'b1;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_D1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_D2 = CLBLM_L_X10Y153_SLICE_X12Y153_CO6;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_D3 = CLBLM_R_X7Y153_SLICE_X9Y153_CO6;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_D4 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_D5 = CLBLM_L_X8Y155_SLICE_X11Y155_DO6;
  assign CLBLM_L_X8Y153_SLICE_X10Y153_D6 = CLBLM_R_X5Y151_SLICE_X7Y151_BQ;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C4 = 1'b1;
  assign RIOI3_X105Y147_ILOGIC_X1Y148_D = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C5 = 1'b1;
  assign RIOI3_X105Y147_ILOGIC_X1Y147_D = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_C6 = CLBLM_L_X8Y147_SLICE_X11Y147_BQ;
  assign LIOB33_X0Y167_IOB_X0Y168_O = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOB33_X0Y167_IOB_X0Y167_O = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_A1 = CLBLM_R_X11Y158_SLICE_X15Y158_BO5;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_A2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_A3 = CLBLM_R_X11Y157_SLICE_X15Y157_AQ;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_A4 = CLBLM_L_X10Y155_SLICE_X13Y155_BQ;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_A6 = CLBLM_L_X12Y157_SLICE_X16Y157_DO6;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_B1 = CLBLM_L_X8Y149_SLICE_X11Y149_CQ;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_B2 = CLBLM_R_X11Y159_SLICE_X15Y159_CO5;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_B3 = CLBLM_L_X12Y156_SLICE_X16Y156_DO6;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_B4 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_B6 = CLBLM_R_X11Y158_SLICE_X14Y158_DO5;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A2 = CLBLM_R_X3Y151_SLICE_X2Y151_AQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A3 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A4 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A5 = CLBLM_L_X10Y149_SLICE_X12Y149_BQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_A6 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_C1 = CLBLM_L_X8Y156_SLICE_X11Y156_DO6;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_C2 = CLBLM_L_X12Y157_SLICE_X16Y157_CQ;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_C3 = CLBLM_L_X10Y157_SLICE_X13Y157_AO5;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B2 = CLBLM_R_X7Y147_SLICE_X9Y147_BQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B4 = CLBLM_R_X7Y147_SLICE_X9Y147_DO5;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B5 = CLBLM_R_X7Y147_SLICE_X8Y147_AQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_B6 = CLBLM_L_X10Y154_SLICE_X13Y154_CQ;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_D1 = CLBLM_L_X10Y159_SLICE_X12Y159_DO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C1 = CLBLM_R_X7Y151_SLICE_X9Y151_AQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C2 = CLBLM_R_X7Y147_SLICE_X9Y147_CQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C4 = CLBLM_L_X10Y154_SLICE_X13Y154_CQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C5 = CLBLM_R_X7Y147_SLICE_X9Y147_DO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D5 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_D4 = CLBLM_L_X8Y156_SLICE_X11Y156_DO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y150_SLICE_X15Y150_D6 = CLBLM_R_X11Y155_SLICE_X14Y155_BQ;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_A1 = CLBLM_L_X12Y157_SLICE_X17Y157_DO6;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_A2 = CLBLM_R_X11Y157_SLICE_X14Y157_AQ;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_A4 = CLBLM_R_X11Y159_SLICE_X15Y159_CO5;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D1 = CLBLM_L_X8Y147_SLICE_X10Y147_BQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D2 = CLBLM_R_X7Y147_SLICE_X9Y147_CQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D3 = CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D4 = CLBLM_R_X7Y147_SLICE_X9Y147_BQ;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D5 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_R_X7Y147_SLICE_X9Y147_D6 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_A5 = CLBLM_L_X8Y157_SLICE_X11Y157_BQ;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_A6 = CLBLM_R_X11Y158_SLICE_X14Y158_DO5;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_B1 = CLBLM_R_X11Y159_SLICE_X15Y159_DO5;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_B2 = CLBLL_L_X4Y152_SLICE_X5Y152_BQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A1 = CLBLM_R_X5Y149_SLICE_X6Y149_AQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A2 = 1'b1;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A3 = CLBLM_R_X7Y147_SLICE_X8Y147_AQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A5 = CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_A6 = CLBLL_L_X4Y147_SLICE_X4Y147_BO6;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_C1 = CLBLM_R_X7Y157_SLICE_X9Y157_AQ;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_C2 = CLBLM_R_X11Y157_SLICE_X14Y157_CQ;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_C3 = CLBLM_R_X11Y157_SLICE_X14Y157_BQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B1 = CLBLM_R_X5Y149_SLICE_X6Y149_AQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B2 = CLBLM_R_X5Y148_SLICE_X7Y148_A5Q;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B3 = CLBLM_R_X5Y147_SLICE_X7Y147_C5Q;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B4 = CLBLM_R_X5Y151_SLICE_X6Y151_C5Q;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B5 = CLBLL_L_X4Y146_SLICE_X5Y146_AQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_B6 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_D1 = CLBLM_L_X10Y159_SLICE_X12Y159_DO6;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_D2 = CLBLM_L_X10Y155_SLICE_X13Y155_CO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C1 = CLBLM_R_X7Y147_SLICE_X9Y147_A5Q;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C2 = CLBLM_R_X5Y149_SLICE_X6Y149_AQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C3 = CLBLM_L_X8Y153_SLICE_X11Y153_C5Q;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C4 = CLBLM_R_X5Y150_SLICE_X7Y150_A5Q;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_C6 = CLBLM_R_X7Y147_SLICE_X8Y147_BO6;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_D3 = CLBLM_R_X3Y153_SLICE_X3Y153_BO6;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_D4 = CLBLM_L_X10Y159_SLICE_X13Y159_CO6;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_D5 = CLBLM_L_X12Y157_SLICE_X17Y157_DO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_D6 = CLBLM_L_X10Y159_SLICE_X12Y159_CO6;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D1 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D2 = CLBLM_R_X7Y147_SLICE_X9Y147_A5Q;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D3 = CLBLM_R_X5Y149_SLICE_X6Y149_AQ;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D4 = CLBLM_L_X8Y153_SLICE_X11Y153_C5Q;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D5 = CLBLM_R_X5Y148_SLICE_X7Y148_A5Q;
  assign CLBLM_R_X7Y147_SLICE_X8Y147_D6 = CLBLM_R_X5Y151_SLICE_X6Y151_C5Q;
  assign LIOI3_X0Y159_OLOGIC_X0Y159_T1 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_A1 = CLBLM_R_X7Y153_SLICE_X9Y153_CO6;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_A2 = CLBLM_L_X10Y156_SLICE_X13Y156_BQ;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_A3 = CLBLM_L_X8Y154_SLICE_X11Y154_AQ;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_A4 = CLBLM_R_X7Y154_SLICE_X8Y154_CQ;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_A5 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOB33_X0Y151_IOB_X0Y152_O = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_AX = CLBLM_R_X11Y154_SLICE_X14Y154_BO6;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_B1 = CLBLM_L_X8Y155_SLICE_X10Y155_BQ;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_B2 = CLBLM_L_X8Y154_SLICE_X11Y154_BQ;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_B3 = CLBLM_R_X7Y153_SLICE_X9Y153_CO6;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_B5 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_B6 = CLBLM_L_X10Y154_SLICE_X12Y154_DQ;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_C1 = CLBLM_L_X10Y157_SLICE_X12Y157_AQ;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_C2 = CLBLM_L_X8Y154_SLICE_X11Y154_CQ;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_C4 = CLBLM_L_X8Y153_SLICE_X10Y153_CO6;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_C5 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOB33_X0Y151_IOB_X0Y151_O = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_D1 = CLBLM_R_X5Y151_SLICE_X7Y151_CQ;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_D2 = CLBLM_R_X7Y157_SLICE_X9Y157_DQ;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_D3 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_D4 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_D5 = CLBLM_R_X5Y150_SLICE_X7Y150_AQ;
  assign CLBLM_L_X8Y154_SLICE_X11Y154_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_D1 = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_A1 = CLBLM_R_X7Y156_SLICE_X9Y156_DO6;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_A2 = CLBLL_L_X4Y152_SLICE_X5Y152_CQ;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_A3 = CLBLM_L_X12Y156_SLICE_X16Y156_CO6;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_A5 = CLBLM_L_X8Y147_SLICE_X11Y147_AQ;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_A6 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_B1 = CLBLM_R_X3Y150_SLICE_X2Y150_A5Q;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_B2 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_B3 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_B5 = CLBLM_L_X10Y158_SLICE_X12Y158_BQ;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_B6 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_C1 = CLBLM_L_X8Y157_SLICE_X11Y157_AQ;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_C2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_C4 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_C5 = CLBLM_L_X8Y154_SLICE_X10Y154_B5Q;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_C6 = 1'b1;
  assign LIOB33_X0Y169_IOB_X0Y170_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_A2 = RIOB33_X105Y139_IOB_X1Y140_I;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_A3 = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_A4 = RIOB33_X105Y137_IOB_X1Y138_I;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_A5 = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_A6 = 1'b1;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_D2 = CLBLM_R_X11Y149_SLICE_X14Y149_DQ;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_D3 = CLBLM_L_X8Y154_SLICE_X10Y154_DQ;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_D4 = CLBLM_L_X10Y150_SLICE_X12Y150_A5Q;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_D5 = CLBLM_L_X12Y155_SLICE_X16Y155_CO6;
  assign CLBLM_L_X8Y154_SLICE_X10Y154_D6 = CLBLM_L_X8Y158_SLICE_X10Y158_BQ;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_A4 = CLBLM_R_X7Y158_SLICE_X8Y158_CO5;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_B1 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_B2 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_B3 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_B4 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_B5 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_B6 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_C1 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_C2 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_C3 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_C4 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_C5 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_C6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y169_T1 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_D1 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_D2 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_D3 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_D4 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_D5 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X163Y141_D6 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_A1 = 1'b1;
  assign CLBLM_R_X11Y158_SLICE_X15Y158_A1 = CLBLM_L_X12Y152_SLICE_X17Y152_AQ;
  assign CLBLM_R_X11Y158_SLICE_X15Y158_A2 = CLBLM_L_X10Y158_SLICE_X13Y158_AQ;
  assign CLBLM_R_X11Y158_SLICE_X15Y158_A3 = CLBLM_R_X11Y158_SLICE_X15Y158_AQ;
  assign CLBLM_R_X11Y158_SLICE_X15Y158_A4 = CLBLM_R_X11Y158_SLICE_X15Y158_BO6;
  assign CLBLM_R_X11Y158_SLICE_X15Y158_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y158_SLICE_X15Y158_A6 = CLBLM_R_X11Y159_SLICE_X15Y159_DO5;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_A2 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_A3 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_B2 = CLBLM_L_X8Y157_SLICE_X11Y157_BQ;
  assign CLBLM_R_X11Y158_SLICE_X15Y158_B1 = CLBLM_R_X11Y159_SLICE_X14Y159_BQ;
  assign CLBLM_R_X11Y158_SLICE_X15Y158_B2 = CLBLM_R_X11Y159_SLICE_X15Y159_AQ;
  assign CLBLM_R_X11Y158_SLICE_X15Y158_B3 = CLBLM_L_X12Y155_SLICE_X16Y155_BO5;
  assign CLBLM_R_X11Y158_SLICE_X15Y158_B4 = CLBLM_L_X12Y158_SLICE_X17Y158_AQ;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y158_SLICE_X15Y158_B5 = CLBLM_L_X12Y158_SLICE_X16Y158_AQ;
  assign CLBLM_R_X11Y158_SLICE_X15Y158_B6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A1 = CLBLM_L_X8Y148_SLICE_X10Y148_CQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A2 = CLBLM_R_X5Y152_SLICE_X6Y152_CO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A3 = CLBLM_R_X7Y148_SLICE_X9Y148_AQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A4 = CLBLM_R_X7Y151_SLICE_X8Y151_BQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_A6 = 1'b1;
  assign CLBLM_R_X11Y158_SLICE_X15Y158_C1 = CLBLM_R_X11Y157_SLICE_X15Y157_AQ;
  assign CLBLM_R_X11Y158_SLICE_X15Y158_C2 = CLBLM_R_X11Y159_SLICE_X15Y159_AQ;
  assign CLBLM_R_X11Y158_SLICE_X15Y158_C3 = CLBLM_L_X8Y157_SLICE_X10Y157_DQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B2 = CLBLM_R_X7Y148_SLICE_X9Y148_BQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B3 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B4 = CLBLM_L_X8Y146_SLICE_X10Y146_AQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B5 = CLBLM_R_X5Y147_SLICE_X7Y147_C5Q;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_B6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y158_SLICE_X15Y158_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y158_SLICE_X15Y158_D1 = CLBLM_R_X11Y157_SLICE_X15Y157_AQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C1 = CLBLL_L_X4Y153_SLICE_X4Y153_AO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C2 = CLBLM_R_X3Y156_SLICE_X2Y156_DO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C3 = CLBLL_L_X4Y154_SLICE_X5Y154_BO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C4 = CLBLL_L_X4Y154_SLICE_X4Y154_BO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C5 = CLBLM_R_X7Y148_SLICE_X9Y148_DO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_C6 = 1'b1;
  assign CLBLM_R_X11Y158_SLICE_X15Y158_D4 = CLBLM_R_X11Y159_SLICE_X14Y159_BQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y158_SLICE_X14Y158_A1 = 1'b1;
  assign CLBLM_R_X11Y158_SLICE_X14Y158_A2 = CLBLM_R_X13Y156_SLICE_X18Y156_BO6;
  assign CLBLM_R_X11Y158_SLICE_X14Y158_A3 = CLBLM_R_X11Y159_SLICE_X15Y159_CO5;
  assign CLBLM_R_X11Y158_SLICE_X14Y158_A4 = CLBLM_R_X11Y158_SLICE_X14Y158_DO5;
  assign CLBLM_R_X11Y158_SLICE_X14Y158_A5 = CLBLM_R_X7Y158_SLICE_X8Y158_AQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D1 = CLBLL_L_X4Y154_SLICE_X5Y154_CO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D2 = CLBLM_R_X5Y155_SLICE_X6Y155_DO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D3 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D4 = CLBLM_R_X3Y155_SLICE_X2Y155_BO6;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D5 = CLBLM_L_X10Y150_SLICE_X13Y150_BQ;
  assign CLBLM_R_X7Y148_SLICE_X9Y148_D6 = CLBLL_L_X4Y153_SLICE_X4Y153_BO6;
  assign CLBLM_R_X11Y158_SLICE_X14Y158_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y158_SLICE_X14Y158_B1 = CLBLM_R_X11Y159_SLICE_X15Y159_DO5;
  assign CLBLM_R_X11Y158_SLICE_X14Y158_B2 = CLBLM_R_X11Y158_SLICE_X15Y158_BO6;
  assign CLBLM_R_X11Y158_SLICE_X14Y158_B3 = CLBLM_R_X11Y156_SLICE_X14Y156_AQ;
  assign CLBLM_R_X11Y158_SLICE_X14Y158_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A2 = CLBLM_R_X7Y148_SLICE_X8Y148_BQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A3 = CLBLM_R_X7Y148_SLICE_X8Y148_AQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A5 = CLBLM_R_X5Y144_SLICE_X6Y144_AQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_A6 = CLBLM_L_X10Y159_SLICE_X12Y159_AO6;
  assign CLBLM_R_X11Y158_SLICE_X14Y158_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y158_SLICE_X14Y158_C2 = CLBLM_L_X10Y154_SLICE_X12Y154_CQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_AX = CLBLM_R_X7Y148_SLICE_X8Y148_DO6;
  assign CLBLM_R_X11Y158_SLICE_X14Y158_C3 = CLBLM_L_X12Y158_SLICE_X16Y158_AQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B2 = CLBLM_R_X7Y148_SLICE_X8Y148_BQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B4 = CLBLM_R_X7Y159_SLICE_X8Y159_BO6;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B5 = CLBLM_R_X7Y146_SLICE_X9Y146_AQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_B6 = CLBLM_R_X7Y158_SLICE_X8Y158_CO5;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_C6 = CLBLM_R_X7Y148_SLICE_X8Y148_BQ;
  assign CLBLM_R_X11Y158_SLICE_X14Y158_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y158_SLICE_X14Y158_D1 = CLBLM_R_X11Y157_SLICE_X15Y157_AQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C1 = CLBLM_L_X10Y149_SLICE_X12Y149_DO5;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C2 = CLBLM_R_X7Y148_SLICE_X8Y148_CQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C4 = CLBLL_L_X4Y148_SLICE_X5Y148_DQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C5 = CLBLM_R_X7Y151_SLICE_X9Y151_CQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_C6 = CLBLM_R_X7Y148_SLICE_X8Y148_DO5;
  assign CLBLM_R_X11Y158_SLICE_X14Y158_D2 = CLBLM_R_X11Y159_SLICE_X14Y159_BQ;
  assign CLBLM_R_X11Y158_SLICE_X14Y158_D3 = CLBLM_L_X12Y158_SLICE_X16Y158_AQ;
  assign CLBLM_R_X11Y158_SLICE_X14Y158_D4 = CLBLM_R_X11Y159_SLICE_X15Y159_AQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y158_SLICE_X14Y158_D6 = 1'b1;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D1 = CLBLM_L_X10Y149_SLICE_X12Y149_DO5;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D2 = CLBLM_L_X10Y149_SLICE_X12Y149_BQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D3 = CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D4 = CLBLM_R_X7Y148_SLICE_X8Y148_A5Q;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y148_SLICE_X8Y148_D6 = 1'b1;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_D1 = RIOB33_X105Y123_IOB_X1Y123_I;
  assign LIOI3_X0Y167_OLOGIC_X0Y168_T1 = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_D1 = CLBLL_L_X2Y140_SLICE_X0Y140_BO5;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_D1 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign LIOI3_X0Y105_OLOGIC_X0Y106_T1 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_D1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_A1 = CLBLM_R_X7Y151_SLICE_X8Y151_CQ;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_A2 = CLBLM_R_X13Y155_SLICE_X18Y155_BQ;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_A3 = CLBLM_L_X8Y155_SLICE_X11Y155_AQ;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_A5 = 1'b1;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_A6 = CLBLM_R_X7Y153_SLICE_X9Y153_CO6;
  assign LIOI3_X0Y167_OLOGIC_X0Y167_T1 = 1'b1;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_D1 = CLBLL_L_X2Y140_SLICE_X0Y140_BO6;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_B1 = CLBLM_L_X10Y153_SLICE_X13Y153_DQ;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_B3 = 1'b1;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_B4 = CLBLM_L_X12Y153_SLICE_X17Y153_DO5;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_B5 = CLBLM_R_X5Y155_SLICE_X7Y155_BQ;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_D1 = CLBLM_L_X8Y146_SLICE_X10Y146_BQ;
  assign LIOI3_X0Y105_OLOGIC_X0Y105_T1 = 1'b1;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_C1 = 1'b1;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_C3 = CLBLM_L_X8Y156_SLICE_X10Y156_CQ;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_C4 = 1'b1;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_C5 = CLBLM_R_X7Y154_SLICE_X9Y154_AQ;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_D1 = LIOB33_X0Y75_IOB_X0Y76_I;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y114_T1 = 1'b1;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign RIOI3_X105Y151_OLOGIC_X1Y151_T1 = 1'b1;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_D1 = 1'b1;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_D2 = CLBLM_L_X8Y157_SLICE_X11Y157_CQ;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_D3 = CLBLM_L_X10Y155_SLICE_X12Y155_DO6;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_D4 = CLBLM_L_X8Y156_SLICE_X11Y156_BQ;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_D5 = CLBLM_L_X8Y154_SLICE_X11Y154_DO6;
  assign CLBLM_L_X8Y155_SLICE_X11Y155_D6 = CLBLM_L_X10Y150_SLICE_X12Y150_DO6;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_D1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign LIOB33_X0Y171_IOB_X0Y172_O = CLBLM_R_X103Y141_SLICE_X163Y141_AO6;
  assign LIOB33_X0Y171_IOB_X0Y171_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_A1 = 1'b1;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_A2 = CLBLM_L_X10Y155_SLICE_X12Y155_CQ;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_A3 = CLBLM_R_X5Y152_SLICE_X6Y152_BQ;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_A4 = CLBLM_L_X8Y155_SLICE_X10Y155_AQ;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_A6 = CLBLM_R_X7Y153_SLICE_X9Y153_CO6;
  assign LIOI3_TBYTETERM_X0Y113_OLOGIC_X0Y113_T1 = 1'b1;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_B1 = CLBLM_L_X8Y149_SLICE_X10Y149_DO6;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_B2 = CLBLM_R_X5Y155_SLICE_X6Y155_AQ;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_B3 = CLBLM_L_X8Y154_SLICE_X11Y154_A5Q;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_B4 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_B6 = 1'b1;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_C1 = CLBLM_L_X10Y150_SLICE_X12Y150_A5Q;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_C2 = CLBLM_L_X8Y155_SLICE_X10Y155_CQ;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_C3 = CLBLM_L_X12Y155_SLICE_X16Y155_CO6;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_C4 = CLBLM_L_X10Y155_SLICE_X12Y155_BQ;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_C6 = CLBLM_L_X8Y155_SLICE_X10Y155_AQ;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_D1 = CLBLM_L_X8Y152_SLICE_X10Y152_CQ;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_D2 = CLBLM_L_X8Y153_SLICE_X10Y153_DO6;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_D3 = CLBLM_L_X8Y149_SLICE_X10Y149_DO6;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_D4 = CLBLL_L_X4Y156_SLICE_X4Y156_CO5;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_D5 = CLBLM_R_X7Y155_SLICE_X9Y155_CO6;
  assign CLBLM_L_X8Y155_SLICE_X10Y155_D6 = CLBLM_R_X13Y152_SLICE_X19Y152_CO6;
  assign CLBLM_R_X11Y159_SLICE_X15Y159_A1 = CLBLM_R_X11Y159_SLICE_X15Y159_AQ;
  assign CLBLM_R_X11Y159_SLICE_X15Y159_A2 = CLBLM_L_X12Y159_SLICE_X17Y159_AO6;
  assign CLBLM_R_X11Y159_SLICE_X15Y159_A3 = CLBLM_L_X12Y158_SLICE_X17Y158_AQ;
  assign CLBLM_R_X11Y159_SLICE_X15Y159_A4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y159_SLICE_X15Y159_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y159_SLICE_X15Y159_A6 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_R_X11Y159_SLICE_X15Y159_B1 = CLBLM_L_X12Y150_SLICE_X16Y150_AQ;
  assign CLBLM_R_X11Y159_SLICE_X15Y159_B2 = CLBLM_R_X11Y159_SLICE_X15Y159_BQ;
  assign CLBLM_R_X11Y159_SLICE_X15Y159_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y159_SLICE_X15Y159_B4 = CLBLM_L_X10Y159_SLICE_X12Y159_CO6;
  assign CLBLM_R_X11Y159_SLICE_X15Y159_B5 = CLBLM_L_X10Y159_SLICE_X12Y159_DO6;
  assign CLBLM_R_X11Y159_SLICE_X15Y159_B6 = CLBLM_L_X10Y159_SLICE_X13Y159_DO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A1 = CLBLM_R_X7Y149_SLICE_X9Y149_CQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A3 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A5 = CLBLM_R_X5Y152_SLICE_X7Y152_AQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_A6 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X11Y159_SLICE_X15Y159_C1 = CLBLM_L_X12Y158_SLICE_X17Y158_AQ;
  assign CLBLM_R_X11Y159_SLICE_X15Y159_C2 = CLBLM_R_X11Y159_SLICE_X14Y159_BQ;
  assign CLBLM_R_X11Y159_SLICE_X15Y159_C3 = CLBLM_L_X12Y159_SLICE_X17Y159_AO5;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B2 = CLBLM_R_X7Y149_SLICE_X9Y149_BQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B3 = CLBLL_L_X4Y151_SLICE_X4Y151_BQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B4 = CLBLM_L_X10Y151_SLICE_X12Y151_CQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B5 = CLBLM_L_X8Y149_SLICE_X10Y149_AQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_B6 = CLBLM_R_X7Y149_SLICE_X9Y149_C5Q;
  assign CLBLM_R_X11Y159_SLICE_X15Y159_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y159_SLICE_X15Y159_D1 = CLBLM_R_X11Y159_SLICE_X14Y159_BQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C1 = CLBLM_R_X7Y149_SLICE_X9Y149_C5Q;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C2 = CLBLM_R_X11Y149_SLICE_X15Y149_A5Q;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C3 = CLBLM_R_X7Y156_SLICE_X9Y156_BQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C4 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_C6 = 1'b1;
  assign CLBLM_R_X11Y159_SLICE_X15Y159_D3 = CLBLM_L_X12Y155_SLICE_X16Y155_BO5;
  assign CLBLM_R_X11Y159_SLICE_X15Y159_D4 = CLBLM_L_X12Y159_SLICE_X17Y159_AO5;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y159_SLICE_X14Y159_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y159_SLICE_X14Y159_A2 = CLBLM_L_X8Y158_SLICE_X11Y158_BQ;
  assign CLBLM_R_X11Y159_SLICE_X14Y159_A3 = CLBLM_R_X11Y159_SLICE_X15Y159_CO5;
  assign CLBLM_R_X11Y159_SLICE_X14Y159_A4 = CLBLM_R_X11Y158_SLICE_X14Y158_DO6;
  assign CLBLM_R_X11Y159_SLICE_X14Y159_A5 = CLBLM_R_X11Y159_SLICE_X14Y159_AQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D1 = CLBLM_R_X3Y156_SLICE_X2Y156_DO6;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D2 = CLBLM_L_X8Y148_SLICE_X10Y148_CQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D3 = CLBLM_L_X8Y155_SLICE_X10Y155_B5Q;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D4 = CLBLM_R_X5Y149_SLICE_X7Y149_A5Q;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D5 = CLBLM_L_X10Y150_SLICE_X13Y150_BQ;
  assign CLBLM_R_X7Y149_SLICE_X9Y149_D6 = 1'b1;
  assign CLBLM_R_X11Y159_SLICE_X14Y159_A6 = CLBLM_L_X12Y159_SLICE_X16Y159_BO6;
  assign CLBLM_R_X11Y159_SLICE_X14Y159_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y159_SLICE_X14Y159_B2 = CLBLM_R_X11Y159_SLICE_X15Y159_DO6;
  assign CLBLM_R_X11Y159_SLICE_X14Y159_B3 = CLBLM_R_X11Y159_SLICE_X14Y159_BQ;
  assign CLBLM_R_X11Y159_SLICE_X14Y159_B4 = CLBLM_L_X12Y159_SLICE_X16Y159_BO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A1 = CLBLM_R_X7Y150_SLICE_X9Y150_CO6;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A3 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A5 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_A6 = CLBLL_L_X4Y149_SLICE_X5Y149_A5Q;
  assign CLBLM_R_X11Y159_SLICE_X14Y159_C1 = CLBLM_R_X11Y157_SLICE_X15Y157_AQ;
  assign CLBLM_R_X11Y159_SLICE_X14Y159_C2 = CLBLM_R_X11Y159_SLICE_X15Y159_AQ;
  assign CLBLM_R_X11Y159_SLICE_X14Y159_C3 = CLBLM_L_X12Y158_SLICE_X16Y158_AQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B2 = CLBLM_R_X7Y149_SLICE_X8Y149_BQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B4 = CLBLM_R_X5Y150_SLICE_X7Y150_CQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B5 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_B6 = CLBLM_L_X8Y149_SLICE_X11Y149_CQ;
  assign CLBLM_R_X11Y159_SLICE_X14Y159_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y159_SLICE_X14Y159_D1 = CLBLM_L_X10Y159_SLICE_X12Y159_DO6;
  assign CLBLM_R_X11Y159_SLICE_X14Y159_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C1 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C2 = CLBLM_R_X5Y149_SLICE_X7Y149_A5Q;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C3 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C4 = CLBLM_R_X5Y151_SLICE_X6Y151_CQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y159_SLICE_X14Y159_D3 = CLBLM_L_X10Y159_SLICE_X12Y159_CO6;
  assign CLBLM_R_X11Y159_SLICE_X14Y159_D4 = CLBLM_L_X12Y152_SLICE_X17Y152_A5Q;
  assign CLBLM_R_X11Y159_SLICE_X14Y159_D5 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y159_SLICE_X14Y159_D6 = CLBLM_L_X8Y159_SLICE_X11Y159_AO6;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A1 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D1 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D2 = CLBLM_R_X5Y149_SLICE_X7Y149_A5Q;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A2 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D4 = CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D6 = 1'b1;
  assign CLBLM_R_X7Y149_SLICE_X8Y149_D5 = CLBLL_L_X4Y154_SLICE_X5Y154_BO6;
  assign CLBLM_L_X8Y156_SLICE_X11Y156_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y156_SLICE_X11Y156_A2 = CLBLM_L_X8Y153_SLICE_X11Y153_C5Q;
  assign CLBLM_L_X8Y156_SLICE_X11Y156_A3 = CLBLM_L_X8Y156_SLICE_X11Y156_AQ;
  assign CLBLM_L_X8Y156_SLICE_X11Y156_A4 = CLBLM_R_X7Y155_SLICE_X8Y155_CO6;
  assign CLBLM_L_X8Y156_SLICE_X11Y156_A5 = CLBLM_L_X10Y153_SLICE_X12Y153_AQ;
  assign CLBLM_L_X8Y156_SLICE_X11Y156_A6 = CLBLM_R_X7Y158_SLICE_X8Y158_CO5;
  assign CLBLM_L_X8Y156_SLICE_X11Y156_B1 = CLBLM_R_X13Y155_SLICE_X18Y155_BQ;
  assign CLBLM_L_X8Y156_SLICE_X11Y156_B2 = CLBLM_L_X8Y156_SLICE_X11Y156_BQ;
  assign CLBLM_L_X8Y156_SLICE_X11Y156_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y156_SLICE_X11Y156_B4 = CLBLL_L_X4Y154_SLICE_X4Y154_BO6;
  assign CLBLM_L_X8Y156_SLICE_X11Y156_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y156_SLICE_X11Y156_B6 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C1 = 1'b1;
  assign LIOB33_X0Y173_IOB_X0Y173_O = CLBLM_R_X103Y141_SLICE_X163Y141_AO5;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C2 = 1'b1;
  assign CLBLM_L_X8Y156_SLICE_X11Y156_C1 = CLBLM_R_X7Y155_SLICE_X8Y155_BO5;
  assign CLBLM_L_X8Y156_SLICE_X11Y156_C2 = CLBLM_L_X8Y154_SLICE_X10Y154_A5Q;
  assign CLBLM_L_X8Y156_SLICE_X11Y156_C3 = CLBLM_L_X8Y158_SLICE_X10Y158_AQ;
  assign CLBLM_L_X8Y156_SLICE_X11Y156_C4 = CLBLM_R_X7Y148_SLICE_X8Y148_AQ;
  assign CLBLM_L_X8Y156_SLICE_X11Y156_C5 = CLBLM_L_X8Y150_SLICE_X11Y150_CQ;
  assign CLBLM_L_X8Y156_SLICE_X11Y156_C6 = CLBLM_R_X7Y148_SLICE_X8Y148_BQ;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C3 = 1'b1;
  assign CLBLM_R_X13Y159_SLICE_X19Y159_C4 = 1'b1;
  assign CLBLM_L_X8Y156_SLICE_X11Y156_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X13Y159_SLICE_X19Y159_C5 = 1'b1;
  assign CLBLM_R_X13Y159_SLICE_X19Y159_C6 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C5 = 1'b1;
  assign CLBLM_L_X8Y156_SLICE_X11Y156_D1 = CLBLM_L_X8Y158_SLICE_X10Y158_AQ;
  assign CLBLM_L_X8Y156_SLICE_X11Y156_D2 = CLBLM_L_X8Y154_SLICE_X10Y154_A5Q;
  assign CLBLM_L_X8Y156_SLICE_X11Y156_D3 = CLBLM_L_X8Y150_SLICE_X11Y150_CQ;
  assign CLBLM_L_X8Y156_SLICE_X11Y156_D4 = CLBLM_L_X10Y156_SLICE_X13Y156_AO6;
  assign CLBLM_L_X8Y156_SLICE_X11Y156_D5 = CLBLM_R_X7Y155_SLICE_X8Y155_AQ;
  assign CLBLM_L_X8Y156_SLICE_X11Y156_D6 = CLBLM_R_X7Y155_SLICE_X8Y155_BO5;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C6 = 1'b1;
  assign CLBLM_L_X8Y156_SLICE_X10Y156_A1 = CLBLM_R_X11Y159_SLICE_X14Y159_DQ;
  assign CLBLM_L_X8Y156_SLICE_X10Y156_A2 = CLBLM_L_X10Y155_SLICE_X12Y155_BQ;
  assign CLBLM_L_X8Y156_SLICE_X10Y156_A3 = CLBLM_L_X8Y156_SLICE_X10Y156_AQ;
  assign CLBLM_L_X8Y156_SLICE_X10Y156_A4 = CLBLL_L_X4Y151_SLICE_X4Y151_BQ;
  assign CLBLM_L_X8Y156_SLICE_X10Y156_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y156_SLICE_X10Y156_A6 = CLBLM_L_X10Y151_SLICE_X12Y151_CQ;
  assign CLBLM_L_X8Y156_SLICE_X10Y156_B1 = CLBLM_L_X12Y157_SLICE_X16Y157_BQ;
  assign CLBLM_L_X8Y156_SLICE_X10Y156_B2 = CLBLM_L_X8Y156_SLICE_X10Y156_BQ;
  assign CLBLM_L_X8Y156_SLICE_X10Y156_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y156_SLICE_X10Y156_B4 = CLBLM_L_X8Y155_SLICE_X10Y155_B5Q;
  assign CLBLM_L_X8Y156_SLICE_X10Y156_B5 = CLBLL_L_X4Y151_SLICE_X4Y151_BQ;
  assign CLBLM_L_X8Y156_SLICE_X10Y156_B6 = CLBLM_L_X10Y151_SLICE_X12Y151_CQ;
  assign CLBLM_L_X8Y156_SLICE_X10Y156_C1 = CLBLM_L_X8Y154_SLICE_X10Y154_BQ;
  assign CLBLM_L_X8Y156_SLICE_X10Y156_C2 = CLBLM_L_X8Y156_SLICE_X10Y156_CQ;
  assign CLBLM_L_X8Y156_SLICE_X10Y156_C3 = CLBLM_L_X10Y154_SLICE_X12Y154_DQ;
  assign CLBLM_L_X8Y156_SLICE_X10Y156_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y156_SLICE_X10Y156_C5 = CLBLM_L_X8Y156_SLICE_X10Y156_DO6;
  assign CLBLM_L_X8Y156_SLICE_X10Y156_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y156_SLICE_X10Y156_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y156_SLICE_X10Y156_D1 = CLBLM_L_X8Y155_SLICE_X11Y155_BQ;
  assign CLBLM_L_X8Y156_SLICE_X10Y156_D2 = 1'b1;
  assign CLBLM_L_X8Y156_SLICE_X10Y156_D3 = 1'b1;
  assign CLBLM_L_X8Y156_SLICE_X10Y156_D4 = CLBLM_L_X12Y158_SLICE_X16Y158_A5Q;
  assign CLBLM_L_X8Y156_SLICE_X10Y156_D5 = 1'b1;
  assign CLBLM_L_X8Y156_SLICE_X10Y156_D6 = 1'b1;
  assign CLBLM_R_X13Y159_SLICE_X19Y159_D3 = 1'b1;
  assign CLBLM_R_X13Y159_SLICE_X19Y159_D4 = 1'b1;
  assign CLBLM_R_X13Y159_SLICE_X19Y159_D5 = 1'b1;
  assign CLBLM_R_X13Y159_SLICE_X19Y159_D6 = 1'b1;
  assign CLBLM_R_X11Y160_SLICE_X15Y160_A1 = 1'b1;
  assign CLBLM_R_X11Y160_SLICE_X15Y160_A2 = 1'b1;
  assign CLBLM_R_X11Y160_SLICE_X15Y160_A3 = 1'b1;
  assign CLBLM_R_X11Y160_SLICE_X15Y160_A4 = 1'b1;
  assign CLBLM_R_X11Y160_SLICE_X15Y160_A5 = 1'b1;
  assign CLBLM_R_X11Y160_SLICE_X15Y160_A6 = 1'b1;
  assign CLBLM_R_X11Y160_SLICE_X15Y160_B1 = 1'b1;
  assign CLBLM_R_X11Y160_SLICE_X15Y160_B2 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_B5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X11Y160_SLICE_X15Y160_B3 = 1'b1;
  assign CLBLM_R_X11Y160_SLICE_X15Y160_B4 = 1'b1;
  assign CLBLM_R_X11Y160_SLICE_X15Y160_B5 = 1'b1;
  assign CLBLM_R_X11Y160_SLICE_X15Y160_B6 = 1'b1;
  assign CLBLM_R_X13Y159_SLICE_X18Y159_A1 = CLBLM_R_X11Y157_SLICE_X14Y157_AQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A1 = CLBLM_R_X11Y151_SLICE_X15Y151_AQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A2 = CLBLM_R_X7Y151_SLICE_X9Y151_AQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A3 = CLBLM_R_X7Y151_SLICE_X8Y151_DQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A4 = CLBLM_L_X10Y151_SLICE_X13Y151_AQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_A6 = 1'b1;
  assign CLBLM_R_X11Y160_SLICE_X15Y160_C1 = 1'b1;
  assign CLBLM_R_X11Y160_SLICE_X15Y160_C2 = 1'b1;
  assign CLBLM_R_X11Y160_SLICE_X15Y160_C3 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B1 = CLBLM_L_X10Y152_SLICE_X12Y152_CO5;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B2 = CLBLM_R_X3Y156_SLICE_X2Y156_DO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B3 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B5 = CLBLM_R_X7Y152_SLICE_X9Y152_CO5;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_B6 = CLBLM_R_X11Y149_SLICE_X15Y149_A5Q;
  assign CLBLM_R_X11Y160_SLICE_X15Y160_D1 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C1 = CLBLM_R_X7Y152_SLICE_X9Y152_CO5;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C2 = CLBLM_R_X7Y154_SLICE_X8Y154_AO5;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_C1 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C3 = CLBLL_L_X4Y153_SLICE_X4Y153_AO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C4 = CLBLM_R_X7Y150_SLICE_X9Y150_AO5;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C5 = CLBLM_L_X10Y152_SLICE_X12Y152_CO5;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y140_SLICE_X0Y140_C2 = 1'b1;
  assign CLBLM_R_X11Y160_SLICE_X14Y160_A1 = 1'b1;
  assign CLBLM_R_X11Y160_SLICE_X14Y160_A2 = CLBLM_L_X10Y158_SLICE_X13Y158_CO6;
  assign CLBLM_R_X11Y160_SLICE_X14Y160_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y160_SLICE_X14Y160_A4 = 1'b1;
  assign CLBLM_R_X11Y160_SLICE_X14Y160_A5 = CLBLM_L_X10Y159_SLICE_X12Y159_CO6;
  assign CLBLM_R_X11Y160_SLICE_X14Y160_A6 = CLBLM_R_X11Y159_SLICE_X14Y159_AQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D1 = CLBLM_R_X5Y147_SLICE_X7Y147_C5Q;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D2 = CLBLM_R_X5Y146_SLICE_X6Y146_A5Q;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D3 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D4 = CLBLM_R_X7Y152_SLICE_X9Y152_BQ;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D5 = CLBLM_L_X10Y156_SLICE_X13Y156_AO6;
  assign CLBLM_R_X7Y150_SLICE_X9Y150_D6 = CLBLM_R_X13Y150_SLICE_X18Y150_DO5;
  assign CLBLM_R_X11Y160_SLICE_X14Y160_B1 = 1'b1;
  assign CLBLM_R_X11Y160_SLICE_X14Y160_B2 = 1'b1;
  assign CLBLM_R_X11Y160_SLICE_X14Y160_B3 = 1'b1;
  assign CLBLM_R_X11Y160_SLICE_X14Y160_B4 = 1'b1;
  assign CLBLM_R_X11Y160_SLICE_X14Y160_B5 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A1 = CLBLM_R_X7Y150_SLICE_X8Y150_DO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A2 = CLBLM_R_X7Y155_SLICE_X9Y155_AQ;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A3 = CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_A6 = 1'b1;
  assign CLBLM_R_X11Y160_SLICE_X14Y160_C1 = 1'b1;
  assign CLBLM_R_X11Y160_SLICE_X14Y160_C2 = 1'b1;
  assign CLBLM_R_X11Y160_SLICE_X14Y160_C3 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B2 = CLBLM_L_X10Y150_SLICE_X13Y150_BQ;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B3 = CLBLM_R_X7Y156_SLICE_X9Y156_BQ;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B5 = CLBLM_R_X7Y150_SLICE_X8Y150_CO5;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_B6 = 1'b1;
  assign CLBLM_R_X11Y160_SLICE_X14Y160_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y160_SLICE_X14Y160_D1 = 1'b1;
  assign CLBLM_R_X11Y160_SLICE_X14Y160_D2 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C1 = CLBLM_L_X8Y150_SLICE_X11Y150_BQ;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C2 = CLBLM_R_X5Y152_SLICE_X6Y152_BQ;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C3 = CLBLL_L_X4Y150_SLICE_X4Y150_BQ;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C4 = CLBLM_L_X10Y149_SLICE_X12Y149_C5Q;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_C6 = 1'b1;
  assign CLBLM_R_X11Y160_SLICE_X14Y160_D3 = 1'b1;
  assign CLBLM_R_X11Y160_SLICE_X14Y160_D4 = 1'b1;
  assign CLBLM_R_X11Y160_SLICE_X14Y160_D5 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y160_SLICE_X14Y160_D6 = 1'b1;
  assign CLBLM_R_X13Y159_SLICE_X18Y159_B5 = CLBLM_R_X13Y157_SLICE_X19Y157_AQ;
  assign CLBLM_R_X13Y159_SLICE_X18Y159_B6 = CLBLM_R_X11Y157_SLICE_X14Y157_AQ;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D1 = 1'b1;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D2 = CLBLL_L_X4Y150_SLICE_X5Y150_DQ;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D3 = CLBLM_R_X7Y152_SLICE_X9Y152_DO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D4 = CLBLM_R_X7Y152_SLICE_X8Y152_A5Q;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D5 = CLBLM_R_X5Y150_SLICE_X7Y150_DO6;
  assign CLBLM_R_X7Y150_SLICE_X8Y150_D6 = CLBLM_R_X7Y151_SLICE_X9Y151_DO6;
  assign CLBLM_R_X13Y159_SLICE_X18Y159_C1 = CLBLM_L_X12Y157_SLICE_X17Y157_BQ;
  assign CLBLM_R_X13Y159_SLICE_X18Y159_C2 = CLBLM_L_X12Y158_SLICE_X17Y158_AQ;
  assign CLBLM_R_X13Y159_SLICE_X18Y159_C3 = CLBLM_L_X12Y156_SLICE_X17Y156_AQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C1 = CLBLM_R_X5Y146_SLICE_X6Y146_AQ;
  assign CLBLM_R_X13Y159_SLICE_X18Y159_C4 = CLBLM_L_X12Y158_SLICE_X16Y158_AQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C2 = CLBLM_R_X5Y146_SLICE_X6Y146_A5Q;
  assign CLBLM_R_X13Y159_SLICE_X18Y159_C5 = CLBLM_R_X11Y159_SLICE_X15Y159_AQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C3 = CLBLM_R_X5Y144_SLICE_X6Y144_BQ;
  assign CLBLM_R_X13Y159_SLICE_X18Y159_C6 = CLBLM_L_X8Y154_SLICE_X10Y154_AQ;
  assign LIOB33_X0Y175_IOB_X0Y176_O = RIOB33_X105Y127_IOB_X1Y128_I;
  assign LIOB33_X0Y175_IOB_X0Y175_O = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_L_X8Y157_SLICE_X11Y157_A1 = CLBLM_R_X11Y149_SLICE_X15Y149_AQ;
  assign CLBLM_L_X8Y157_SLICE_X11Y157_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y157_SLICE_X11Y157_A3 = CLBLM_R_X7Y158_SLICE_X8Y158_CO5;
  assign CLBLM_L_X8Y157_SLICE_X11Y157_A4 = CLBLM_R_X7Y155_SLICE_X8Y155_CO6;
  assign CLBLM_L_X8Y157_SLICE_X11Y157_A5 = CLBLM_L_X8Y158_SLICE_X11Y158_AQ;
  assign CLBLM_L_X8Y157_SLICE_X11Y157_A6 = CLBLM_L_X8Y157_SLICE_X11Y157_AQ;
  assign CLBLM_L_X8Y157_SLICE_X11Y157_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y157_SLICE_X11Y157_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y157_SLICE_X11Y157_B3 = 1'b1;
  assign CLBLM_L_X8Y157_SLICE_X11Y157_B4 = CLBLM_L_X10Y156_SLICE_X13Y156_BQ;
  assign CLBLM_L_X8Y157_SLICE_X11Y157_B5 = 1'b1;
  assign CLBLM_L_X8Y157_SLICE_X11Y157_B6 = CLBLM_L_X10Y157_SLICE_X12Y157_AQ;
  assign CLBLM_L_X8Y157_SLICE_X11Y157_C1 = 1'b1;
  assign CLBLM_L_X8Y157_SLICE_X11Y157_C2 = CLBLM_L_X8Y157_SLICE_X11Y157_CQ;
  assign CLBLM_L_X8Y157_SLICE_X11Y157_C3 = CLBLM_R_X13Y158_SLICE_X18Y158_BQ;
  assign CLBLM_L_X8Y157_SLICE_X11Y157_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y157_SLICE_X11Y157_C5 = 1'b1;
  assign CLBLM_L_X8Y157_SLICE_X11Y157_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y159_SLICE_X18Y159_D1 = CLBLM_L_X12Y157_SLICE_X17Y157_BQ;
  assign CLBLM_R_X13Y159_SLICE_X18Y159_D2 = CLBLM_L_X12Y158_SLICE_X17Y158_AQ;
  assign CLBLM_L_X8Y157_SLICE_X11Y157_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X13Y159_SLICE_X18Y159_D3 = CLBLM_L_X12Y156_SLICE_X17Y156_AQ;
  assign CLBLM_L_X8Y157_SLICE_X11Y157_D1 = CLBLM_R_X7Y148_SLICE_X8Y148_AQ;
  assign CLBLM_L_X8Y157_SLICE_X11Y157_D2 = CLBLM_L_X8Y158_SLICE_X10Y158_AQ;
  assign CLBLM_L_X8Y157_SLICE_X11Y157_D3 = CLBLM_R_X7Y155_SLICE_X8Y155_BO5;
  assign CLBLM_L_X8Y157_SLICE_X11Y157_D4 = CLBLM_L_X8Y154_SLICE_X10Y154_A5Q;
  assign CLBLM_L_X8Y157_SLICE_X11Y157_D5 = CLBLM_R_X7Y155_SLICE_X8Y155_AQ;
  assign CLBLM_L_X8Y157_SLICE_X11Y157_D6 = CLBLM_R_X7Y148_SLICE_X8Y148_BQ;
  assign CLBLM_R_X13Y159_SLICE_X18Y159_D5 = CLBLM_R_X11Y159_SLICE_X15Y159_AQ;
  assign CLBLM_L_X8Y157_SLICE_X10Y157_A1 = CLBLM_R_X11Y158_SLICE_X14Y158_CQ;
  assign CLBLM_L_X8Y157_SLICE_X10Y157_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X8Y157_SLICE_X10Y157_A3 = CLBLL_L_X4Y158_SLICE_X4Y158_AO6;
  assign CLBLM_L_X8Y157_SLICE_X10Y157_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y157_SLICE_X10Y157_A5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X8Y157_SLICE_X10Y157_A6 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X8Y157_SLICE_X10Y157_B1 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X8Y157_SLICE_X10Y157_B2 = CLBLM_L_X8Y157_SLICE_X10Y157_BQ;
  assign CLBLM_L_X8Y157_SLICE_X10Y157_B3 = CLBLM_L_X8Y156_SLICE_X11Y156_AQ;
  assign CLBLM_L_X8Y157_SLICE_X10Y157_B4 = CLBLM_R_X7Y155_SLICE_X8Y155_CO6;
  assign CLBLM_L_X8Y157_SLICE_X10Y157_B5 = CLBLM_R_X7Y158_SLICE_X8Y158_CO5;
  assign CLBLM_L_X8Y157_SLICE_X10Y157_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y157_SLICE_X10Y157_C1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y157_SLICE_X10Y157_C2 = CLBLM_L_X8Y157_SLICE_X10Y157_CQ;
  assign CLBLM_L_X8Y157_SLICE_X10Y157_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y157_SLICE_X10Y157_C4 = CLBLM_L_X12Y149_SLICE_X16Y149_CQ;
  assign CLBLM_L_X8Y157_SLICE_X10Y157_C5 = CLBLM_L_X8Y150_SLICE_X11Y150_CQ;
  assign CLBLM_L_X8Y157_SLICE_X10Y157_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y157_SLICE_X10Y157_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_D1 = CLBLM_R_X103Y141_SLICE_X163Y141_AO6;
  assign CLBLM_L_X8Y157_SLICE_X10Y157_D1 = CLBLM_R_X5Y149_SLICE_X6Y149_BQ;
  assign CLBLM_L_X8Y157_SLICE_X10Y157_D2 = CLBLM_R_X11Y158_SLICE_X14Y158_CQ;
  assign CLBLM_L_X8Y157_SLICE_X10Y157_D3 = 1'b1;
  assign CLBLM_L_X8Y157_SLICE_X10Y157_D4 = CLBLM_R_X11Y159_SLICE_X15Y159_CO6;
  assign CLBLM_L_X8Y157_SLICE_X10Y157_D5 = 1'b1;
  assign CLBLM_L_X8Y157_SLICE_X10Y157_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_D = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y172_T1 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_D1 = CLBLM_R_X3Y142_SLICE_X3Y142_BO6;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_D1 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_X0Y109_OLOGIC_X0Y110_T1 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_D1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign LIOI3_X0Y171_OLOGIC_X0Y171_T1 = 1'b1;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_D1 = CLBLM_R_X3Y142_SLICE_X3Y142_DO6;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_D3 = 1'b1;
  assign RIOI3_X105Y153_OLOGIC_X1Y154_T1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = CLBLM_R_X5Y146_SLICE_X6Y146_BQ;
  assign LIOI3_X0Y109_OLOGIC_X0Y109_T1 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C5 = CLBLM_R_X11Y159_SLICE_X14Y159_CQ;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_D1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A1 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_D4 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A3 = CLBLM_R_X7Y151_SLICE_X9Y151_AQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A4 = CLBLM_L_X8Y153_SLICE_X10Y153_BO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_A6 = CLBLM_L_X8Y152_SLICE_X10Y152_CQ;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = CLBLM_R_X5Y144_SLICE_X6Y144_BQ;
  assign RIOI3_X105Y153_OLOGIC_X1Y153_T1 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B1 = CLBLM_L_X8Y151_SLICE_X10Y151_CQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B3 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B4 = CLBLM_L_X8Y151_SLICE_X11Y151_CO6;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B5 = CLBLM_L_X10Y152_SLICE_X12Y152_AQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C1 = CLBLM_R_X7Y155_SLICE_X9Y155_AQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C2 = CLBLM_R_X5Y151_SLICE_X6Y151_BQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C3 = CLBLM_R_X11Y151_SLICE_X15Y151_AQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_C6 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D1 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D2 = CLBLL_L_X4Y150_SLICE_X4Y150_CQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D3 = CLBLM_R_X7Y151_SLICE_X9Y151_BQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D4 = CLBLM_R_X7Y154_SLICE_X9Y154_CQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D5 = CLBLM_R_X7Y152_SLICE_X9Y152_BQ;
  assign CLBLM_R_X7Y151_SLICE_X9Y151_D6 = CLBLM_R_X7Y151_SLICE_X8Y151_BQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A1 = CLBLM_L_X10Y151_SLICE_X13Y151_DO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A3 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A5 = CLBLM_L_X8Y151_SLICE_X11Y151_AQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_A6 = CLBLM_R_X7Y148_SLICE_X8Y148_CQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B1 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B2 = CLBLM_R_X7Y149_SLICE_X8Y149_BQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B3 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B4 = CLBLM_L_X8Y153_SLICE_X10Y153_BO6;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C1 = CLBLM_R_X7Y150_SLICE_X8Y150_BQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C2 = CLBLM_R_X7Y151_SLICE_X8Y151_CQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C4 = CLBLM_R_X7Y151_SLICE_X9Y151_CQ;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_C4 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C5 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D1 = CLBLM_R_X7Y157_SLICE_X8Y157_BQ;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D3 = CLBLM_R_X7Y151_SLICE_X9Y151_C5Q;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D4 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D5 = 1'b1;
  assign CLBLM_R_X7Y151_SLICE_X8Y151_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOB33_X0Y177_IOB_X0Y178_O = RIOB33_X105Y129_IOB_X1Y130_I;
  assign LIOB33_X0Y177_IOB_X0Y177_O = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_D1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D3 = 1'b1;
  assign LIOB33_X0Y131_IOB_X0Y132_O = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D4 = 1'b1;
  assign CLBLL_L_X2Y140_SLICE_X1Y140_D4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D6 = 1'b1;
  assign CLBLM_L_X8Y158_SLICE_X11Y158_A1 = CLBLM_L_X8Y157_SLICE_X10Y157_BQ;
  assign CLBLM_L_X8Y158_SLICE_X11Y158_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y158_SLICE_X11Y158_A3 = CLBLM_L_X8Y158_SLICE_X11Y158_AQ;
  assign CLBLM_L_X8Y158_SLICE_X11Y158_A4 = CLBLM_R_X7Y155_SLICE_X8Y155_CO6;
  assign CLBLM_L_X8Y158_SLICE_X11Y158_A5 = CLBLM_R_X7Y158_SLICE_X8Y158_CO5;
  assign CLBLM_L_X8Y158_SLICE_X11Y158_A6 = CLBLM_R_X7Y156_SLICE_X8Y156_DQ;
  assign LIOB33_X0Y131_IOB_X0Y131_O = CLBLM_L_X10Y144_SLICE_X12Y144_AO5;
  assign CLBLM_L_X8Y158_SLICE_X11Y158_B1 = 1'b1;
  assign CLBLM_L_X8Y158_SLICE_X11Y158_B2 = CLBLM_L_X8Y158_SLICE_X11Y158_BQ;
  assign CLBLM_L_X8Y158_SLICE_X11Y158_B3 = CLBLM_L_X10Y153_SLICE_X12Y153_BQ;
  assign CLBLM_L_X8Y158_SLICE_X11Y158_B4 = CLBLM_R_X11Y152_SLICE_X14Y152_B5Q;
  assign CLBLM_L_X8Y158_SLICE_X11Y158_B5 = CLBLM_R_X5Y152_SLICE_X6Y152_CO5;
  assign CLBLM_L_X8Y158_SLICE_X11Y158_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y158_SLICE_X11Y158_C1 = 1'b1;
  assign CLBLM_L_X8Y158_SLICE_X11Y158_C2 = 1'b1;
  assign CLBLM_L_X8Y158_SLICE_X11Y158_C3 = 1'b1;
  assign CLBLM_L_X8Y158_SLICE_X11Y158_C4 = 1'b1;
  assign CLBLM_L_X8Y158_SLICE_X11Y158_C5 = 1'b1;
  assign CLBLM_L_X8Y158_SLICE_X11Y158_C6 = 1'b1;
  assign CLBLM_L_X8Y158_SLICE_X11Y158_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y158_SLICE_X11Y158_D1 = 1'b1;
  assign CLBLM_L_X8Y158_SLICE_X11Y158_D2 = 1'b1;
  assign CLBLM_L_X8Y158_SLICE_X11Y158_D3 = 1'b1;
  assign CLBLM_L_X8Y158_SLICE_X11Y158_D4 = 1'b1;
  assign CLBLM_L_X8Y158_SLICE_X11Y158_D5 = 1'b1;
  assign CLBLM_L_X8Y158_SLICE_X11Y158_D6 = 1'b1;
  assign CLBLM_L_X8Y158_SLICE_X10Y158_A1 = CLBLM_L_X8Y159_SLICE_X10Y159_BO5;
  assign CLBLM_L_X8Y158_SLICE_X10Y158_A2 = CLBLM_L_X10Y159_SLICE_X12Y159_AO6;
  assign CLBLM_L_X8Y158_SLICE_X10Y158_A3 = CLBLM_L_X8Y158_SLICE_X10Y158_AQ;
  assign CLBLM_L_X8Y158_SLICE_X10Y158_A4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X8Y158_SLICE_X10Y158_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y158_SLICE_X10Y158_A6 = CLBLM_L_X8Y156_SLICE_X10Y156_CQ;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A6 = 1'b1;
  assign CLBLM_L_X8Y158_SLICE_X10Y158_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y158_SLICE_X10Y158_B2 = CLBLM_L_X8Y158_SLICE_X10Y158_BQ;
  assign CLBLM_L_X8Y158_SLICE_X10Y158_B3 = 1'b1;
  assign CLBLM_L_X8Y158_SLICE_X10Y158_B4 = CLBLM_R_X7Y158_SLICE_X9Y158_AQ;
  assign CLBLM_L_X8Y158_SLICE_X10Y158_B5 = 1'b1;
  assign CLBLM_L_X8Y158_SLICE_X10Y158_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y158_SLICE_X10Y158_C1 = 1'b1;
  assign CLBLM_L_X8Y158_SLICE_X10Y158_C2 = 1'b1;
  assign CLBLM_L_X8Y158_SLICE_X10Y158_C3 = 1'b1;
  assign CLBLM_L_X8Y158_SLICE_X10Y158_C4 = 1'b1;
  assign CLBLM_L_X8Y158_SLICE_X10Y158_C5 = 1'b1;
  assign CLBLM_L_X8Y158_SLICE_X10Y158_C6 = 1'b1;
  assign CLBLM_L_X8Y158_SLICE_X10Y158_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y158_SLICE_X10Y158_D1 = 1'b1;
  assign CLBLM_L_X8Y158_SLICE_X10Y158_D2 = 1'b1;
  assign CLBLM_L_X8Y158_SLICE_X10Y158_D3 = 1'b1;
  assign CLBLM_L_X8Y158_SLICE_X10Y158_D4 = 1'b1;
  assign CLBLM_L_X8Y158_SLICE_X10Y158_D5 = 1'b1;
  assign CLBLM_L_X8Y158_SLICE_X10Y158_D6 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C2 = CLBLM_R_X11Y150_SLICE_X14Y150_BO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B4 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_C5 = CLBLM_L_X12Y151_SLICE_X17Y151_A5Q;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B6 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X54Y150_A1 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X54Y150_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X36Y150_SLICE_X54Y150_A3 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X54Y150_A4 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLL_L_X36Y150_SLICE_X54Y150_A5 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X54Y150_A6 = CLBLM_R_X7Y149_SLICE_X9Y149_CQ;
  assign CLBLM_R_X11Y151_SLICE_X15Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLL_L_X36Y150_SLICE_X54Y150_B1 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X54Y150_B2 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X54Y150_B3 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X54Y150_B4 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X54Y150_B5 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X54Y150_B6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D3 = 1'b1;
  assign RIOI3_SING_X105Y149_ILOGIC_X1Y149_D = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLL_L_X36Y150_SLICE_X54Y150_C1 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X54Y150_C2 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X54Y150_C3 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X54Y150_C4 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X54Y150_C5 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X54Y150_C6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_A1 = CLBLM_R_X5Y152_SLICE_X6Y152_CO6;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_A2 = CLBLM_R_X7Y152_SLICE_X9Y152_BQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_A3 = CLBLM_R_X7Y152_SLICE_X9Y152_AQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_A4 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_A6 = CLBLM_L_X12Y152_SLICE_X16Y152_BQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_B1 = CLBLM_L_X8Y152_SLICE_X10Y152_DO6;
  assign CLBLL_L_X36Y150_SLICE_X54Y150_D1 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X54Y150_D2 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X54Y150_D3 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X54Y150_D4 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X54Y150_D5 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X54Y150_D6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_B4 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_B5 = CLBLM_R_X13Y154_SLICE_X19Y154_AQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_B6 = CLBLM_R_X7Y154_SLICE_X9Y154_CQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_C1 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_C2 = CLBLM_R_X3Y155_SLICE_X2Y155_BO6;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_C4 = CLBLM_R_X7Y150_SLICE_X8Y150_CO6;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_C5 = CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_C6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_D1 = CLBLM_R_X5Y154_SLICE_X6Y154_AQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_D2 = CLBLM_R_X7Y153_SLICE_X9Y153_CO5;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_D3 = CLBLM_L_X10Y157_SLICE_X12Y157_AQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_D5 = CLBLM_L_X8Y151_SLICE_X11Y151_AQ;
  assign CLBLM_R_X7Y152_SLICE_X9Y152_D6 = CLBLM_L_X8Y157_SLICE_X11Y157_BQ;
  assign CLBLL_L_X36Y150_SLICE_X55Y150_A1 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X55Y150_A2 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X55Y150_A3 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X55Y150_A4 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X55Y150_A5 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X55Y150_A6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_A1 = CLBLM_R_X7Y155_SLICE_X8Y155_DO6;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_A2 = CLBLM_R_X7Y151_SLICE_X8Y151_BQ;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_A3 = CLBLM_R_X7Y152_SLICE_X8Y152_AQ;
  assign CLBLL_L_X36Y150_SLICE_X55Y150_B1 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X55Y150_B2 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X55Y150_B3 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X55Y150_B4 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X55Y150_B5 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X55Y150_B6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_A6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_AX = CLBLM_R_X7Y152_SLICE_X8Y152_BO6;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_B1 = CLBLM_L_X8Y157_SLICE_X10Y157_DQ;
  assign CLBLL_L_X36Y150_SLICE_X55Y150_C1 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X55Y150_C2 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X55Y150_C3 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X55Y150_C4 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X55Y150_C5 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X55Y150_C6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_B5 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_B6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_C1 = CLBLM_R_X7Y148_SLICE_X8Y148_AQ;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_C2 = CLBLM_R_X7Y150_SLICE_X9Y150_DO6;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_C3 = CLBLM_L_X8Y158_SLICE_X10Y158_AQ;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_C4 = CLBLM_L_X8Y148_SLICE_X10Y148_DO6;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_C5 = CLBLM_R_X7Y152_SLICE_X8Y152_DO6;
  assign CLBLL_L_X36Y150_SLICE_X55Y150_D1 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X55Y150_D2 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X55Y150_D3 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X55Y150_D4 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X55Y150_D5 = 1'b1;
  assign CLBLL_L_X36Y150_SLICE_X55Y150_D6 = 1'b1;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_D1 = CLBLM_R_X5Y150_SLICE_X7Y150_AQ;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_D2 = CLBLM_R_X7Y157_SLICE_X9Y157_DQ;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_D3 = CLBLM_L_X10Y150_SLICE_X13Y150_BQ;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_D4 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y152_SLICE_X8Y152_D6 = CLBLM_R_X5Y151_SLICE_X7Y151_CQ;
  assign LIOB33_X0Y179_IOB_X0Y179_O = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOB33_X0Y179_IOB_X0Y180_O = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0 = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_A1 = CLBLM_L_X8Y157_SLICE_X11Y157_DO6;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_A2 = CLBLM_L_X10Y159_SLICE_X12Y159_BO6;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_A3 = CLBLM_L_X8Y157_SLICE_X11Y157_AQ;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_A4 = CLBLM_L_X10Y159_SLICE_X13Y159_BO5;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_A5 = CLBLM_L_X8Y156_SLICE_X11Y156_DO6;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_A6 = CLBLM_R_X11Y159_SLICE_X14Y159_DQ;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_T1 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_B1 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_B2 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_B3 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_B4 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_B5 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_B6 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_C1 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_C2 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_C3 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_C4 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_C5 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_C6 = 1'b1;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_B1 = CLBLM_L_X12Y156_SLICE_X17Y156_AQ;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_D1 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_D2 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_D3 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_D4 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_D5 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X11Y159_D6 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_A1 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_A2 = CLBLM_R_X7Y149_SLICE_X9Y149_DO6;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_A3 = CLBLM_R_X7Y158_SLICE_X8Y158_CO5;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_A4 = CLBLM_R_X7Y159_SLICE_X9Y159_AO6;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_A6 = CLBLM_R_X11Y159_SLICE_X15Y159_AQ;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_B1 = CLBLM_R_X7Y148_SLICE_X8Y148_AQ;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_B2 = CLBLM_R_X7Y148_SLICE_X8Y148_BQ;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_B3 = CLBLM_L_X8Y154_SLICE_X10Y154_A5Q;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_B4 = CLBLM_R_X7Y155_SLICE_X8Y155_AQ;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_B5 = CLBLM_L_X8Y158_SLICE_X10Y158_AQ;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_B6 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_C1 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_C2 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_C3 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_C4 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_C5 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_C6 = 1'b1;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_D1 = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_D1 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_D2 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_D3 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_D4 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_D5 = 1'b1;
  assign CLBLM_L_X8Y159_SLICE_X10Y159_D6 = 1'b1;
  assign RIOI3_SING_X105Y150_OLOGIC_X1Y150_T1 = 1'b1;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D4 = CLBLM_L_X12Y153_SLICE_X17Y153_BQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D5 = 1'b1;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_B1 = CLBLM_R_X3Y156_SLICE_X3Y156_AO5;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B4 = CLBLM_L_X10Y146_SLICE_X12Y146_AQ;
  assign CLBLM_R_X11Y151_SLICE_X14Y151_D6 = CLBLM_L_X10Y151_SLICE_X12Y151_AQ;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_B2 = CLBLM_R_X7Y155_SLICE_X8Y155_A5Q;
  assign CLBLM_L_X8Y147_SLICE_X11Y147_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_A1 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_A2 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_A3 = CLBLM_R_X7Y153_SLICE_X9Y153_AQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_A6 = CLBLL_L_X4Y156_SLICE_X4Y156_AQ;
  assign CLBLM_L_X10Y163_SLICE_X12Y163_A6 = 1'b1;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_B2 = CLBLM_R_X11Y158_SLICE_X15Y158_DO6;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_B1 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_B2 = CLBLM_R_X7Y153_SLICE_X9Y153_BQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_B4 = CLBLM_R_X5Y150_SLICE_X7Y150_A5Q;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_B5 = CLBLM_L_X10Y158_SLICE_X13Y158_AQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_B6 = CLBLL_L_X4Y147_SLICE_X4Y147_BO6;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_C1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_C3 = CLBLM_L_X12Y149_SLICE_X16Y149_CQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_C4 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_C5 = CLBLM_R_X13Y150_SLICE_X18Y150_AQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_C6 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_D1 = CLBLL_L_X4Y153_SLICE_X5Y153_AQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_D2 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_D3 = CLBLM_R_X5Y150_SLICE_X6Y150_AQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_D4 = CLBLM_L_X10Y150_SLICE_X13Y150_CQ;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_D5 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X9Y153_D6 = CLBLM_L_X10Y153_SLICE_X12Y153_BQ;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_A1 = CLBLM_L_X8Y157_SLICE_X10Y157_AQ;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_A2 = CLBLL_L_X4Y148_SLICE_X5Y148_DQ;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_A4 = CLBLM_L_X8Y158_SLICE_X10Y158_AQ;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_A5 = CLBLM_L_X12Y150_SLICE_X16Y150_CQ;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_A6 = 1'b1;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_D1 = CLBLM_L_X10Y163_SLICE_X13Y163_AO6;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_B1 = CLBLM_R_X7Y156_SLICE_X8Y156_CQ;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_B2 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_B4 = CLBLM_L_X10Y151_SLICE_X13Y151_BQ;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_B5 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOB33_X0Y181_IOB_X0Y181_O = RIOB33_X105Y133_IOB_X1Y133_I;
  assign LIOB33_X0Y181_IOB_X0Y182_O = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_D1 = CLBLM_L_X12Y151_SLICE_X16Y151_C5Q;
  assign LIOI3_X0Y173_OLOGIC_X0Y174_T1 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_C1 = CLBLM_L_X10Y148_SLICE_X13Y148_AQ;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_C2 = CLBLM_R_X7Y153_SLICE_X8Y153_CQ;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_C3 = CLBLM_R_X7Y155_SLICE_X9Y155_A5Q;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_C4 = CLBLM_L_X10Y150_SLICE_X12Y150_A5Q;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_C5 = CLBLM_L_X12Y155_SLICE_X16Y155_CO6;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y111_OLOGIC_X0Y112_T1 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_D1 = CLBLM_R_X103Y141_SLICE_X163Y141_AO5;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_D1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign LIOI3_X0Y173_OLOGIC_X0Y173_T1 = 1'b1;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_D1 = CLBLM_R_X3Y151_SLICE_X2Y151_CO5;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_D2 = CLBLM_R_X7Y152_SLICE_X8Y152_CO6;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_D3 = CLBLM_R_X13Y156_SLICE_X18Y156_CO6;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_D4 = CLBLM_R_X7Y155_SLICE_X8Y155_BO6;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_D5 = CLBLM_L_X8Y155_SLICE_X11Y155_DO6;
  assign CLBLM_R_X7Y153_SLICE_X8Y153_D6 = CLBLM_R_X7Y153_SLICE_X9Y153_BQ;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_D1 = 1'b0;
  assign RIOI3_X105Y155_OLOGIC_X1Y156_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_D1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_T1 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_D1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y164_T1 = 1'b1;
  assign RIOI3_X105Y155_OLOGIC_X1Y155_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_D1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X4Y153_SLICE_X5Y153_D5 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y163_OLOGIC_X0Y163_T1 = 1'b1;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_D1 = CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign CLBLM_L_X10Y163_SLICE_X12Y163_B4 = 1'b1;
  assign CLBLM_L_X10Y163_SLICE_X12Y163_B5 = 1'b1;
  assign LIOI3_X0Y51_ILOGIC_X0Y52_D = LIOB33_X0Y51_IOB_X0Y52_I;
  assign CLBLM_L_X10Y163_SLICE_X12Y163_B6 = 1'b1;
  assign LIOI3_X0Y51_ILOGIC_X0Y51_D = LIOB33_X0Y51_IOB_X0Y51_I;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_D1 = CLBLM_R_X13Y156_SLICE_X19Y156_AQ;
  assign RIOB33_X105Y151_IOB_X1Y152_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOB33_X105Y151_IOB_X1Y151_O = LIOB33_X0Y75_IOB_X0Y76_I;
  assign RIOI3_SING_X105Y199_OLOGIC_X1Y199_T1 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_A1 = CLBLM_R_X7Y154_SLICE_X9Y154_AQ;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_A2 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_A4 = CLBLM_R_X11Y146_SLICE_X15Y146_AQ;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_A5 = CLBLM_R_X5Y152_SLICE_X6Y152_CO5;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_A6 = CLBLL_L_X4Y150_SLICE_X4Y150_CQ;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y58_D = LIOB33_X0Y57_IOB_X0Y58_I;
  assign LIOI3_TBYTESRC_X0Y57_ILOGIC_X0Y57_D = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_A1 = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_A2 = CLBLL_L_X4Y157_SLICE_X4Y157_CO6;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_A5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_A6 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_B1 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_B2 = CLBLM_R_X7Y154_SLICE_X9Y154_BQ;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_B1 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_B2 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A3 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A4 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A5 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_A6 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_B3 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_B4 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_B5 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_B6 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_C1 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_C2 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_C3 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_C4 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_C5 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_C6 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B1 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B2 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B3 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B4 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B5 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_B6 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_D1 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_D2 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_D3 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_D4 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_D5 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X0Y153_D6 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_C4 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D1 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D2 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D3 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D4 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D5 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X7Y144_D6 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_A5 = CLBLL_L_X4Y150_SLICE_X4Y150_CQ;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_A6 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_B1 = CLBLM_R_X7Y155_SLICE_X8Y155_CO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_B2 = CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_B3 = CLBLM_L_X8Y157_SLICE_X11Y157_AQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A1 = CLBLM_R_X5Y144_SLICE_X6Y144_DO6;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A3 = CLBLM_R_X5Y144_SLICE_X6Y144_AQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A4 = CLBLM_R_X11Y155_SLICE_X14Y155_CQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_A6 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_C1 = CLBLM_R_X7Y148_SLICE_X8Y148_AQ;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_C2 = CLBLM_R_X7Y148_SLICE_X8Y148_BQ;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B5 = CLBLM_R_X5Y144_SLICE_X6Y144_CO5;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_A4 = CLBLL_L_X4Y157_SLICE_X4Y157_CO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_A5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_A6 = 1'b1;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B2 = CLBLM_R_X5Y144_SLICE_X6Y144_BQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B3 = CLBLM_R_X5Y153_SLICE_X7Y153_AQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_B4 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_B1 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C4 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C5 = CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_C6 = 1'b1;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_B2 = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_B3 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_B4 = CLBLM_R_X3Y153_SLICE_X2Y153_CO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_B5 = CLBLL_L_X2Y153_SLICE_X1Y153_AO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_B6 = CLBLL_L_X2Y154_SLICE_X1Y154_AO5;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_C1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_C2 = CLBLM_R_X3Y152_SLICE_X2Y152_AO5;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_C3 = CLBLL_L_X4Y157_SLICE_X4Y157_CO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_C4 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_C6 = CLBLM_R_X5Y156_SLICE_X7Y156_AQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D1 = CLBLM_R_X5Y146_SLICE_X6Y146_AQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D2 = CLBLM_R_X5Y146_SLICE_X6Y146_BQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D3 = CLBLM_R_X5Y144_SLICE_X6Y144_BQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D4 = CLBLM_R_X5Y146_SLICE_X6Y146_A5Q;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D5 = CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  assign CLBLM_R_X5Y144_SLICE_X6Y144_D6 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_D1 = CLBLM_R_X3Y153_SLICE_X2Y153_AO6;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_D2 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_D3 = CLBLM_R_X3Y151_SLICE_X2Y151_CO5;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_D4 = CLBLL_L_X2Y154_SLICE_X1Y154_AO5;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_D5 = CLBLL_L_X4Y155_SLICE_X4Y155_AQ;
  assign CLBLL_L_X2Y153_SLICE_X1Y153_D6 = CLBLM_R_X5Y156_SLICE_X7Y156_AQ;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_D1 = CLBLM_R_X13Y155_SLICE_X18Y155_CO5;
  assign RIOB33_X105Y153_IOB_X1Y154_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOB33_X105Y153_IOB_X1Y153_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y161_OLOGIC_X1Y161_T1 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_D2 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_D3 = 1'b1;
  assign LIOB33_X0Y185_IOB_X0Y186_O = RIOB33_X105Y143_IOB_X1Y143_I;
  assign LIOB33_X0Y185_IOB_X0Y185_O = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_A1 = CLBLM_L_X10Y154_SLICE_X12Y154_A5Q;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_A4 = CLBLL_L_X4Y158_SLICE_X4Y158_AO6;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_A5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_A1 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_A2 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_A3 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_A4 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_A5 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_A6 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_A6 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_AX = CLBLM_R_X7Y155_SLICE_X9Y155_CO5;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_B1 = CLBLM_R_X7Y155_SLICE_X8Y155_CO6;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_B1 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_B2 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_B3 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_B4 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_B5 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_B6 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_D4 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_B4 = CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_B6 = CLBLM_R_X5Y149_SLICE_X7Y149_CQ;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_C1 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_C2 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_C3 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_C4 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_C5 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_C6 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_C3 = CLBLM_L_X8Y156_SLICE_X11Y156_AQ;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_C4 = CLBLM_R_X7Y155_SLICE_X9Y155_A5Q;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_C5 = CLBLM_R_X7Y155_SLICE_X8Y155_CO6;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_C6 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_D1 = CLBLM_L_X8Y155_SLICE_X10Y155_AQ;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_D2 = CLBLM_L_X8Y156_SLICE_X10Y156_AQ;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_D1 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_D2 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_D3 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_D4 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_D5 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X0Y154_D6 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_D3 = CLBLM_R_X3Y153_SLICE_X3Y153_AO6;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_D4 = CLBLM_R_X3Y157_SLICE_X2Y157_AO5;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_A1 = CLBLM_R_X7Y158_SLICE_X8Y158_DO6;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_A2 = CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_A4 = CLBLM_L_X8Y154_SLICE_X11Y154_A5Q;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_A5 = CLBLL_L_X4Y153_SLICE_X4Y153_AO6;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_A6 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_B1 = CLBLM_R_X7Y156_SLICE_X8Y156_CQ;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_B2 = CLBLM_R_X7Y156_SLICE_X8Y156_BQ;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_B3 = CLBLM_R_X7Y158_SLICE_X8Y158_CO5;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_B4 = CLBLM_R_X7Y158_SLICE_X8Y158_BQ;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_B5 = CLBLM_R_X7Y152_SLICE_X8Y152_AQ;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_B6 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_C1 = CLBLM_R_X7Y152_SLICE_X8Y152_AQ;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_C2 = CLBLM_R_X7Y155_SLICE_X8Y155_AQ;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_C3 = CLBLM_R_X7Y158_SLICE_X8Y158_BQ;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_C4 = CLBLM_R_X7Y156_SLICE_X8Y156_CQ;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_C5 = CLBLM_L_X8Y154_SLICE_X10Y154_A5Q;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_A1 = CLBLL_L_X4Y157_SLICE_X4Y157_CO6;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_A2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_A6 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_C6 = CLBLM_R_X7Y156_SLICE_X8Y156_BQ;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_B1 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_B2 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_B3 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_B4 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_B5 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_B6 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_D1 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_D2 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_D3 = CLBLM_R_X7Y158_SLICE_X8Y158_BQ;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_C1 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_C2 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_C3 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_C4 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_C5 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_C6 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_C4 = CLBLM_L_X12Y154_SLICE_X17Y154_A5Q;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_C5 = CLBLM_R_X11Y158_SLICE_X15Y158_BO6;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_C6 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_D1 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_D2 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_D3 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_D4 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_D5 = 1'b1;
  assign CLBLL_L_X2Y154_SLICE_X1Y154_D6 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_D2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_D1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign LIOI3_X0Y175_OLOGIC_X0Y176_T1 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_D5 = CLBLM_L_X10Y148_SLICE_X12Y148_DO6;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_D1 = CLBLM_R_X11Y144_SLICE_X15Y144_AQ;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_D6 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_D1 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign LIOI3_X0Y115_OLOGIC_X0Y116_T1 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_D1 = CLBLM_R_X13Y155_SLICE_X18Y155_CO6;
  assign LIOI3_X0Y175_OLOGIC_X0Y175_T1 = 1'b1;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_D1 = CLBLM_L_X12Y151_SLICE_X16Y151_CQ;
  assign RIOI3_X105Y159_OLOGIC_X1Y160_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_D1 = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOI3_X0Y115_OLOGIC_X0Y115_T1 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_D1 = CLBLM_R_X13Y154_SLICE_X18Y154_DO6;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y188_T1 = 1'b1;
  assign RIOI3_X105Y159_OLOGIC_X1Y159_T1 = 1'b1;
  assign RIOB33_X105Y155_IOB_X1Y156_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOB33_X105Y155_IOB_X1Y155_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_D1 = RIOB33_X105Y143_IOB_X1Y144_I;
  assign LIOI3_TBYTETERM_X0Y187_OLOGIC_X0Y187_T1 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_D1 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_C4 = CLBLM_R_X7Y148_SLICE_X8Y148_AQ;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_C5 = CLBLM_L_X8Y158_SLICE_X10Y158_AQ;
  assign CLBLM_R_X11Y158_SLICE_X14Y158_D5 = CLBLM_L_X12Y158_SLICE_X17Y158_AQ;
  assign LIOB33_X0Y187_IOB_X0Y188_O = RIOB33_X105Y145_IOB_X1Y145_I;
  assign LIOB33_X0Y187_IOB_X0Y187_O = RIOB33_X105Y143_IOB_X1Y144_I;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_C6 = CLBLM_R_X7Y148_SLICE_X8Y148_BQ;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_B6 = CLBLM_L_X12Y154_SLICE_X16Y154_BQ;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_A1 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_A2 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_A3 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_A4 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_A5 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_A6 = 1'b1;
  assign CLBLM_R_X7Y156_SLICE_X9Y156_A1 = CLBLM_R_X5Y152_SLICE_X6Y152_CO5;
  assign CLBLM_R_X7Y156_SLICE_X9Y156_A2 = CLBLM_L_X10Y157_SLICE_X12Y157_AQ;
  assign CLBLM_R_X7Y156_SLICE_X9Y156_A3 = CLBLM_R_X7Y156_SLICE_X9Y156_AQ;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_B1 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_B2 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_B3 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_B4 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_B5 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_B6 = 1'b1;
  assign CLBLM_R_X7Y156_SLICE_X9Y156_B1 = 1'b1;
  assign CLBLM_R_X7Y156_SLICE_X9Y156_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_C1 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_C2 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_C3 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_C4 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_C5 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_C6 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_D2 = CLBLM_R_X13Y151_SLICE_X18Y151_CQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A1 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A2 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A3 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A4 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A5 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_A6 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_C4 = CLBLM_L_X8Y153_SLICE_X11Y153_BQ;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_D1 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_D2 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_D3 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_D4 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_D5 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X0Y155_D6 = 1'b1;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_D5 = CLBLM_R_X13Y155_SLICE_X18Y155_BQ;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y156_SLICE_X13Y156_D6 = CLBLM_R_X11Y154_SLICE_X14Y154_CQ;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_C6 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C1 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C2 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C3 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C4 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C5 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_C6 = 1'b1;
  assign CLBLM_R_X7Y156_SLICE_X8Y156_A1 = CLBLM_L_X10Y151_SLICE_X12Y151_CQ;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D1 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D2 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D3 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D4 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D5 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_D6 = 1'b1;
  assign CLBLM_R_X7Y156_SLICE_X8Y156_B4 = CLBLM_R_X7Y158_SLICE_X8Y158_BQ;
  assign CLBLM_R_X7Y156_SLICE_X8Y156_B5 = CLBLM_R_X7Y156_SLICE_X9Y156_AQ;
  assign CLBLM_R_X7Y156_SLICE_X8Y156_B6 = CLBLM_R_X7Y155_SLICE_X8Y155_BO6;
  assign CLBLM_R_X7Y156_SLICE_X8Y156_B1 = CLBLM_R_X7Y156_SLICE_X8Y156_CQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A1 = CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A2 = CLBLM_R_X5Y147_SLICE_X6Y147_BQ;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_A1 = CLBLM_R_X3Y158_SLICE_X2Y158_AO6;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_A3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_A4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_A5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_A6 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A3 = CLBLM_R_X5Y146_SLICE_X6Y146_AQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A5 = CLBLM_R_X5Y146_SLICE_X6Y146_CO5;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_B1 = CLBLM_R_X3Y158_SLICE_X2Y158_AO6;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_B2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_B3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_B4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_B5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_B6 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_AX = CLBLM_R_X5Y146_SLICE_X6Y146_CO6;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B2 = CLBLM_R_X5Y146_SLICE_X6Y146_BQ;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_C1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_C2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_C3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_C4 = 1'b1;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_C5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_C6 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C1 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C3 = CLBLM_R_X7Y152_SLICE_X8Y152_AQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C4 = CLBLM_R_X5Y146_SLICE_X6Y146_A5Q;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_C6 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_D1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_D2 = CLBLM_R_X3Y155_SLICE_X2Y155_DO6;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_D3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_D4 = CLBLM_R_X3Y158_SLICE_X2Y158_AO6;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_D5 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLL_L_X2Y155_SLICE_X1Y155_D6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D1 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D2 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D3 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D4 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D5 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y70_D = LIOB33_X0Y69_IOB_X0Y70_I;
  assign LIOI3_TBYTESRC_X0Y69_ILOGIC_X0Y69_D = LIOB33_X0Y69_IOB_X0Y69_I;
  assign RIOB33_SING_X105Y199_IOB_X1Y199_O = CLBLM_R_X13Y156_SLICE_X19Y156_AQ;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_B5 = CLBLM_L_X10Y156_SLICE_X12Y156_CO6;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_B6 = CLBLM_L_X10Y155_SLICE_X12Y155_CQ;
  assign CLBLM_L_X12Y157_SLICE_X16Y157_D2 = CLBLM_R_X11Y158_SLICE_X14Y158_BQ;
  assign RIOB33_X105Y157_IOB_X1Y158_O = CLBLL_L_X36Y150_SLICE_X54Y150_AO6;
  assign RIOB33_X105Y157_IOB_X1Y157_O = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_C4 = CLBLM_L_X12Y158_SLICE_X16Y158_A5Q;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B1 = CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_C5 = CLBLM_L_X10Y153_SLICE_X13Y153_DQ;
  assign CLBLM_L_X12Y157_SLICE_X16Y157_D3 = CLBLM_R_X11Y157_SLICE_X14Y157_CQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B2 = CLBLM_R_X11Y152_SLICE_X15Y152_BQ;
  assign CLBLM_L_X10Y156_SLICE_X12Y156_C6 = CLBLM_L_X8Y155_SLICE_X11Y155_BQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y157_SLICE_X16Y157_D4 = CLBLM_R_X11Y159_SLICE_X15Y159_DO5;
  assign LIOB33_X0Y189_IOB_X0Y190_O = RIOB33_X105Y147_IOB_X1Y147_I;
  assign LIOB33_X0Y189_IOB_X0Y189_O = RIOB33_X105Y145_IOB_X1Y146_I;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C1 = CLBLM_L_X12Y153_SLICE_X17Y153_BQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C2 = CLBLM_R_X11Y152_SLICE_X15Y152_CQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C5 = CLBLM_R_X11Y154_SLICE_X14Y154_DQ;
  assign CLBLM_R_X11Y152_SLICE_X15Y152_C6 = CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_A1 = CLBLM_R_X7Y158_SLICE_X8Y158_CO5;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_A2 = CLBLM_R_X7Y155_SLICE_X9Y155_BQ;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_A3 = CLBLM_R_X7Y157_SLICE_X9Y157_AQ;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_A5 = CLBLL_L_X4Y155_SLICE_X4Y155_BQ;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_A6 = CLBLM_R_X7Y155_SLICE_X8Y155_CO6;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_B1 = CLBLM_R_X5Y157_SLICE_X7Y157_DQ;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_B2 = CLBLM_R_X7Y157_SLICE_X9Y157_BQ;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_B4 = CLBLM_R_X5Y152_SLICE_X6Y152_CO5;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_B5 = CLBLM_L_X12Y156_SLICE_X16Y156_BQ;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_B6 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A1 = CLBLM_R_X5Y152_SLICE_X6Y152_CO6;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A2 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A3 = CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A5 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_A6 = CLBLM_R_X5Y148_SLICE_X6Y148_A5Q;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_C2 = CLBLM_R_X7Y157_SLICE_X9Y157_CQ;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_C3 = CLBLM_R_X7Y152_SLICE_X8Y152_A5Q;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B1 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B3 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B5 = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_B6 = CLBLM_L_X10Y150_SLICE_X12Y150_CO6;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C1 = CLBLM_R_X5Y148_SLICE_X7Y148_AQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C2 = CLBLM_R_X5Y147_SLICE_X7Y147_CQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C3 = CLBLM_R_X7Y148_SLICE_X8Y148_CQ;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C5 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_C6 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_D3 = CLBLM_R_X7Y157_SLICE_X9Y157_DQ;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_A1 = CLBLM_R_X7Y159_SLICE_X8Y159_BO5;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_A2 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_A4 = CLBLM_R_X7Y158_SLICE_X8Y158_BQ;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_A5 = CLBLM_L_X8Y156_SLICE_X11Y156_B5Q;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D1 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D2 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D3 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D4 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D5 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X7Y147_D6 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_A6 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_B1 = CLBLM_R_X7Y159_SLICE_X8Y159_BO5;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_B2 = CLBLM_L_X10Y145_SLICE_X12Y145_CQ;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_B3 = CLBLM_R_X7Y157_SLICE_X8Y157_AQ;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_B4 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A1 = CLBLM_R_X7Y152_SLICE_X8Y152_BO5;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A2 = CLBLM_R_X5Y149_SLICE_X6Y149_AQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A3 = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A4 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_A6 = CLBLL_L_X4Y146_SLICE_X5Y146_AO5;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_C1 = CLBLM_R_X11Y155_SLICE_X14Y155_AQ;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_C3 = CLBLM_R_X7Y157_SLICE_X8Y157_BQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B1 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B2 = CLBLM_R_X5Y147_SLICE_X6Y147_BQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B3 = CLBLL_L_X4Y147_SLICE_X4Y147_BO6;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B5 = CLBLM_L_X8Y155_SLICE_X11Y155_BQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_B6 = CLBLM_R_X5Y148_SLICE_X7Y148_A5Q;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_B4 = CLBLM_R_X5Y152_SLICE_X7Y152_CQ;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_D1 = CLBLM_L_X8Y157_SLICE_X11Y157_BQ;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C1 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C2 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C3 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C4 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C5 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_C6 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_B5 = CLBLM_R_X5Y152_SLICE_X6Y152_CO5;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_B6 = CLBLM_L_X8Y154_SLICE_X10Y154_B5Q;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_D4 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_D6 = CLBLM_R_X5Y152_SLICE_X6Y152_CO5;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D1 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D2 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D3 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D4 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D5 = 1'b1;
  assign CLBLM_R_X5Y147_SLICE_X6Y147_D6 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_C2 = CLBLL_L_X4Y150_SLICE_X4Y150_CQ;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_C3 = CLBLM_L_X8Y153_SLICE_X10Y153_CO6;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_C5 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_C6 = CLBLM_L_X10Y154_SLICE_X12Y154_AQ;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOB33_X0Y183_IOB_X0Y184_O = RIOB33_X105Y135_IOB_X1Y136_I;
  assign LIOB33_X0Y183_IOB_X0Y183_O = RIOB33_X105Y135_IOB_X1Y135_I;
  assign RIOB33_X105Y159_IOB_X1Y160_O = CLBLM_R_X13Y155_SLICE_X18Y155_CO6;
  assign RIOB33_X105Y159_IOB_X1Y159_O = CLBLM_R_X13Y154_SLICE_X18Y154_DO6;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_D1 = CLBLM_R_X3Y155_SLICE_X3Y155_AO6;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_D2 = CLBLM_R_X13Y155_SLICE_X19Y155_AO6;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_D3 = CLBLM_R_X7Y148_SLICE_X9Y148_BQ;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_D4 = CLBLM_R_X7Y155_SLICE_X9Y155_DO6;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_D5 = CLBLM_R_X5Y156_SLICE_X6Y156_AO6;
  assign LIOB33_X0Y191_IOB_X0Y192_O = LIOB33_X0Y51_IOB_X0Y52_I;
  assign LIOB33_X0Y191_IOB_X0Y191_O = RIOB33_X105Y147_IOB_X1Y148_I;
  assign CLBLM_R_X7Y154_SLICE_X9Y154_D6 = CLBLM_R_X13Y154_SLICE_X19Y154_AQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A2 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_A5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_A1 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_A2 = CLBLM_R_X7Y154_SLICE_X8Y154_DO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_AX = CLBLM_L_X10Y148_SLICE_X12Y148_BO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_D1 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y177_OLOGIC_X0Y178_T1 = 1'b1;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_B4 = CLBLM_R_X5Y155_SLICE_X7Y155_DO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B2 = CLBLM_L_X8Y148_SLICE_X11Y148_A5Q;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_D1 = CLBLM_R_X5Y148_SLICE_X7Y148_BQ;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_B5 = CLBLM_R_X5Y157_SLICE_X6Y157_DO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B3 = CLBLM_R_X7Y148_SLICE_X9Y148_AQ;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_D1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B4 = 1'b1;
  assign CLBLM_R_X11Y152_SLICE_X14Y152_D6 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_T1 = 1'b1;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B5 = CLBLL_L_X4Y151_SLICE_X5Y151_CQ;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_D1 = CLBLM_L_X12Y155_SLICE_X17Y155_DO6;
  assign CLBLM_L_X8Y148_SLICE_X11Y148_B6 = 1'b1;
  assign LIOI3_X0Y177_OLOGIC_X0Y177_T1 = 1'b1;
  assign CLBLM_R_X7Y158_SLICE_X9Y158_A1 = CLBLM_L_X8Y154_SLICE_X10Y154_A5Q;
  assign CLBLM_R_X7Y158_SLICE_X9Y158_A2 = CLBLM_R_X5Y152_SLICE_X6Y152_CO5;
  assign CLBLM_R_X7Y158_SLICE_X9Y158_A3 = CLBLM_R_X7Y158_SLICE_X9Y158_AQ;
  assign CLBLM_R_X7Y158_SLICE_X9Y158_A4 = 1'b1;
  assign CLBLM_R_X7Y158_SLICE_X9Y158_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y158_SLICE_X9Y158_A6 = CLBLM_R_X7Y154_SLICE_X9Y154_CQ;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_D1 = CLBLM_R_X5Y147_SLICE_X7Y147_CQ;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_D1 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign RIOI3_X105Y161_OLOGIC_X1Y162_T1 = 1'b1;
  assign CLBLM_R_X7Y158_SLICE_X9Y158_B1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X7Y158_SLICE_X9Y158_B2 = CLBLM_R_X13Y150_SLICE_X18Y150_AQ;
  assign CLBLM_R_X7Y158_SLICE_X9Y158_B3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X7Y158_SLICE_X9Y158_B4 = CLBLL_L_X4Y157_SLICE_X4Y157_CO5;
  assign CLBLM_R_X7Y158_SLICE_X9Y158_B5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y158_SLICE_X9Y158_B6 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOI3_X0Y117_OLOGIC_X0Y117_T1 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_B4 = CLBLM_R_X7Y158_SLICE_X8Y158_CO5;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A2 = CLBLM_L_X8Y148_SLICE_X10Y148_BQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A3 = CLBLM_R_X5Y148_SLICE_X7Y148_AQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A4 = CLBLM_R_X7Y147_SLICE_X9Y147_BQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A5 = CLBLM_L_X10Y151_SLICE_X12Y151_CQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_A6 = CLBLL_L_X4Y151_SLICE_X4Y151_BQ;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_B5 = CLBLM_R_X5Y154_SLICE_X6Y154_AQ;
  assign CLBLM_R_X7Y158_SLICE_X9Y158_C1 = CLBLM_L_X10Y158_SLICE_X12Y158_AQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_AX = CLBLM_R_X5Y149_SLICE_X7Y149_DO5;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B1 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B2 = CLBLM_L_X8Y148_SLICE_X10Y148_AQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B5 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_B6 = 1'b1;
  assign CLBLM_R_X7Y158_SLICE_X9Y158_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_C6 = CLBLL_L_X4Y151_SLICE_X5Y151_DO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C1 = CLBLM_R_X5Y149_SLICE_X7Y149_AQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C2 = CLBLM_L_X8Y148_SLICE_X10Y148_AQ;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C5 = CLBLM_R_X5Y148_SLICE_X7Y148_DO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_C6 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X7Y158_SLICE_X9Y158_D3 = CLBLM_R_X7Y158_SLICE_X9Y158_BO6;
  assign CLBLM_R_X7Y158_SLICE_X9Y158_D4 = CLBLM_R_X7Y158_SLICE_X9Y158_CO6;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y158_SLICE_X8Y158_A1 = 1'b1;
  assign CLBLM_R_X7Y158_SLICE_X8Y158_A2 = CLBLM_R_X7Y156_SLICE_X8Y156_AQ;
  assign CLBLM_R_X7Y158_SLICE_X8Y158_A3 = CLBLM_R_X7Y158_SLICE_X8Y158_AQ;
  assign CLBLL_L_X4Y154_SLICE_X5Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y158_SLICE_X8Y158_A4 = CLBLM_R_X5Y152_SLICE_X6Y152_CO5;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D2 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D4 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X5Y148_SLICE_X7Y148_D6 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X7Y158_SLICE_X8Y158_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y158_SLICE_X8Y158_A6 = CLBLM_L_X8Y153_SLICE_X11Y153_DQ;
  assign CLBLM_R_X7Y158_SLICE_X8Y158_B1 = CLBLM_R_X7Y159_SLICE_X8Y159_BO5;
  assign CLBLM_R_X7Y158_SLICE_X8Y158_B2 = CLBLL_L_X4Y155_SLICE_X5Y155_BQ;
  assign CLBLM_R_X7Y158_SLICE_X8Y158_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A1 = CLBLM_R_X5Y148_SLICE_X6Y148_AQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A3 = CLBLM_L_X10Y149_SLICE_X12Y149_DO5;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A4 = CLBLM_L_X10Y149_SLICE_X12Y149_CQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A5 = CLBLM_R_X5Y148_SLICE_X6Y148_CO5;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_A6 = CLBLM_R_X5Y148_SLICE_X6Y148_BQ;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_C4 = CLBLL_L_X4Y151_SLICE_X4Y151_CQ;
  assign CLBLM_R_X7Y158_SLICE_X8Y158_C3 = CLBLM_L_X8Y154_SLICE_X10Y154_A5Q;
  assign CLBLM_R_X7Y158_SLICE_X8Y158_C4 = CLBLM_R_X7Y155_SLICE_X8Y155_BO5;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_AX = CLBLM_L_X8Y148_SLICE_X11Y148_DO5;
  assign CLBLM_R_X7Y158_SLICE_X8Y158_C5 = CLBLM_L_X8Y158_SLICE_X10Y158_AQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B1 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B3 = CLBLM_L_X10Y149_SLICE_X12Y149_DO5;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B4 = CLBLM_R_X5Y158_SLICE_X6Y158_BQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B5 = CLBLM_R_X5Y148_SLICE_X6Y148_CO5;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_B6 = CLBLM_R_X5Y148_SLICE_X6Y148_BQ;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_C5 = CLBLM_L_X8Y154_SLICE_X10Y154_A5Q;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_C6 = CLBLM_L_X8Y158_SLICE_X10Y158_AQ;
  assign CLBLM_R_X7Y158_SLICE_X8Y158_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C1 = CLBLM_R_X7Y148_SLICE_X8Y148_CQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C2 = CLBLM_R_X7Y148_SLICE_X8Y148_A5Q;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C3 = CLBLM_L_X10Y149_SLICE_X12Y149_BQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C4 = CLBLL_L_X4Y148_SLICE_X5Y148_DQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C5 = CLBLM_R_X5Y148_SLICE_X6Y148_DO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_C6 = 1'b1;
  assign CLBLM_R_X7Y158_SLICE_X8Y158_D2 = CLBLM_R_X7Y155_SLICE_X8Y155_CO6;
  assign CLBLM_R_X7Y158_SLICE_X8Y158_D3 = CLBLM_R_X7Y155_SLICE_X8Y155_AQ;
  assign CLBLM_R_X7Y158_SLICE_X8Y158_D4 = CLBLM_R_X7Y158_SLICE_X8Y158_CO6;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y158_SLICE_X8Y158_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D1 = 1'b1;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D2 = CLBLL_L_X4Y150_SLICE_X5Y150_BQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D3 = CLBLM_R_X5Y148_SLICE_X6Y148_AQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D4 = CLBLM_R_X5Y148_SLICE_X6Y148_BQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D5 = CLBLM_R_X5Y149_SLICE_X7Y149_CQ;
  assign CLBLM_R_X5Y148_SLICE_X6Y148_D6 = CLBLL_L_X4Y150_SLICE_X5Y150_AQ;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_D1 = LIOB33_X0Y71_IOB_X0Y71_I;
  assign RIOB33_X105Y161_IOB_X1Y162_O = CLBLM_L_X12Y155_SLICE_X17Y155_DO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_D1 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign RIOB33_X105Y161_IOB_X1Y161_O = CLBLM_R_X13Y155_SLICE_X18Y155_CO5;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_D3 = 1'b1;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_D4 = CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_D5 = CLBLL_L_X4Y153_SLICE_X4Y153_AO6;
  assign CLBLM_R_X7Y154_SLICE_X8Y154_D6 = CLBLM_R_X7Y154_SLICE_X8Y154_AQ;
  assign LIOB33_X0Y193_IOB_X0Y194_O = LIOB33_X0Y59_IOB_X0Y60_I;
  assign LIOB33_X0Y193_IOB_X0Y193_O = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_T1 = 1'b1;
  assign LIOI3_X0Y55_ILOGIC_X0Y56_D = LIOB33_X0Y55_IOB_X0Y56_I;
  assign LIOI3_X0Y55_ILOGIC_X0Y55_D = LIOB33_X0Y55_IOB_X0Y55_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_D = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_D = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A1 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X9Y144_A2 = 1'b1;
  assign RIOI3_X105Y151_OLOGIC_X1Y152_T1 = 1'b1;
  assign CLBLM_R_X7Y159_SLICE_X9Y159_A1 = CLBLM_R_X7Y159_SLICE_X9Y159_BO6;
  assign CLBLM_R_X7Y159_SLICE_X9Y159_A2 = CLBLM_R_X7Y148_SLICE_X8Y148_AQ;
  assign CLBLM_R_X7Y159_SLICE_X9Y159_A3 = CLBLM_L_X8Y159_SLICE_X10Y159_AQ;
  assign CLBLM_R_X7Y159_SLICE_X9Y159_A4 = CLBLM_L_X8Y158_SLICE_X10Y158_AQ;
  assign CLBLM_R_X7Y159_SLICE_X9Y159_A5 = CLBLM_R_X7Y148_SLICE_X8Y148_BQ;
  assign CLBLM_R_X7Y159_SLICE_X9Y159_A6 = CLBLM_R_X7Y159_SLICE_X9Y159_CO6;
  assign CLBLM_R_X7Y159_SLICE_X9Y159_B1 = CLBLM_L_X8Y154_SLICE_X10Y154_A5Q;
  assign CLBLM_R_X7Y159_SLICE_X9Y159_B2 = CLBLM_R_X7Y148_SLICE_X8Y148_AQ;
  assign CLBLM_R_X7Y159_SLICE_X9Y159_B3 = CLBLM_R_X7Y155_SLICE_X8Y155_AQ;
  assign CLBLM_R_X7Y159_SLICE_X9Y159_B4 = CLBLM_R_X7Y148_SLICE_X8Y148_BQ;
  assign CLBLM_R_X7Y159_SLICE_X9Y159_B5 = CLBLM_L_X8Y158_SLICE_X10Y158_AQ;
  assign CLBLM_R_X7Y159_SLICE_X9Y159_B6 = CLBLM_R_X7Y157_SLICE_X8Y157_CQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A2 = CLBLL_L_X4Y153_SLICE_X4Y153_AO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A3 = CLBLM_R_X5Y149_SLICE_X6Y149_CO5;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A4 = CLBLM_R_X7Y148_SLICE_X8Y148_BQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A5 = CLBLM_R_X5Y149_SLICE_X7Y149_AQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y159_SLICE_X9Y159_C1 = CLBLM_R_X7Y148_SLICE_X8Y148_AQ;
  assign CLBLM_R_X7Y159_SLICE_X9Y159_C2 = CLBLM_R_X7Y148_SLICE_X8Y148_BQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_AX = CLBLM_R_X5Y149_SLICE_X6Y149_CO6;
  assign CLBLM_R_X7Y159_SLICE_X9Y159_C3 = CLBLM_L_X8Y150_SLICE_X11Y150_CQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B1 = CLBLM_L_X8Y151_SLICE_X10Y151_CQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B2 = CLBLM_R_X5Y149_SLICE_X7Y149_BQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B3 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B4 = CLBLM_R_X5Y152_SLICE_X6Y152_CO6;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_B6 = CLBLM_L_X12Y149_SLICE_X16Y149_BQ;
  assign CLBLM_R_X7Y159_SLICE_X9Y159_D1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X7Y159_SLICE_X9Y159_D2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C2 = CLBLM_R_X5Y149_SLICE_X7Y149_CQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C3 = CLBLM_L_X8Y155_SLICE_X10Y155_B5Q;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C4 = CLBLL_L_X4Y149_SLICE_X5Y149_BO5;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C5 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_C6 = CLBLM_L_X10Y149_SLICE_X12Y149_DO5;
  assign CLBLM_R_X7Y159_SLICE_X9Y159_D3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X7Y159_SLICE_X9Y159_D4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y159_SLICE_X8Y159_A1 = CLBLM_R_X7Y159_SLICE_X8Y159_BO5;
  assign CLBLM_R_X7Y159_SLICE_X8Y159_A2 = CLBLM_R_X11Y158_SLICE_X15Y158_AQ;
  assign CLBLM_R_X7Y159_SLICE_X8Y159_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y159_SLICE_X8Y159_A4 = 1'b1;
  assign CLBLM_R_X7Y159_SLICE_X8Y159_A5 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D2 = CLBLM_R_X11Y149_SLICE_X15Y149_A5Q;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D3 = CLBLL_L_X4Y150_SLICE_X5Y150_BQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D4 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D5 = CLBLM_L_X8Y151_SLICE_X10Y151_AQ;
  assign CLBLM_R_X5Y149_SLICE_X7Y149_D6 = 1'b1;
  assign CLBLM_R_X7Y159_SLICE_X8Y159_A6 = CLBLM_R_X7Y157_SLICE_X8Y157_CQ;
  assign CLBLM_R_X7Y159_SLICE_X8Y159_B1 = CLBLM_L_X8Y154_SLICE_X10Y154_A5Q;
  assign CLBLM_R_X7Y159_SLICE_X8Y159_B2 = CLBLM_L_X8Y158_SLICE_X10Y158_AQ;
  assign CLBLM_R_X7Y159_SLICE_X8Y159_B3 = CLBLM_L_X10Y159_SLICE_X12Y159_AO6;
  assign CLBLM_R_X7Y159_SLICE_X8Y159_B4 = CLBLM_R_X7Y148_SLICE_X8Y148_BQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A2 = CLBLM_R_X5Y150_SLICE_X6Y150_BQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A3 = CLBLL_L_X4Y148_SLICE_X4Y148_AQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A4 = CLBLM_R_X5Y147_SLICE_X7Y147_BQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A5 = CLBLM_R_X5Y148_SLICE_X6Y148_BQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_A6 = 1'b1;
  assign CLBLM_R_X7Y159_SLICE_X8Y159_C1 = 1'b1;
  assign CLBLM_R_X7Y159_SLICE_X8Y159_C2 = 1'b1;
  assign CLBLM_R_X7Y159_SLICE_X8Y159_C3 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B1 = CLBLM_R_X7Y151_SLICE_X9Y151_BQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B3 = CLBLM_L_X8Y147_SLICE_X11Y147_BQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B4 = CLBLM_L_X8Y147_SLICE_X11Y147_CO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B5 = CLBLL_L_X4Y153_SLICE_X4Y153_BO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_B6 = 1'b1;
  assign CLBLM_R_X7Y159_SLICE_X8Y159_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y159_SLICE_X8Y159_D1 = 1'b1;
  assign CLBLM_R_X7Y159_SLICE_X8Y159_D2 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C2 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C3 = CLBLM_L_X10Y149_SLICE_X13Y149_A5Q;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C5 = CLBLM_R_X7Y149_SLICE_X8Y149_DO6;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_C6 = 1'b1;
  assign CLBLM_R_X7Y159_SLICE_X8Y159_D3 = 1'b1;
  assign CLBLM_R_X7Y159_SLICE_X8Y159_D4 = 1'b1;
  assign CLBLM_R_X7Y159_SLICE_X8Y159_D5 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X7Y159_SLICE_X8Y159_D6 = 1'b1;
  assign CLBLM_R_X13Y157_SLICE_X19Y157_C4 = 1'b1;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D1 = CLBLM_R_X5Y148_SLICE_X6Y148_BQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D2 = CLBLM_R_X7Y148_SLICE_X8Y148_A5Q;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D3 = CLBLM_R_X5Y148_SLICE_X6Y148_AQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D4 = CLBLL_L_X4Y148_SLICE_X5Y148_DQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D5 = CLBLM_L_X10Y149_SLICE_X12Y149_BQ;
  assign CLBLM_R_X5Y149_SLICE_X6Y149_D6 = CLBLM_R_X7Y148_SLICE_X8Y148_CQ;
  assign RIOB33_X105Y163_IOB_X1Y163_O = CLBLM_L_X12Y155_SLICE_X17Y155_DO5;
  assign RIOB33_X105Y163_IOB_X1Y164_O = CLBLM_R_X7Y149_SLICE_X9Y149_DO5;
  assign CLBLM_R_X13Y157_SLICE_X19Y157_C5 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B1 = 1'b1;
  assign CLBLM_R_X13Y157_SLICE_X19Y157_C6 = 1'b1;
  assign LIOB33_X0Y195_IOB_X0Y196_O = LIOB33_X0Y69_IOB_X0Y69_I;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B2 = 1'b1;
  assign LIOB33_X0Y195_IOB_X0Y195_O = LIOB33_X0Y63_IOB_X0Y64_I;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B3 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B4 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B5 = 1'b1;
  assign CLBLM_R_X5Y146_SLICE_X7Y146_B6 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOB33_X0Y161_IOB_X0Y162_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign LIOB33_X0Y161_IOB_X0Y161_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X13Y159_SLICE_X18Y159_A2 = CLBLM_R_X13Y158_SLICE_X18Y158_BQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B3 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B4 = 1'b1;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B5 = CLBLM_R_X5Y146_SLICE_X6Y146_AQ;
  assign CLBLM_R_X7Y144_SLICE_X8Y144_B6 = CLBLM_R_X5Y146_SLICE_X6Y146_A5Q;
  assign CLBLM_R_X13Y159_SLICE_X18Y159_A3 = CLBLM_R_X11Y158_SLICE_X14Y158_AQ;
  assign CLBLM_R_X13Y159_SLICE_X18Y159_A4 = CLBLM_R_X11Y157_SLICE_X15Y157_BQ;
  assign CLBLM_R_X13Y159_SLICE_X18Y159_A5 = CLBLM_R_X13Y157_SLICE_X19Y157_AQ;
  assign CLBLM_R_X13Y159_SLICE_X18Y159_A6 = CLBLM_R_X13Y159_SLICE_X18Y159_CO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A1 = CLBLM_R_X5Y156_SLICE_X7Y156_AQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A2 = CLBLL_L_X4Y150_SLICE_X5Y150_AQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A3 = CLBLM_R_X5Y150_SLICE_X7Y150_AQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_A6 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B1 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B2 = CLBLM_R_X7Y150_SLICE_X8Y150_BQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B4 = CLBLL_L_X4Y149_SLICE_X4Y149_BQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B5 = CLBLM_R_X7Y150_SLICE_X9Y150_AO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C1 = CLBLM_R_X5Y151_SLICE_X6Y151_C5Q;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C2 = CLBLM_R_X5Y150_SLICE_X7Y150_CQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C3 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C4 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C5 = CLBLL_L_X4Y147_SLICE_X4Y147_BO6;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_A6 = CLBLM_R_X5Y146_SLICE_X6Y146_A5Q;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D1 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D2 = CLBLM_R_X5Y148_SLICE_X6Y148_A5Q;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D3 = CLBLM_L_X8Y151_SLICE_X10Y151_CQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D4 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D5 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X7Y150_D6 = CLBLM_L_X10Y150_SLICE_X12Y150_CQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A1 = CLBLM_R_X5Y150_SLICE_X7Y150_BQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A3 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A5 = CLBLM_R_X5Y149_SLICE_X6Y149_A5Q;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_A6 = CLBLM_R_X7Y150_SLICE_X9Y150_AO5;
  assign LIOI3_X0Y179_OLOGIC_X0Y180_D1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign RIOB33_X105Y165_IOB_X1Y165_O = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B1 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B2 = CLBLM_R_X5Y150_SLICE_X6Y150_BQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B3 = CLBLM_L_X12Y155_SLICE_X16Y155_CO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B5 = CLBLM_L_X10Y150_SLICE_X12Y150_A5Q;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_B6 = CLBLM_L_X8Y149_SLICE_X10Y149_AQ;
  assign RIOB33_X105Y165_IOB_X1Y166_O = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X13Y157_SLICE_X19Y157_D1 = 1'b1;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C1 = CLBLM_L_X10Y150_SLICE_X12Y150_A5Q;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C2 = CLBLM_R_X5Y150_SLICE_X6Y150_CQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C3 = CLBLM_L_X8Y148_SLICE_X10Y148_BQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C4 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B3 = CLBLM_R_X5Y144_SLICE_X6Y144_CO6;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_C6 = CLBLM_L_X12Y155_SLICE_X16Y155_CO6;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = CLBLL_L_X4Y149_SLICE_X5Y149_A5Q;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_D1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B5 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D1 = CLBLM_L_X10Y150_SLICE_X12Y150_A5Q;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D2 = CLBLM_L_X8Y148_SLICE_X10Y148_BQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D3 = CLBLM_R_X5Y150_SLICE_X6Y150_DQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D4 = CLBLM_L_X8Y148_SLICE_X11Y148_BQ;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y150_SLICE_X6Y150_D6 = CLBLM_L_X12Y155_SLICE_X16Y155_CO6;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_C4 = CLBLM_L_X8Y156_SLICE_X10Y156_BQ;
  assign CLBLM_R_X5Y146_SLICE_X6Y146_B6 = CLBLM_L_X10Y149_SLICE_X13Y149_BQ;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_C5 = CLBLM_L_X12Y150_SLICE_X17Y150_CO6;
  assign CLBLM_R_X13Y157_SLICE_X19Y157_D2 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = CLBLM_R_X11Y144_SLICE_X15Y144_A5Q;
  assign LIOI3_X0Y179_OLOGIC_X0Y179_T1 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_T1 = 1'b1;
  assign LIOB33_X0Y197_IOB_X0Y198_O = LIOB33_X0Y73_IOB_X0Y73_I;
  assign LIOB33_X0Y197_IOB_X0Y197_O = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_D1 = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLM_R_X13Y157_SLICE_X19Y157_D3 = 1'b1;
  assign RIOI3_X105Y165_OLOGIC_X1Y165_T1 = 1'b1;
  assign CLBLM_R_X13Y159_SLICE_X18Y159_B1 = CLBLM_R_X13Y159_SLICE_X18Y159_DO6;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_D2 = CLBLM_R_X11Y155_SLICE_X14Y155_DQ;
  assign CLBLM_R_X13Y159_SLICE_X18Y159_B2 = CLBLM_R_X11Y157_SLICE_X15Y157_BQ;
  assign CLBLM_L_X10Y157_SLICE_X13Y157_A5 = CLBLM_L_X12Y157_SLICE_X16Y157_CQ;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_D5 = CLBLM_L_X10Y150_SLICE_X13Y150_BQ;
  assign CLBLM_L_X10Y157_SLICE_X13Y157_A6 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_D6 = 1'b1;
  assign CLBLM_R_X13Y159_SLICE_X18Y159_B3 = CLBLM_R_X11Y158_SLICE_X14Y158_AQ;
  assign CLBLM_L_X10Y157_SLICE_X13Y157_B2 = CLBLM_R_X7Y157_SLICE_X9Y157_AQ;
  assign CLBLM_L_X10Y157_SLICE_X13Y157_B3 = CLBLM_L_X10Y159_SLICE_X12Y159_DO6;
  assign CLBLM_L_X10Y157_SLICE_X13Y157_B4 = CLBLM_L_X10Y157_SLICE_X12Y157_BQ;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_A1 = CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  assign CLBLM_R_X13Y159_SLICE_X18Y159_B4 = CLBLM_R_X13Y158_SLICE_X18Y158_BQ;
  assign CLBLM_L_X10Y157_SLICE_X13Y157_B5 = CLBLM_L_X10Y157_SLICE_X13Y157_AO6;
  assign CLBLM_L_X10Y157_SLICE_X13Y157_B6 = CLBLM_L_X8Y156_SLICE_X11Y156_DO6;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_D1 = CLBLM_R_X13Y153_SLICE_X19Y153_BQ;
  assign CLBLM_L_X10Y157_SLICE_X13Y157_C1 = CLBLM_R_X11Y156_SLICE_X14Y156_BQ;
  assign CLBLM_L_X10Y157_SLICE_X13Y157_C2 = CLBLM_L_X10Y155_SLICE_X12Y155_AQ;
  assign CLBLM_L_X10Y157_SLICE_X13Y157_C3 = CLBLM_L_X8Y157_SLICE_X11Y157_DO6;
  assign CLBLM_L_X10Y157_SLICE_X13Y157_C4 = CLBLM_L_X8Y156_SLICE_X11Y156_DO6;
  assign CLBLM_L_X10Y157_SLICE_X13Y157_C5 = CLBLM_L_X10Y157_SLICE_X13Y157_DO6;
  assign CLBLM_L_X10Y157_SLICE_X13Y157_C6 = CLBLM_L_X10Y156_SLICE_X13Y156_CO6;
  assign LIOI3_X0Y59_ILOGIC_X0Y60_D = LIOB33_X0Y59_IOB_X0Y60_I;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_B6 = 1'b1;
  assign LIOI3_X0Y59_ILOGIC_X0Y59_D = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOB33_X0Y79_IOB_X0Y80_O = CLBLL_L_X2Y140_SLICE_X0Y140_AO6;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_D = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_D = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A1 = CLBLM_R_X3Y152_SLICE_X3Y152_BO5;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A3 = CLBLM_R_X5Y151_SLICE_X7Y151_AQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A5 = CLBLL_L_X4Y151_SLICE_X4Y151_BQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_A6 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X10Y157_SLICE_X13Y157_D1 = CLBLM_R_X7Y148_SLICE_X8Y148_AQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B2 = CLBLM_R_X5Y151_SLICE_X7Y151_BQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B3 = CLBLM_R_X5Y149_SLICE_X6Y149_CO5;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B4 = CLBLM_L_X12Y154_SLICE_X16Y154_BQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_B6 = CLBLM_R_X3Y156_SLICE_X2Y156_DO6;
  assign CLBLM_L_X10Y157_SLICE_X13Y157_D2 = CLBLM_R_X7Y148_SLICE_X8Y148_BQ;
  assign CLBLM_L_X10Y157_SLICE_X13Y157_D3 = CLBLM_L_X8Y158_SLICE_X10Y158_AQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C2 = CLBLM_R_X5Y151_SLICE_X7Y151_CQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C4 = CLBLM_L_X8Y151_SLICE_X10Y151_CQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C5 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_C6 = 1'b1;
  assign CLBLM_L_X10Y157_SLICE_X13Y157_D4 = CLBLM_L_X12Y157_SLICE_X16Y157_CQ;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_C4 = CLBLM_L_X12Y154_SLICE_X16Y154_AQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y157_SLICE_X13Y157_D5 = CLBLM_R_X11Y156_SLICE_X15Y156_AQ;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_C5 = CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  assign RIOB33_X105Y167_IOB_X1Y167_O = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign RIOB33_X105Y167_IOB_X1Y168_O = CLBLM_L_X10Y163_SLICE_X13Y163_AO6;
  assign CLBLM_L_X10Y157_SLICE_X13Y157_D6 = CLBLM_L_X10Y157_SLICE_X12Y157_BQ;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_C6 = CLBLM_L_X12Y152_SLICE_X16Y152_DO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D3 = CLBLM_R_X5Y151_SLICE_X7Y151_DQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D4 = CLBLL_L_X4Y154_SLICE_X5Y154_BO6;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D5 = CLBLM_R_X5Y150_SLICE_X7Y150_BQ;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y151_SLICE_X7Y151_D2 = CLBLM_R_X5Y149_SLICE_X6Y149_CO5;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A1 = CLBLM_R_X5Y152_SLICE_X6Y152_CO6;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A2 = CLBLM_R_X7Y150_SLICE_X8Y150_BQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A3 = CLBLM_R_X5Y151_SLICE_X6Y151_AQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A5 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_A6 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B1 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B2 = CLBLM_R_X5Y151_SLICE_X6Y151_BQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B3 = CLBLM_R_X5Y152_SLICE_X6Y152_CO5;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B5 = CLBLM_R_X5Y150_SLICE_X7Y150_BQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_B6 = CLBLM_R_X5Y150_SLICE_X6Y150_CQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C2 = CLBLM_R_X5Y148_SLICE_X6Y148_AQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C3 = CLBLM_R_X7Y153_SLICE_X8Y153_CQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C4 = CLBLM_R_X7Y153_SLICE_X8Y153_BQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_C6 = 1'b1;
  assign CLBLM_L_X10Y157_SLICE_X12Y157_A2 = 1'b1;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y157_SLICE_X12Y157_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D1 = CLBLM_R_X5Y149_SLICE_X6Y149_CO5;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D2 = CLBLM_L_X12Y149_SLICE_X17Y149_A5Q;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D3 = CLBLM_R_X5Y151_SLICE_X6Y151_DQ;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y151_SLICE_X6Y151_D6 = CLBLL_L_X4Y154_SLICE_X4Y154_BO6;
  assign CLBLM_L_X10Y157_SLICE_X12Y157_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_D5 = CLBLM_R_X7Y153_SLICE_X8Y153_AQ;
  assign CLBLM_L_X10Y157_SLICE_X12Y157_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y157_SLICE_X12Y157_B5 = 1'b1;
  assign CLBLM_L_X10Y157_SLICE_X12Y157_B6 = CLBLM_R_X7Y157_SLICE_X9Y157_DQ;
  assign CLBLM_L_X10Y157_SLICE_X12Y157_C4 = CLBLM_R_X11Y156_SLICE_X14Y156_BQ;
  assign CLBLM_L_X10Y157_SLICE_X12Y157_C5 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B2 = CLBLM_R_X11Y153_SLICE_X15Y153_BQ;
  assign CLBLM_L_X10Y157_SLICE_X12Y157_C6 = 1'b1;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_A6 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B3 = CLBLM_R_X11Y153_SLICE_X15Y153_CQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y159_SLICE_X15Y159_C4 = CLBLM_L_X12Y158_SLICE_X16Y158_AQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C2 = CLBLM_R_X11Y153_SLICE_X15Y153_CQ;
  assign CLBLM_L_X10Y157_SLICE_X12Y157_D2 = CLBLM_L_X8Y156_SLICE_X11Y156_AQ;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_C5 = CLBLM_L_X10Y152_SLICE_X13Y152_AQ;
  assign CLBLM_L_X10Y157_SLICE_X12Y157_D3 = CLBLM_L_X10Y158_SLICE_X12Y158_BQ;
  assign CLBLM_R_X11Y159_SLICE_X15Y159_C5 = CLBLM_R_X11Y159_SLICE_X15Y159_AQ;
  assign CLBLM_R_X11Y159_SLICE_X15Y159_C6 = 1'b1;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_AX = CLBLM_R_X11Y158_SLICE_X14Y158_BQ;
  assign RIOB33_X105Y169_IOB_X1Y170_O = CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  assign RIOB33_X105Y169_IOB_X1Y169_O = CLBLM_R_X103Y169_SLICE_X163Y169_AO6;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_A1 = CLBLM_R_X5Y152_SLICE_X6Y152_CO6;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_A3 = CLBLM_R_X5Y152_SLICE_X7Y152_AQ;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_A4 = CLBLM_R_X5Y149_SLICE_X7Y149_AQ;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_A5 = CLBLM_L_X8Y151_SLICE_X11Y151_AQ;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_A6 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_B1 = CLBLM_R_X7Y149_SLICE_X8Y149_CQ;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_B2 = CLBLM_R_X5Y152_SLICE_X7Y152_BQ;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_B3 = CLBLM_R_X5Y152_SLICE_X6Y152_CO5;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_B5 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_B6 = CLBLM_L_X10Y152_SLICE_X12Y152_AQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A1 = LIOB33_X0Y51_IOB_X0Y51_I;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A3 = CLBLL_L_X4Y151_SLICE_X4Y151_CQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A4 = CLBLL_L_X4Y152_SLICE_X4Y152_AQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A5 = CLBLL_L_X4Y153_SLICE_X4Y153_AO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_A6 = CLBLM_R_X3Y156_SLICE_X2Y156_DO6;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_C1 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_C2 = CLBLM_R_X7Y150_SLICE_X8Y150_CO6;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_C3 = CLBLM_R_X5Y152_SLICE_X7Y152_DQ;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B1 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B2 = CLBLL_L_X4Y148_SLICE_X4Y148_CO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B3 = CLBLL_L_X4Y147_SLICE_X4Y147_AO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B4 = CLBLL_L_X4Y154_SLICE_X4Y154_BO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B5 = CLBLM_R_X3Y142_SLICE_X3Y142_AO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_D1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C1 = CLBLM_R_X3Y142_SLICE_X3Y142_AO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C2 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C4 = CLBLL_L_X4Y147_SLICE_X4Y147_AO6;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C5 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_C6 = CLBLL_L_X4Y154_SLICE_X4Y154_BO6;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_D4 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_D5 = CLBLM_R_X5Y151_SLICE_X7Y151_DQ;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_A1 = CLBLM_L_X10Y150_SLICE_X13Y150_CQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_A2 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D1 = CLBLM_R_X3Y152_SLICE_X3Y152_AO5;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D2 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D3 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D4 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X3Y142_D6 = CLBLL_L_X4Y148_SLICE_X4Y148_CO6;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_B1 = CLBLM_R_X7Y149_SLICE_X8Y149_CQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_B2 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_B4 = CLBLL_L_X4Y152_SLICE_X5Y152_AQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_B5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A2 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A3 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A4 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_A6 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_C6 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B3 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B2 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B6 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_D1 = CLBLM_R_X5Y150_SLICE_X6Y150_BQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_D2 = CLBLL_L_X2Y155_SLICE_X1Y155_CO6;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_D3 = CLBLM_R_X5Y151_SLICE_X6Y151_BQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_D4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_D5 = CLBLM_R_X3Y156_SLICE_X3Y156_AO5;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_D6 = CLBLM_R_X3Y158_SLICE_X2Y158_AO5;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C3 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C2 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C4 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_C6 = 1'b1;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_B3 = CLBLM_L_X12Y158_SLICE_X16Y158_CO5;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D1 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D2 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D3 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D4 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D5 = 1'b1;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_D6 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_C2 = CLBLL_L_X4Y149_SLICE_X4Y149_CO6;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_D1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign LIOI3_X0Y183_OLOGIC_X0Y184_T1 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = CLBLM_R_X5Y148_SLICE_X7Y148_B5Q;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_D1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_D1 = CLBLM_L_X10Y163_SLICE_X13Y163_AO6;
  assign LIOI3_X0Y183_OLOGIC_X0Y183_T1 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_D5 = CLBLL_L_X2Y155_SLICE_X1Y155_BO5;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = CLBLM_L_X8Y146_SLICE_X10Y146_B5Q;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_D6 = CLBLM_L_X8Y156_SLICE_X10Y156_BQ;
  assign RIOI3_X105Y167_OLOGIC_X1Y168_T1 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_D1 = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_D1 = CLBLM_R_X3Y151_SLICE_X3Y151_BO6;
  assign RIOI3_X105Y167_OLOGIC_X1Y167_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y108_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_D1 = CLBLM_R_X3Y142_SLICE_X3Y142_CO6;
  assign CLBLM_R_X11Y159_SLICE_X15Y159_D2 = CLBLM_R_X11Y157_SLICE_X15Y157_AQ;
  assign LIOI3_TBYTESRC_X0Y107_OLOGIC_X0Y107_T1 = 1'b1;
  assign RIOB33_X105Y171_IOB_X1Y172_O = CLBLM_R_X103Y172_SLICE_X163Y172_AO6;
  assign RIOB33_X105Y171_IOB_X1Y171_O = CLBLM_L_X12Y159_SLICE_X16Y159_CO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D4 = CLBLM_R_X11Y153_SLICE_X14Y153_CO6;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D5 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X14Y153_D6 = CLBLM_R_X5Y147_SLICE_X7Y147_BQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_A1 = CLBLM_L_X12Y154_SLICE_X16Y154_AQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_A3 = CLBLM_R_X5Y153_SLICE_X7Y153_AQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_A4 = CLBLM_R_X5Y153_SLICE_X7Y153_BO6;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_A5 = CLBLM_R_X5Y153_SLICE_X7Y153_CO6;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_C1 = CLBLM_R_X13Y157_SLICE_X19Y157_AQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_B1 = CLBLM_R_X5Y152_SLICE_X7Y152_DQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_B3 = CLBLM_L_X8Y150_SLICE_X11Y150_AQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_B4 = CLBLM_R_X7Y156_SLICE_X9Y156_BQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_B5 = CLBLM_L_X8Y153_SLICE_X11Y153_DQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_B6 = CLBLM_R_X5Y152_SLICE_X7Y152_CQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_C1 = CLBLM_R_X5Y157_SLICE_X7Y157_DQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_C2 = CLBLM_R_X7Y150_SLICE_X8Y150_BQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_C3 = CLBLM_R_X7Y153_SLICE_X9Y153_DO6;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_C4 = CLBLM_R_X5Y150_SLICE_X7Y150_BQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_C5 = CLBLM_R_X5Y153_SLICE_X7Y153_DO6;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_C6 = CLBLM_R_X5Y152_SLICE_X6Y152_AQ;
  assign CLBLM_R_X11Y159_SLICE_X15Y159_D5 = CLBLM_L_X12Y158_SLICE_X16Y158_AQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_C2 = CLBLM_R_X11Y157_SLICE_X14Y157_BQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_D1 = CLBLM_R_X5Y154_SLICE_X6Y154_AQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_D2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_D3 = 1'b1;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_D4 = CLBLM_L_X12Y149_SLICE_X16Y149_CQ;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_D5 = 1'b1;
  assign CLBLM_R_X5Y153_SLICE_X7Y153_D6 = CLBLM_L_X10Y152_SLICE_X12Y152_AQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_A1 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_A3 = CLBLM_R_X5Y153_SLICE_X6Y153_AQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_A4 = CLBLM_L_X12Y150_SLICE_X16Y150_CQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_A5 = CLBLL_L_X4Y151_SLICE_X5Y151_AQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y159_SLICE_X15Y159_D6 = 1'b1;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_B2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_B3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_B4 = CLBLL_L_X4Y157_SLICE_X4Y157_CO5;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_B5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_B6 = 1'b1;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_C3 = CLBLM_R_X13Y157_SLICE_X19Y157_BO6;
  assign LIOB33_X0Y155_IOB_X0Y155_O = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_C1 = CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_C2 = CLBLM_R_X5Y148_SLICE_X7Y148_CO6;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_C3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_C4 = CLBLM_R_X3Y153_SLICE_X3Y153_AO5;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_C5 = 1'b1;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_C6 = CLBLM_L_X8Y157_SLICE_X10Y157_CQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_C4 = CLBLM_R_X11Y158_SLICE_X15Y158_DO6;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_D1 = CLBLM_R_X3Y157_SLICE_X2Y157_AO6;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_D2 = CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_D3 = CLBLM_R_X3Y154_SLICE_X3Y154_AO6;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_D4 = 1'b1;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_D5 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y153_SLICE_X6Y153_D6 = CLBLM_R_X5Y152_SLICE_X6Y152_DO6;
  assign LIOI3_X0Y61_ILOGIC_X0Y62_D = LIOB33_X0Y61_IOB_X0Y62_I;
  assign LIOI3_X0Y61_ILOGIC_X0Y61_D = LIOB33_X0Y61_IOB_X0Y61_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_D = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_C5 = CLBLM_R_X13Y157_SLICE_X18Y157_DO6;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_D = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A4 = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_A6 = 1'b1;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_C6 = CLBLM_L_X12Y158_SLICE_X16Y158_BO5;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y114_D = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_B6 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_D4 = CLBLM_R_X7Y156_SLICE_X8Y156_CQ;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_D5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_C6 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X8Y155_D6 = CLBLM_R_X7Y156_SLICE_X8Y156_BQ;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X78Y126_D6 = 1'b1;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_T1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_A6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_B6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_C6 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D1 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D2 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D3 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D4 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D5 = 1'b1;
  assign CLBLL_L_X52Y126_SLICE_X79Y126_D6 = 1'b1;
  assign RIOB33_X105Y173_IOB_X1Y174_O = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign RIOB33_X105Y173_IOB_X1Y173_O = CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_A1 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_A2 = CLBLM_L_X10Y146_SLICE_X12Y146_C5Q;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_A3 = CLBLM_R_X5Y154_SLICE_X7Y154_AQ;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_A5 = CLBLM_R_X5Y152_SLICE_X6Y152_CO5;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_A6 = CLBLM_R_X5Y152_SLICE_X6Y152_AQ;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_B2 = CLBLL_L_X4Y157_SLICE_X4Y157_CO5;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_B3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_B4 = CLBLM_R_X11Y153_SLICE_X15Y153_BQ;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_B5 = CLBLM_L_X8Y153_SLICE_X11Y153_AQ;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_B6 = CLBLL_L_X4Y157_SLICE_X4Y157_AO5;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_C1 = CLBLL_L_X2Y155_SLICE_X1Y155_BO5;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_C2 = CLBLM_R_X5Y155_SLICE_X7Y155_AQ;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_C3 = CLBLM_R_X3Y153_SLICE_X3Y153_AO6;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_C4 = CLBLM_R_X3Y154_SLICE_X3Y154_AO5;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_C5 = CLBLM_R_X7Y149_SLICE_X9Y149_BQ;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_C6 = CLBLM_L_X10Y154_SLICE_X12Y154_AQ;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOB33_X0Y163_IOB_X0Y164_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_D1 = CLBLL_L_X2Y155_SLICE_X1Y155_BO5;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_D2 = CLBLM_R_X3Y157_SLICE_X2Y157_AO5;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_D3 = CLBLM_R_X5Y151_SLICE_X7Y151_AQ;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_D4 = CLBLM_R_X5Y148_SLICE_X7Y148_AQ;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_D5 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X7Y154_D6 = CLBLM_R_X5Y154_SLICE_X7Y154_BO6;
  assign LIOB33_X0Y163_IOB_X0Y163_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_A1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_A3 = CLBLM_R_X5Y154_SLICE_X6Y154_AQ;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_A4 = CLBLM_R_X5Y151_SLICE_X6Y151_DQ;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_A6 = CLBLM_L_X12Y149_SLICE_X16Y149_CQ;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_B1 = CLBLM_R_X11Y155_SLICE_X14Y155_AQ;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_B2 = CLBLL_L_X2Y155_SLICE_X1Y155_BO5;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_B3 = CLBLM_R_X3Y157_SLICE_X2Y157_AO5;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_B4 = CLBLM_R_X3Y154_SLICE_X3Y154_AO5;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_B5 = CLBLL_L_X4Y148_SLICE_X5Y148_AQ;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_B6 = CLBLM_R_X5Y151_SLICE_X6Y151_DQ;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_C1 = CLBLM_R_X3Y157_SLICE_X2Y157_AO6;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_C2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_C3 = CLBLM_R_X7Y154_SLICE_X9Y154_AQ;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_C4 = CLBLM_R_X5Y150_SLICE_X6Y150_CQ;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_C5 = CLBLL_L_X4Y156_SLICE_X4Y156_CO6;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_C6 = CLBLM_R_X5Y153_SLICE_X6Y153_BO6;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_D1 = CLBLM_R_X5Y154_SLICE_X7Y154_AQ;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_D2 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_D3 = CLBLL_L_X4Y151_SLICE_X5Y151_AQ;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_D4 = 1'b1;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_D5 = CLBLL_L_X4Y157_SLICE_X4Y157_BO5;
  assign CLBLM_R_X5Y154_SLICE_X6Y154_D6 = CLBLM_R_X5Y153_SLICE_X6Y153_BO6;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_D1 = CLBLM_R_X11Y158_SLICE_X14Y158_AQ;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_D2 = CLBLM_R_X13Y158_SLICE_X18Y158_BQ;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_D3 = CLBLM_R_X13Y159_SLICE_X18Y159_DO6;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_D4 = CLBLM_R_X11Y157_SLICE_X15Y157_BQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_D5 = CLBLM_R_X11Y157_SLICE_X14Y157_AQ;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_D1 = CLBLM_L_X12Y156_SLICE_X16Y156_AQ;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B1 = 1'b1;
  assign RIOB33_X105Y175_IOB_X1Y176_O = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign RIOB33_X105Y175_IOB_X1Y175_O = CLBLM_R_X13Y157_SLICE_X18Y157_AO5;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B2 = 1'b1;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_D6 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B3 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B4 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B5 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_B6 = 1'b1;
  assign CLBLM_R_X7Y145_SLICE_X8Y145_C1 = 1'b1;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_D1 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign LIOI3_X0Y185_OLOGIC_X0Y186_T1 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_D1 = CLBLL_L_X4Y147_SLICE_X5Y147_AQ;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_D1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_T1 = 1'b1;
  assign CLBLM_R_X11Y159_SLICE_X14Y159_B5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_A1 = CLBLL_L_X4Y151_SLICE_X4Y151_DQ;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_A2 = CLBLM_R_X7Y153_SLICE_X9Y153_CO6;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_A3 = CLBLM_R_X5Y155_SLICE_X7Y155_AQ;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_A4 = 1'b1;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_A6 = CLBLM_L_X8Y156_SLICE_X10Y156_CQ;
  assign LIOI3_X0Y185_OLOGIC_X0Y185_T1 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_D1 = CLBLM_L_X8Y154_SLICE_X10Y154_C5Q;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_B1 = CLBLM_R_X5Y151_SLICE_X7Y151_CQ;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_B2 = CLBLM_R_X5Y155_SLICE_X7Y155_BQ;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_B4 = CLBLM_L_X10Y150_SLICE_X12Y150_A5Q;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_B5 = CLBLM_L_X12Y155_SLICE_X16Y155_CO6;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_B6 = CLBLM_L_X8Y155_SLICE_X10Y155_B5Q;
  assign RIOI3_X105Y171_OLOGIC_X1Y172_T1 = 1'b1;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_C1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_C2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_C3 = CLBLL_L_X4Y157_SLICE_X4Y157_CO5;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_C4 = CLBLM_L_X8Y155_SLICE_X11Y155_AQ;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_C5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_C6 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X11Y159_SLICE_X14Y159_B6 = CLBLM_L_X8Y155_SLICE_X10Y155_CQ;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_T1 = 1'b1;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_SR = CLBLM_R_X13Y155_SLICE_X18Y155_DO6;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_D1 = CLBLM_L_X12Y159_SLICE_X16Y159_CO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = CLBLM_L_X12Y149_SLICE_X16Y149_BQ;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_D1 = CLBLM_R_X5Y155_SLICE_X6Y155_AQ;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_D2 = CLBLM_R_X5Y151_SLICE_X7Y151_DQ;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_D3 = CLBLM_R_X3Y153_SLICE_X3Y153_AO6;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_D4 = CLBLM_R_X5Y155_SLICE_X7Y155_CO6;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_D5 = CLBLM_R_X3Y157_SLICE_X2Y157_AO5;
  assign CLBLM_R_X5Y155_SLICE_X7Y155_D6 = CLBLM_R_X7Y159_SLICE_X9Y159_DO6;
  assign RIOI3_X105Y171_OLOGIC_X1Y171_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_A2 = CLBLM_L_X8Y155_SLICE_X11Y155_BQ;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_A3 = CLBLM_R_X5Y155_SLICE_X6Y155_AQ;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_A4 = CLBLM_R_X7Y153_SLICE_X9Y153_CO6;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_A5 = CLBLM_R_X3Y151_SLICE_X3Y151_AQ;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = CLBLM_R_X11Y149_SLICE_X15Y149_AQ;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_B1 = CLBLM_R_X7Y155_SLICE_X9Y155_DO6;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_B2 = CLBLM_R_X3Y154_SLICE_X3Y154_DO6;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_B3 = CLBLM_R_X13Y155_SLICE_X19Y155_AO6;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_B4 = CLBLM_R_X5Y156_SLICE_X6Y156_BO6;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_B5 = CLBLL_L_X4Y156_SLICE_X4Y156_CO5;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_B6 = CLBLM_R_X5Y155_SLICE_X6Y155_CO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_C1 = CLBLM_R_X3Y157_SLICE_X2Y157_AO6;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_C2 = CLBLL_L_X4Y155_SLICE_X5Y155_CO6;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_C3 = CLBLL_L_X4Y156_SLICE_X4Y156_CO5;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_C4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_C5 = CLBLL_L_X4Y156_SLICE_X5Y156_DO6;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_C6 = CLBLM_L_X8Y155_SLICE_X10Y155_CQ;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_D1 = CLBLM_R_X7Y155_SLICE_X9Y155_DO6;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_D2 = 1'b1;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_D3 = CLBLL_L_X4Y156_SLICE_X4Y156_CO5;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_D4 = CLBLM_R_X5Y155_SLICE_X6Y155_CO6;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_D5 = CLBLM_R_X3Y154_SLICE_X3Y154_DO6;
  assign CLBLM_R_X5Y155_SLICE_X6Y155_D6 = CLBLM_R_X5Y156_SLICE_X6Y156_BO6;
  assign CLBLM_L_X12Y156_SLICE_X17Y156_C3 = CLBLM_L_X12Y158_SLICE_X16Y158_BO5;
  assign CLBLM_L_X12Y156_SLICE_X17Y156_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X12Y156_SLICE_X17Y156_D3 = CLBLM_L_X12Y157_SLICE_X16Y157_CQ;
  assign CLBLM_L_X10Y158_SLICE_X13Y158_A6 = CLBLM_R_X11Y157_SLICE_X14Y157_CQ;
  assign CLBLM_L_X12Y156_SLICE_X17Y156_D6 = CLBLM_R_X13Y149_SLICE_X18Y149_A5Q;
  assign RIOB33_X105Y177_IOB_X1Y178_O = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign RIOB33_X105Y177_IOB_X1Y177_O = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y193_T1 = 1'b1;
  assign LIOI3_X0Y65_ILOGIC_X0Y66_D = LIOB33_X0Y65_IOB_X0Y66_I;
  assign CLBLM_L_X10Y158_SLICE_X13Y158_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_X0Y65_ILOGIC_X0Y65_D = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLM_L_X10Y158_SLICE_X13Y158_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y158_SLICE_X13Y158_B3 = CLBLM_L_X12Y152_SLICE_X17Y152_AQ;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_D = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X10Y158_SLICE_X13Y158_B4 = 1'b1;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_D = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X12Y156_SLICE_X16Y156_A6 = CLBLM_L_X10Y157_SLICE_X12Y157_DO6;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y138_D = RIOB33_X105Y137_IOB_X1Y138_I;
  assign RIOI3_TBYTETERM_X105Y137_ILOGIC_X1Y137_D = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X5Y156_SLICE_X7Y156_A1 = CLBLM_R_X7Y153_SLICE_X8Y153_A5Q;
  assign CLBLM_R_X5Y156_SLICE_X7Y156_A2 = CLBLM_L_X12Y158_SLICE_X16Y158_A5Q;
  assign CLBLM_R_X5Y156_SLICE_X7Y156_A3 = CLBLM_R_X5Y156_SLICE_X7Y156_AQ;
  assign CLBLM_R_X5Y156_SLICE_X7Y156_A4 = CLBLL_L_X4Y147_SLICE_X4Y147_BO6;
  assign CLBLM_R_X5Y156_SLICE_X7Y156_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y156_SLICE_X7Y156_A6 = 1'b1;
  assign CLBLM_L_X12Y156_SLICE_X16Y156_BX = CLBLM_R_X11Y146_SLICE_X15Y146_BQ;
  assign CLBLM_R_X5Y156_SLICE_X7Y156_B1 = CLBLM_R_X7Y157_SLICE_X9Y157_BQ;
  assign CLBLM_R_X3Y142_SLICE_X2Y142_B4 = 1'b1;
  assign CLBLM_R_X5Y156_SLICE_X7Y156_B2 = CLBLM_R_X5Y152_SLICE_X7Y152_BQ;
  assign CLBLM_R_X5Y156_SLICE_X7Y156_B3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y156_SLICE_X7Y156_B4 = CLBLL_L_X4Y157_SLICE_X4Y157_CO5;
  assign CLBLM_R_X5Y156_SLICE_X7Y156_B5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X5Y156_SLICE_X7Y156_B6 = CLBLL_L_X4Y157_SLICE_X4Y157_AO5;
  assign CLBLM_R_X7Y159_SLICE_X9Y159_C4 = CLBLM_R_X3Y152_SLICE_X3Y152_BO5;
  assign CLBLM_R_X5Y156_SLICE_X7Y156_C1 = CLBLL_L_X2Y155_SLICE_X1Y155_CO6;
  assign CLBLM_R_X5Y156_SLICE_X7Y156_C2 = 1'b1;
  assign CLBLM_R_X5Y156_SLICE_X7Y156_C3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X5Y156_SLICE_X7Y156_C4 = CLBLM_R_X3Y156_SLICE_X3Y156_AO5;
  assign CLBLM_R_X5Y156_SLICE_X7Y156_C5 = CLBLM_R_X3Y158_SLICE_X2Y158_AO6;
  assign CLBLM_R_X5Y156_SLICE_X7Y156_C6 = CLBLM_L_X8Y154_SLICE_X10Y154_DQ;
  assign CLBLM_R_X5Y156_SLICE_X7Y156_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X12Y156_SLICE_X16Y156_C3 = CLBLM_L_X8Y154_SLICE_X10Y154_AQ;
  assign CLBLM_R_X5Y156_SLICE_X7Y156_D1 = CLBLM_R_X7Y156_SLICE_X9Y156_AQ;
  assign CLBLM_R_X5Y156_SLICE_X7Y156_D2 = 1'b1;
  assign CLBLM_R_X5Y156_SLICE_X7Y156_D3 = CLBLM_R_X5Y157_SLICE_X6Y157_BO6;
  assign CLBLM_R_X5Y156_SLICE_X7Y156_D4 = CLBLM_R_X5Y156_SLICE_X7Y156_CO6;
  assign CLBLM_R_X5Y156_SLICE_X7Y156_D5 = CLBLM_R_X3Y154_SLICE_X3Y154_AO6;
  assign CLBLM_R_X5Y156_SLICE_X7Y156_D6 = CLBLM_R_X5Y156_SLICE_X7Y156_BO6;
  assign CLBLM_R_X7Y159_SLICE_X9Y159_C5 = CLBLM_L_X8Y154_SLICE_X10Y154_A5Q;
  assign RIOI3_X105Y165_OLOGIC_X1Y166_D1 = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign CLBLM_R_X5Y156_SLICE_X6Y156_A1 = CLBLM_R_X5Y156_SLICE_X6Y156_DO6;
  assign CLBLM_L_X12Y156_SLICE_X16Y156_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y156_SLICE_X6Y156_A2 = CLBLM_R_X5Y155_SLICE_X7Y155_BQ;
  assign CLBLM_R_X5Y156_SLICE_X6Y156_A3 = CLBLL_L_X4Y156_SLICE_X5Y156_DO6;
  assign CLBLM_R_X5Y156_SLICE_X6Y156_A4 = CLBLL_L_X4Y156_SLICE_X4Y156_CO6;
  assign CLBLM_R_X5Y156_SLICE_X6Y156_A5 = CLBLL_L_X4Y155_SLICE_X5Y155_CO6;
  assign CLBLM_R_X5Y156_SLICE_X6Y156_A6 = CLBLM_R_X5Y156_SLICE_X6Y156_CO6;
  assign CLBLM_R_X5Y156_SLICE_X6Y156_B1 = CLBLL_L_X4Y156_SLICE_X4Y156_CO6;
  assign CLBLM_R_X5Y156_SLICE_X6Y156_B2 = CLBLM_R_X5Y155_SLICE_X7Y155_BQ;
  assign CLBLM_R_X5Y156_SLICE_X6Y156_B3 = CLBLM_R_X5Y151_SLICE_X6Y151_AQ;
  assign CLBLM_R_X5Y156_SLICE_X6Y156_B4 = CLBLL_L_X4Y157_SLICE_X4Y157_BO6;
  assign CLBLM_R_X5Y156_SLICE_X6Y156_B5 = CLBLM_R_X7Y148_SLICE_X9Y148_AQ;
  assign CLBLM_R_X5Y156_SLICE_X6Y156_B6 = CLBLM_R_X3Y154_SLICE_X3Y154_AO6;
  assign CLBLM_R_X7Y159_SLICE_X9Y159_C6 = CLBLM_L_X8Y158_SLICE_X10Y158_AQ;
  assign LIOB33_X0Y139_IOB_X0Y140_O = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLM_R_X5Y156_SLICE_X6Y156_C1 = CLBLM_R_X7Y148_SLICE_X9Y148_AQ;
  assign CLBLM_R_X5Y156_SLICE_X6Y156_C2 = CLBLM_R_X5Y151_SLICE_X6Y151_AQ;
  assign CLBLM_R_X5Y156_SLICE_X6Y156_C3 = CLBLL_L_X4Y157_SLICE_X4Y157_CO5;
  assign CLBLM_R_X5Y156_SLICE_X6Y156_C4 = CLBLL_L_X2Y155_SLICE_X1Y155_CO6;
  assign CLBLM_R_X5Y156_SLICE_X6Y156_C5 = 1'b1;
  assign CLBLM_R_X5Y156_SLICE_X6Y156_C6 = CLBLL_L_X2Y155_SLICE_X1Y155_CO5;
  assign LIOB33_X0Y139_IOB_X0Y139_O = CLBLM_R_X5Y144_SLICE_X6Y144_AQ;
  assign CLBLM_R_X5Y156_SLICE_X6Y156_D1 = CLBLM_L_X8Y155_SLICE_X10Y155_CQ;
  assign CLBLM_R_X5Y156_SLICE_X6Y156_D2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X5Y156_SLICE_X6Y156_D3 = CLBLM_R_X3Y158_SLICE_X2Y158_AO6;
  assign CLBLM_R_X5Y156_SLICE_X6Y156_D4 = CLBLL_L_X2Y155_SLICE_X1Y155_CO6;
  assign CLBLM_R_X5Y156_SLICE_X6Y156_D5 = 1'b1;
  assign CLBLM_R_X5Y156_SLICE_X6Y156_D6 = CLBLL_L_X2Y155_SLICE_X1Y155_CO5;
  assign CLBLM_L_X10Y158_SLICE_X12Y158_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y158_SLICE_X12Y158_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y156_SLICE_X16Y156_D2 = CLBLM_R_X13Y156_SLICE_X18Y156_CO6;
  assign CLBLM_L_X10Y158_SLICE_X12Y158_A6 = 1'b1;
  assign CLBLM_L_X12Y156_SLICE_X16Y156_D3 = CLBLM_L_X12Y158_SLICE_X16Y158_BO5;
  assign CLBLM_L_X12Y156_SLICE_X16Y156_D4 = CLBLM_R_X11Y158_SLICE_X15Y158_DO6;
  assign CLBLM_R_X13Y155_SLICE_X18Y155_D6 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign RIOI3_X105Y139_ILOGIC_X1Y140_D = RIOB33_X105Y139_IOB_X1Y140_I;
  assign CLBLM_L_X10Y158_SLICE_X12Y158_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOB33_X105Y179_IOB_X1Y180_O = CLBLM_R_X13Y154_SLICE_X18Y154_DO6;
  assign RIOB33_X105Y179_IOB_X1Y179_O = CLBLM_L_X12Y159_SLICE_X16Y159_AO5;
  assign CLBLM_L_X10Y158_SLICE_X12Y158_B5 = CLBLM_R_X11Y153_SLICE_X15Y153_AQ;
  assign CLBLM_L_X10Y158_SLICE_X12Y158_B6 = CLBLM_L_X10Y158_SLICE_X12Y158_CO6;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y139_ILOGIC_X1Y139_D = RIOB33_X105Y139_IOB_X1Y139_I;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_A4 = 1'b1;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_A6 = CLBLM_R_X13Y151_SLICE_X18Y151_CQ;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_B4 = CLBLM_R_X11Y158_SLICE_X15Y158_BO6;
  assign CLBLM_L_X10Y158_SLICE_X12Y158_C4 = CLBLM_L_X10Y153_SLICE_X12Y153_AQ;
  assign CLBLM_L_X10Y158_SLICE_X12Y158_C5 = CLBLM_L_X10Y157_SLICE_X12Y157_CO5;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_B5 = CLBLM_R_X11Y158_SLICE_X14Y158_BQ;
  assign CLBLM_L_X10Y158_SLICE_X12Y158_C6 = CLBLM_L_X10Y156_SLICE_X13Y156_CO6;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_B4 = CLBLM_R_X7Y153_SLICE_X8Y153_AQ;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_B6 = CLBLM_L_X8Y150_SLICE_X10Y150_BQ;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_B6 = CLBLM_R_X11Y157_SLICE_X14Y157_BQ;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_C2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_C3 = CLBLM_R_X11Y154_SLICE_X14Y154_D5Q;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_C4 = CLBLM_L_X10Y155_SLICE_X13Y155_BQ;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_C5 = CLBLM_R_X11Y151_SLICE_X15Y151_AQ;
  assign CLBLM_L_X10Y158_SLICE_X12Y158_D3 = 1'b1;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_C6 = 1'b1;
  assign CLBLM_L_X10Y158_SLICE_X12Y158_D6 = 1'b1;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X5Y157_SLICE_X7Y157_A1 = CLBLM_R_X5Y157_SLICE_X7Y157_CQ;
  assign CLBLM_R_X5Y157_SLICE_X7Y157_A2 = 1'b1;
  assign CLBLM_R_X5Y157_SLICE_X7Y157_A3 = CLBLM_R_X5Y157_SLICE_X7Y157_AQ;
  assign CLBLM_R_X5Y157_SLICE_X7Y157_A4 = CLBLM_L_X10Y153_SLICE_X13Y153_CQ;
  assign CLBLM_R_X5Y157_SLICE_X7Y157_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y157_SLICE_X7Y157_A6 = CLBLM_R_X7Y153_SLICE_X9Y153_CO6;
  assign CLBLM_R_X5Y157_SLICE_X7Y157_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y157_SLICE_X7Y157_B2 = CLBLM_R_X5Y157_SLICE_X7Y157_BQ;
  assign CLBLM_R_X5Y157_SLICE_X7Y157_B3 = CLBLM_R_X7Y151_SLICE_X8Y151_AQ;
  assign CLBLM_R_X5Y157_SLICE_X7Y157_B4 = CLBLM_R_X5Y152_SLICE_X6Y152_CO5;
  assign CLBLM_R_X5Y157_SLICE_X7Y157_B5 = CLBLM_L_X8Y157_SLICE_X10Y157_AQ;
  assign CLBLM_R_X5Y157_SLICE_X7Y157_B6 = 1'b1;
  assign CLBLM_R_X5Y157_SLICE_X7Y157_C1 = CLBLM_R_X5Y152_SLICE_X6Y152_CO5;
  assign CLBLM_R_X5Y157_SLICE_X7Y157_C2 = CLBLM_R_X5Y157_SLICE_X7Y157_CQ;
  assign CLBLM_R_X5Y157_SLICE_X7Y157_C3 = 1'b1;
  assign CLBLM_R_X5Y157_SLICE_X7Y157_C4 = CLBLM_R_X7Y156_SLICE_X9Y156_BQ;
  assign CLBLM_R_X5Y157_SLICE_X7Y157_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y157_SLICE_X7Y157_C6 = CLBLM_R_X5Y154_SLICE_X7Y154_AQ;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_D1 = CLBLM_R_X11Y146_SLICE_X15Y146_AQ;
  assign CLBLM_R_X5Y157_SLICE_X7Y157_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_D2 = CLBLL_L_X4Y155_SLICE_X4Y155_CO6;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_D3 = CLBLM_R_X11Y156_SLICE_X15Y156_DO6;
  assign CLBLM_R_X5Y157_SLICE_X7Y157_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y157_SLICE_X7Y157_D2 = 1'b1;
  assign CLBLM_R_X5Y157_SLICE_X7Y157_D3 = CLBLM_R_X5Y149_SLICE_X7Y149_DO6;
  assign CLBLM_R_X5Y157_SLICE_X7Y157_D4 = CLBLM_R_X5Y157_SLICE_X7Y157_BQ;
  assign CLBLM_R_X5Y157_SLICE_X7Y157_D5 = CLBLM_L_X8Y153_SLICE_X11Y153_DQ;
  assign CLBLM_R_X5Y157_SLICE_X7Y157_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y156_SLICE_X9Y156_A4 = CLBLM_L_X12Y155_SLICE_X17Y155_BQ;
  assign CLBLM_R_X7Y156_SLICE_X9Y156_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_D4 = CLBLM_R_X11Y155_SLICE_X15Y155_CO6;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_D5 = CLBLM_R_X13Y152_SLICE_X18Y152_BO5;
  assign CLBLM_R_X7Y156_SLICE_X9Y156_A6 = 1'b1;
  assign CLBLM_R_X5Y157_SLICE_X6Y157_A1 = CLBLM_L_X12Y158_SLICE_X16Y158_A5Q;
  assign CLBLM_R_X5Y157_SLICE_X6Y157_A2 = CLBLM_R_X7Y157_SLICE_X8Y157_AQ;
  assign CLBLM_R_X5Y157_SLICE_X6Y157_A3 = CLBLM_R_X5Y157_SLICE_X6Y157_AQ;
  assign CLBLM_R_X5Y157_SLICE_X6Y157_A4 = 1'b1;
  assign CLBLM_R_X5Y157_SLICE_X6Y157_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y157_SLICE_X6Y157_A6 = CLBLM_R_X7Y153_SLICE_X9Y153_CO6;
  assign CLBLM_R_X11Y154_SLICE_X15Y154_D6 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_R_X5Y157_SLICE_X6Y157_B1 = CLBLL_L_X4Y157_SLICE_X5Y157_AO5;
  assign CLBLM_R_X5Y157_SLICE_X6Y157_B2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y157_SLICE_X6Y157_B3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y157_SLICE_X6Y157_B4 = CLBLM_R_X3Y150_SLICE_X3Y150_AQ;
  assign CLBLM_R_X5Y157_SLICE_X6Y157_B5 = CLBLM_R_X7Y158_SLICE_X9Y158_AQ;
  assign CLBLM_R_X5Y157_SLICE_X6Y157_B6 = CLBLM_R_X3Y158_SLICE_X2Y158_AO5;
  assign CLBLM_R_X5Y157_SLICE_X6Y157_C1 = CLBLM_R_X5Y152_SLICE_X7Y152_AQ;
  assign CLBLM_R_X5Y157_SLICE_X6Y157_C2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X5Y157_SLICE_X6Y157_C3 = CLBLM_R_X7Y157_SLICE_X9Y157_CQ;
  assign CLBLM_R_X5Y157_SLICE_X6Y157_C4 = 1'b1;
  assign CLBLM_R_X5Y157_SLICE_X6Y157_C5 = CLBLL_L_X4Y157_SLICE_X5Y157_AO5;
  assign CLBLM_R_X5Y157_SLICE_X6Y157_C6 = CLBLL_L_X4Y157_SLICE_X4Y157_CO5;
  assign CLBLM_R_X5Y157_SLICE_X6Y157_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y156_SLICE_X9Y156_B3 = CLBLM_L_X8Y152_SLICE_X11Y152_AO6;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_D1 = RIOB33_X105Y147_IOB_X1Y147_I;
  assign CLBLM_R_X5Y157_SLICE_X6Y157_D1 = CLBLL_L_X4Y156_SLICE_X4Y156_AQ;
  assign CLBLM_R_X5Y157_SLICE_X6Y157_D2 = CLBLM_R_X5Y158_SLICE_X7Y158_AO6;
  assign CLBLM_R_X5Y157_SLICE_X6Y157_D3 = CLBLL_L_X4Y156_SLICE_X4Y156_CO5;
  assign CLBLM_R_X5Y157_SLICE_X6Y157_D4 = CLBLM_R_X7Y158_SLICE_X8Y158_AQ;
  assign CLBLM_R_X5Y157_SLICE_X6Y157_D5 = 1'b1;
  assign CLBLM_R_X5Y157_SLICE_X6Y157_D6 = CLBLL_L_X4Y157_SLICE_X4Y157_BO5;
  assign CLBLM_R_X7Y156_SLICE_X9Y156_B4 = CLBLM_L_X8Y156_SLICE_X10Y156_AQ;
  assign CLBLM_R_X7Y156_SLICE_X9Y156_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y189_OLOGIC_X0Y190_T1 = 1'b1;
  assign CLBLM_R_X7Y156_SLICE_X9Y156_B6 = 1'b1;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_A3 = CLBLM_R_X11Y154_SLICE_X14Y154_AQ;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_D1 = CLBLM_R_X3Y151_SLICE_X2Y151_AQ;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_A4 = CLBLM_R_X7Y150_SLICE_X9Y150_BO6;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_D1 = RIOB33_X105Y145_IOB_X1Y146_I;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_T1 = 1'b1;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_D1 = CLBLM_R_X103Y174_SLICE_X163Y174_AO6;
  assign LIOI3_X0Y189_OLOGIC_X0Y189_T1 = 1'b1;
  assign CLBLM_R_X7Y156_SLICE_X9Y156_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_D1 = CLBLL_L_X4Y152_SLICE_X4Y152_AQ;
  assign RIOB33_X105Y181_IOB_X1Y182_O = CLBLM_R_X13Y155_SLICE_X18Y155_CO5;
  assign RIOB33_X105Y181_IOB_X1Y181_O = CLBLM_R_X13Y155_SLICE_X18Y155_CO6;
  assign RIOI3_X105Y173_OLOGIC_X1Y174_T1 = 1'b1;
  assign CLBLM_R_X7Y156_SLICE_X9Y156_C2 = CLBLM_R_X7Y156_SLICE_X9Y156_CQ;
  assign CLBLM_R_X7Y156_SLICE_X9Y156_C3 = CLBLM_R_X5Y147_SLICE_X7Y147_C5Q;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_T1 = 1'b1;
  assign CLBLM_R_X7Y156_SLICE_X9Y156_C4 = CLBLM_R_X11Y157_SLICE_X14Y157_AQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A3 = CLBLM_L_X12Y146_SLICE_X16Y146_AQ;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_D1 = CLBLM_R_X103Y172_SLICE_X163Y172_AO5;
  assign CLBLM_R_X7Y156_SLICE_X9Y156_C5 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A4 = CLBLM_R_X7Y146_SLICE_X9Y146_DO6;
  assign CLBLM_R_X7Y156_SLICE_X9Y156_C6 = CLBLL_L_X4Y147_SLICE_X4Y147_BO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y173_OLOGIC_X1Y173_T1 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A6 = CLBLM_L_X10Y147_SLICE_X13Y147_BQ;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_B4 = CLBLM_L_X10Y154_SLICE_X13Y154_DQ;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1 = 1'b1;
  assign CLBLM_R_X7Y156_SLICE_X9Y156_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_D1 = CLBLM_R_X7Y149_SLICE_X9Y149_DO5;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_B5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1 = CLBLM_L_X10Y144_SLICE_X12Y144_AO5;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y164_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_D1 = CLBLM_L_X12Y155_SLICE_X17Y155_DO5;
  assign CLBLM_R_X7Y156_SLICE_X9Y156_D1 = CLBLM_R_X7Y155_SLICE_X8Y155_AQ;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_TBYTETERM_X105Y163_OLOGIC_X1Y163_T1 = 1'b1;
  assign CLBLM_R_X7Y156_SLICE_X9Y156_D2 = CLBLM_L_X10Y159_SLICE_X12Y159_AO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_C2 = CLBLM_L_X12Y152_SLICE_X16Y152_AQ;
  assign CLBLM_R_X7Y156_SLICE_X9Y156_D3 = CLBLM_L_X8Y154_SLICE_X10Y154_A5Q;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B6 = CLBLM_L_X12Y153_SLICE_X16Y153_AQ;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_C3 = CLBLM_R_X13Y151_SLICE_X18Y151_CQ;
  assign CLBLM_R_X7Y156_SLICE_X9Y156_D4 = CLBLM_R_X7Y155_SLICE_X8Y155_BO5;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y156_SLICE_X9Y156_D5 = CLBLL_L_X4Y156_SLICE_X4Y156_AO5;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_C5 = CLBLM_R_X11Y154_SLICE_X14Y154_BO5;
  assign CLBLM_R_X7Y156_SLICE_X9Y156_D6 = CLBLM_L_X8Y158_SLICE_X10Y158_AQ;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_C6 = 1'b1;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y156_SLICE_X8Y156_A2 = CLBLM_L_X8Y157_SLICE_X11Y157_CQ;
  assign CLBLM_R_X7Y156_SLICE_X8Y156_A3 = CLBLM_R_X7Y156_SLICE_X8Y156_AQ;
  assign CLBLM_R_X7Y156_SLICE_X8Y156_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y156_SLICE_X8Y156_A5 = CLBLL_L_X4Y151_SLICE_X4Y151_BQ;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_D2 = CLBLM_R_X11Y154_SLICE_X14Y154_CQ;
  assign CLBLM_R_X7Y156_SLICE_X8Y156_A6 = CLBLM_L_X10Y148_SLICE_X13Y148_AQ;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_D3 = CLBLM_L_X8Y159_SLICE_X10Y159_AQ;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_D4 = CLBLM_R_X11Y148_SLICE_X14Y148_CQ;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_D5 = CLBLM_L_X12Y157_SLICE_X17Y157_AQ;
  assign CLBLM_R_X11Y154_SLICE_X14Y154_D6 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_A1 = CLBLM_L_X8Y158_SLICE_X11Y158_BQ;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_A2 = CLBLL_L_X4Y157_SLICE_X4Y157_CO5;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_A3 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_A4 = CLBLM_R_X5Y158_SLICE_X6Y158_BQ;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_A5 = CLBLL_L_X2Y155_SLICE_X1Y155_CO5;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_A6 = CLBLL_L_X2Y155_SLICE_X1Y155_CO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D3 = CLBLM_R_X11Y153_SLICE_X15Y153_DQ;
  assign LIOI3_X0Y67_ILOGIC_X0Y68_D = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_R_X7Y156_SLICE_X8Y156_B2 = CLBLM_R_X7Y156_SLICE_X8Y156_BQ;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_B1 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_B2 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_B3 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_B4 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_B5 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_B6 = 1'b1;
  assign CLBLM_R_X7Y156_SLICE_X8Y156_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_D = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_C1 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_C2 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_C3 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_C4 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_C5 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_C6 = 1'b1;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_D = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_D1 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_D2 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_D3 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_D4 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_D5 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X7Y158_D6 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_A1 = CLBLL_L_X4Y153_SLICE_X5Y153_AQ;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_A2 = CLBLM_L_X8Y153_SLICE_X11Y153_AQ;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_A3 = CLBLM_R_X5Y158_SLICE_X6Y158_AQ;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_A5 = CLBLM_R_X5Y152_SLICE_X6Y152_CO5;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_A6 = 1'b1;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D5 = CLBLM_L_X8Y154_SLICE_X10Y154_DQ;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_B1 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_B2 = CLBLM_R_X5Y158_SLICE_X6Y158_BQ;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_B3 = CLBLM_R_X5Y158_SLICE_X6Y158_AQ;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_B5 = CLBLM_R_X5Y152_SLICE_X6Y152_CO5;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_B6 = CLBLM_L_X10Y150_SLICE_X12Y150_CQ;
  assign CLBLM_R_X7Y156_SLICE_X8Y156_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y156_SLICE_X8Y156_C2 = CLBLM_R_X7Y156_SLICE_X8Y156_CQ;
  assign CLBLM_R_X7Y156_SLICE_X8Y156_C3 = CLBLM_R_X7Y157_SLICE_X8Y157_DQ;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_C1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_C2 = CLBLM_R_X3Y158_SLICE_X2Y158_AO5;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_C3 = CLBLM_R_X5Y158_SLICE_X6Y158_AQ;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_C4 = CLBLL_L_X2Y155_SLICE_X1Y155_CO6;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_C5 = CLBLM_R_X7Y153_SLICE_X8Y153_CQ;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_C6 = CLBLM_R_X3Y156_SLICE_X3Y156_AO5;
  assign CLBLM_R_X7Y156_SLICE_X8Y156_C4 = CLBLM_R_X7Y155_SLICE_X8Y155_BO6;
  assign CLBLM_R_X11Y153_SLICE_X15Y153_D6 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y156_SLICE_X8Y156_C5 = 1'b1;
  assign CLBLM_R_X7Y156_SLICE_X8Y156_C6 = CLBLM_R_X7Y158_SLICE_X8Y158_BQ;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_D1 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_D2 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_D3 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_D4 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_D5 = 1'b1;
  assign CLBLM_R_X5Y158_SLICE_X6Y158_D6 = 1'b1;
  assign RIOB33_X105Y183_IOB_X1Y184_O = CLBLM_L_X12Y155_SLICE_X17Y155_DO5;
  assign RIOB33_X105Y183_IOB_X1Y183_O = CLBLM_L_X12Y155_SLICE_X17Y155_DO6;
  assign CLBLM_R_X7Y156_SLICE_X8Y156_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X7Y156_SLICE_X8Y156_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y156_SLICE_X8Y156_D2 = 1'b1;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_B2 = CLBLM_R_X7Y155_SLICE_X9Y155_BQ;
  assign CLBLM_R_X7Y156_SLICE_X8Y156_D3 = CLBLM_R_X7Y156_SLICE_X8Y156_DQ;
  assign CLBLM_R_X7Y156_SLICE_X8Y156_D4 = CLBLL_L_X4Y147_SLICE_X4Y147_BO6;
  assign CLBLM_R_X7Y156_SLICE_X8Y156_D5 = CLBLM_L_X8Y159_SLICE_X10Y159_AQ;
  assign CLBLM_R_X7Y156_SLICE_X8Y156_D6 = CLBLM_R_X7Y147_SLICE_X9Y147_A5Q;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y155_SLICE_X9Y155_B5 = CLBLM_R_X7Y158_SLICE_X8Y158_CO5;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A6 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_D1 = CLBLM_R_X13Y156_SLICE_X18Y156_AQ;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B3 = 1'b1;
  assign RIOB33_X105Y185_IOB_X1Y186_O = CLBLM_R_X13Y154_SLICE_X18Y154_AQ;
  assign RIOB33_X105Y185_IOB_X1Y185_O = CLBLM_R_X7Y149_SLICE_X9Y149_DO5;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B4 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B5 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B6 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y190_T1 = 1'b1;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_D1 = CLBLM_L_X12Y159_SLICE_X16Y159_BQ;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_D1 = LIOB33_X0Y51_IOB_X0Y52_I;
  assign RIOI3_X105Y189_OLOGIC_X1Y189_T1 = 1'b1;
  assign LIOI3_X0Y191_OLOGIC_X0Y192_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_D1 = CLBLL_L_X52Y126_SLICE_X78Y126_AO6;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_D1 = RIOB33_X105Y147_IOB_X1Y148_I;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_D1 = CLBLM_R_X103Y174_SLICE_X163Y174_AO5;
  assign LIOI3_X0Y191_OLOGIC_X0Y191_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_D1 = CLBLL_L_X4Y151_SLICE_X5Y151_CQ;
  assign RIOI3_X105Y175_OLOGIC_X1Y176_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_T1 = 1'b1;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_D1 = CLBLM_R_X13Y157_SLICE_X18Y157_AO5;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign RIOI3_X105Y175_OLOGIC_X1Y175_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_D1 = CLBLM_R_X11Y156_SLICE_X15Y156_BQ;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y188_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_D1 = CLBLM_L_X12Y155_SLICE_X16Y155_AQ;
  assign LIOB33_X0Y101_IOB_X0Y102_O = CLBLL_L_X2Y139_SLICE_X0Y139_AO5;
  assign LIOB33_X0Y101_IOB_X0Y101_O = CLBLL_L_X2Y139_SLICE_X0Y139_AO6;
  assign RIOI3_TBYTETERM_X105Y187_OLOGIC_X1Y187_T1 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A1 = CLBLL_L_X4Y149_SLICE_X5Y149_CO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A2 = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A3 = CLBLM_R_X3Y150_SLICE_X3Y150_AQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A4 = CLBLM_R_X11Y154_SLICE_X15Y154_AQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_A6 = CLBLM_R_X3Y151_SLICE_X3Y151_AO5;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B1 = CLBLL_L_X4Y149_SLICE_X5Y149_CO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B2 = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B3 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B5 = CLBLM_L_X10Y148_SLICE_X12Y148_AQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_B6 = CLBLM_R_X3Y151_SLICE_X3Y151_AO5;
  assign RIOB33_X105Y187_IOB_X1Y187_O = CLBLM_L_X12Y155_SLICE_X16Y155_AQ;
  assign RIOB33_X105Y187_IOB_X1Y188_O = CLBLM_R_X11Y156_SLICE_X15Y156_BQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C1 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C2 = CLBLM_R_X3Y150_SLICE_X3Y150_CQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C3 = CLBLM_R_X3Y150_SLICE_X2Y150_BO5;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C4 = CLBLL_L_X4Y149_SLICE_X4Y149_DO6;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_C6 = CLBLL_L_X4Y149_SLICE_X4Y149_AQ;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOB33_X0Y153_IOB_X0Y154_O = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D1 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D2 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D3 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D4 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D5 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X3Y150_D6 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A1 = CLBLM_R_X3Y150_SLICE_X2Y150_BO5;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A3 = CLBLM_R_X3Y150_SLICE_X2Y150_AQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A4 = CLBLL_L_X4Y149_SLICE_X4Y149_DO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A5 = CLBLM_L_X12Y153_SLICE_X17Y153_CQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_A6 = CLBLM_R_X3Y150_SLICE_X3Y150_CQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_AX = CLBLM_R_X3Y150_SLICE_X2Y150_BO6;
  assign LIOB33_X0Y153_IOB_X0Y153_O = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B1 = CLBLL_L_X4Y149_SLICE_X4Y149_DO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B2 = CLBLM_R_X3Y150_SLICE_X2Y150_A5Q;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B4 = CLBLM_R_X3Y151_SLICE_X2Y151_BQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B5 = CLBLM_L_X8Y147_SLICE_X11Y147_CO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_B6 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C2 = CLBLM_R_X3Y152_SLICE_X2Y152_AO5;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C3 = CLBLL_L_X4Y157_SLICE_X4Y157_CO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C4 = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_C6 = CLBLM_R_X3Y151_SLICE_X2Y151_BQ;
  assign CLBLM_L_X12Y157_SLICE_X17Y157_C1 = CLBLM_R_X7Y157_SLICE_X9Y157_CQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D1 = CLBLM_L_X8Y147_SLICE_X11Y147_CO6;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D2 = 1'b1;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D3 = CLBLM_R_X3Y150_SLICE_X2Y150_AQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D4 = CLBLM_R_X3Y150_SLICE_X3Y150_CQ;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D5 = CLBLM_R_X3Y150_SLICE_X2Y150_A5Q;
  assign CLBLM_R_X3Y150_SLICE_X2Y150_D6 = 1'b1;
  assign LIOI3_X0Y71_ILOGIC_X0Y72_D = LIOB33_X0Y71_IOB_X0Y72_I;
  assign LIOI3_X0Y71_ILOGIC_X0Y71_D = LIOB33_X0Y71_IOB_X0Y71_I;
  assign CLBLM_L_X12Y157_SLICE_X17Y157_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign RIOI3_X105Y115_ILOGIC_X1Y116_D = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y115_ILOGIC_X1Y115_D = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_L_X12Y157_SLICE_X17Y157_D3 = CLBLM_R_X11Y158_SLICE_X15Y158_DO6;
  assign CLBLM_L_X12Y157_SLICE_X17Y157_D4 = 1'b1;
  assign LIOB33_X0Y141_IOB_X0Y142_O = LIOB33_X0Y53_IOB_X0Y54_I;
  assign LIOB33_X0Y141_IOB_X0Y141_O = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign LIOB33_X0Y103_IOB_X0Y104_O = CLBLL_L_X2Y139_SLICE_X0Y139_BO5;
  assign LIOB33_X0Y103_IOB_X0Y103_O = CLBLL_L_X2Y139_SLICE_X0Y139_BO6;
  assign CLBLM_L_X10Y159_SLICE_X13Y159_C4 = CLBLM_L_X8Y156_SLICE_X11Y156_DO6;
  assign CLBLM_L_X10Y159_SLICE_X13Y159_C5 = CLBLM_L_X8Y157_SLICE_X11Y157_DO6;
  assign CLBLM_L_X10Y159_SLICE_X13Y159_C6 = CLBLM_L_X10Y159_SLICE_X13Y159_BO6;
  assign CLBLM_L_X12Y157_SLICE_X16Y157_B4 = CLBLM_R_X11Y159_SLICE_X15Y159_DO5;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_D1 = CLBLM_R_X13Y156_SLICE_X19Y156_AQ;
  assign RIOB33_X105Y189_IOB_X1Y190_O = CLBLM_R_X13Y156_SLICE_X18Y156_AQ;
  assign RIOB33_X105Y189_IOB_X1Y189_O = CLBLM_L_X12Y159_SLICE_X16Y159_BQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A2 = CLBLM_L_X12Y155_SLICE_X16Y155_CO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A3 = CLBLM_R_X3Y151_SLICE_X3Y151_AQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A4 = CLBLM_R_X5Y151_SLICE_X6Y151_C5Q;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A5 = CLBLL_L_X4Y150_SLICE_X4Y150_DO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_A6 = 1'b1;
  assign CLBLM_L_X12Y157_SLICE_X16Y157_C1 = CLBLM_R_X11Y151_SLICE_X15Y151_BQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B1 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B2 = CLBLM_R_X3Y152_SLICE_X3Y152_AO5;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B3 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B4 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B5 = CLBLL_L_X4Y151_SLICE_X4Y151_D5Q;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_B6 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C1 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C2 = CLBLM_R_X5Y150_SLICE_X7Y150_CQ;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C3 = CLBLM_R_X3Y152_SLICE_X2Y152_CO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C4 = CLBLM_R_X3Y150_SLICE_X2Y150_CO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C5 = CLBLM_R_X3Y152_SLICE_X3Y152_DO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_C6 = CLBLM_R_X3Y151_SLICE_X2Y151_CO5;
  assign CLBLM_L_X10Y159_SLICE_X13Y159_D5 = CLBLM_L_X8Y157_SLICE_X11Y157_DO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y159_SLICE_X13Y159_D6 = CLBLM_L_X10Y159_SLICE_X13Y159_BO6;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D1 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D2 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D3 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D4 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D5 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X3Y151_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y193_OLOGIC_X1Y194_T1 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A2 = CLBLM_R_X3Y151_SLICE_X2Y151_BQ;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A3 = CLBLM_R_X3Y150_SLICE_X3Y150_CQ;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A4 = CLBLM_R_X3Y150_SLICE_X2Y150_A5Q;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A5 = CLBLM_R_X3Y150_SLICE_X2Y150_AQ;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_A6 = 1'b1;
  assign CLBLM_L_X12Y157_SLICE_X16Y157_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B1 = CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B2 = CLBLM_R_X3Y151_SLICE_X2Y151_BQ;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B3 = CLBLL_L_X4Y149_SLICE_X4Y149_DO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B4 = CLBLM_R_X3Y150_SLICE_X2Y150_DO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_B6 = CLBLM_R_X3Y151_SLICE_X2Y151_AO5;
  assign LIOI3_X0Y155_OLOGIC_X0Y156_D1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C2 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X16Y156_SLICE_X23Y156_A1 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X23Y156_A2 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X23Y156_A3 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X23Y156_A4 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X23Y156_A5 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X23Y156_A6 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C5 = CLBLL_L_X4Y157_SLICE_X4Y157_CO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_C6 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X23Y156_B1 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X23Y156_B2 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X23Y156_B3 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X23Y156_B4 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X23Y156_B5 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X23Y156_B6 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D1 = CLBLM_R_X3Y150_SLICE_X2Y150_AQ;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D2 = CLBLL_L_X2Y154_SLICE_X1Y154_AO5;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A1 = CLBLM_R_X11Y146_SLICE_X15Y146_DO5;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A2 = CLBLM_R_X7Y148_SLICE_X9Y148_CO5;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A3 = CLBLM_L_X10Y145_SLICE_X13Y145_CQ;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A4 = CLBLM_L_X10Y145_SLICE_X13Y145_BQ;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A5 = CLBLM_R_X7Y146_SLICE_X8Y146_BO6;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_A6 = CLBLM_R_X7Y146_SLICE_X9Y146_BO6;
  assign CLBLM_L_X16Y156_SLICE_X23Y156_C1 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X23Y156_C2 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X23Y156_C3 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B1 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B2 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B3 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B4 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B5 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_B6 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X23Y156_D1 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X23Y156_D2 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C1 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C2 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C3 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C4 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C5 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_C6 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X23Y156_D3 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X23Y156_D4 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X22Y156_A1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_L_X16Y156_SLICE_X22Y156_A2 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X22Y156_A3 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_L_X16Y156_SLICE_X22Y156_A4 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_L_X16Y156_SLICE_X22Y156_A5 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_L_X16Y156_SLICE_X22Y156_A6 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D1 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D2 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D3 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D4 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D5 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X17Y146_D6 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X22Y156_B1 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X22Y156_B2 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X22Y156_B3 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X22Y156_B4 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X22Y156_B5 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A1 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_A2 = CLBLM_L_X12Y146_SLICE_X16Y146_BQ;
  assign CLBLM_L_X16Y156_SLICE_X22Y156_B6 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X22Y156_C1 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X22Y156_C2 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X22Y156_C3 = 1'b1;
  assign CLBLM_L_X10Y159_SLICE_X12Y159_B5 = CLBLM_L_X10Y158_SLICE_X12Y158_BQ;
  assign CLBLM_L_X16Y156_SLICE_X22Y156_C4 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X22Y156_C5 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B1 = 1'b1;
  assign CLBLM_L_X10Y159_SLICE_X12Y159_B6 = CLBLM_R_X11Y159_SLICE_X15Y159_BQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B2 = CLBLM_L_X12Y146_SLICE_X16Y146_BQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B3 = CLBLM_R_X7Y146_SLICE_X8Y146_DO6;
  assign CLBLM_L_X16Y156_SLICE_X22Y156_C6 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_B4 = CLBLM_L_X12Y146_SLICE_X16Y146_CQ;
  assign CLBLM_L_X16Y156_SLICE_X22Y156_D1 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X22Y156_D2 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X22Y156_D3 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C2 = CLBLM_L_X12Y146_SLICE_X16Y146_CQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C3 = CLBLM_L_X12Y146_SLICE_X16Y146_DQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C4 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C5 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_C6 = CLBLM_L_X12Y146_SLICE_X16Y146_AQ;
  assign CLBLM_L_X16Y156_SLICE_X22Y156_D4 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X22Y156_D5 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X22Y156_D6 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D2 = 1'b1;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D3 = CLBLM_L_X12Y146_SLICE_X16Y146_DQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D4 = CLBLM_L_X8Y146_SLICE_X11Y146_CQ;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D5 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_L_X12Y146_SLICE_X16Y146_D6 = CLBLM_R_X11Y150_SLICE_X14Y150_AQ;
  assign CLBLM_L_X10Y159_SLICE_X12Y159_C4 = CLBLM_L_X8Y156_SLICE_X11Y156_DO6;
  assign CLBLM_R_X11Y155_SLICE_X15Y155_B1 = CLBLM_R_X11Y156_SLICE_X14Y156_DO6;
  assign CLBLM_L_X10Y159_SLICE_X12Y159_C5 = CLBLM_L_X8Y159_SLICE_X10Y159_BO6;
  assign CLBLM_R_X11Y155_SLICE_X15Y155_B2 = CLBLM_R_X7Y149_SLICE_X8Y149_DO5;
  assign CLBLM_L_X10Y159_SLICE_X12Y159_C6 = CLBLM_L_X10Y159_SLICE_X12Y159_BO6;
  assign CLBLM_R_X11Y155_SLICE_X15Y155_B3 = CLBLM_L_X8Y155_SLICE_X10Y155_DO6;
  assign CLBLM_R_X11Y155_SLICE_X15Y155_B4 = CLBLM_L_X12Y156_SLICE_X16Y156_DO6;
  assign CLBLM_R_X11Y155_SLICE_X15Y155_B5 = CLBLM_R_X13Y156_SLICE_X18Y156_BO6;
  assign LIOB33_X0Y105_IOB_X0Y106_O = CLBLL_L_X2Y140_SLICE_X0Y140_BO5;
  assign LIOB33_X0Y105_IOB_X0Y105_O = CLBLL_L_X2Y140_SLICE_X0Y140_BO6;
  assign CLBLM_R_X11Y155_SLICE_X15Y155_B6 = CLBLM_L_X10Y159_SLICE_X12Y159_CO6;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE = 1'b1;
  assign CLBLM_R_X11Y155_SLICE_X15Y155_C1 = CLBLM_R_X11Y157_SLICE_X15Y157_AQ;
  assign CLBLM_R_X11Y155_SLICE_X15Y155_C2 = CLBLM_R_X3Y157_SLICE_X2Y157_AO5;
  assign CLBLM_R_X11Y155_SLICE_X15Y155_C3 = CLBLM_L_X12Y155_SLICE_X16Y155_BO5;
  assign RIOB33_X105Y191_IOB_X1Y192_O = CLBLM_R_X13Y153_SLICE_X19Y153_BQ;
  assign RIOB33_X105Y191_IOB_X1Y191_O = CLBLM_L_X12Y156_SLICE_X16Y156_BQ;
  assign CLBLM_R_X11Y155_SLICE_X15Y155_C4 = CLBLM_L_X12Y155_SLICE_X16Y155_DO6;
  assign CLBLM_R_X11Y155_SLICE_X15Y155_C5 = CLBLM_R_X5Y149_SLICE_X7Y149_AQ;
  assign CLBLM_R_X11Y155_SLICE_X15Y155_C6 = CLBLM_R_X11Y155_SLICE_X15Y155_DO6;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_D1 = LIOB33_X0Y69_IOB_X0Y69_I;
  assign CLBLM_R_X11Y155_SLICE_X15Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOI3_X0Y195_OLOGIC_X0Y196_T1 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_D1 = CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A1 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A2 = CLBLM_R_X3Y152_SLICE_X2Y152_DO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A3 = CLBLL_L_X4Y158_SLICE_X5Y158_AQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A4 = CLBLM_R_X3Y152_SLICE_X3Y152_BO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_A6 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_T1 = 1'b1;
  assign LIOI3_X0Y195_OLOGIC_X0Y195_D1 = LIOB33_X0Y63_IOB_X0Y64_I;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B2 = CLBLL_L_X4Y154_SLICE_X5Y154_BO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B3 = CLBLM_R_X5Y155_SLICE_X6Y155_DO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B4 = CLBLL_L_X4Y153_SLICE_X4Y153_BO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B5 = CLBLL_L_X4Y154_SLICE_X5Y154_CO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_B6 = 1'b1;
  assign CLBLM_R_X11Y155_SLICE_X15Y155_D1 = CLBLM_L_X12Y155_SLICE_X17Y155_BQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_D1 = CLBLM_R_X5Y146_SLICE_X6Y146_A5Q;
  assign CLBLM_R_X11Y155_SLICE_X15Y155_D2 = CLBLM_L_X12Y153_SLICE_X16Y153_DO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C1 = CLBLL_L_X4Y155_SLICE_X4Y155_BQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C2 = CLBLM_R_X3Y152_SLICE_X2Y152_AO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C3 = CLBLL_L_X2Y155_SLICE_X1Y155_CO5;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C5 = CLBLL_L_X4Y157_SLICE_X4Y157_CO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_C6 = CLBLM_R_X3Y150_SLICE_X3Y150_CQ;
  assign CLBLM_R_X11Y155_SLICE_X15Y155_D3 = CLBLM_L_X8Y157_SLICE_X11Y157_DO6;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_T1 = 1'b1;
  assign CLBLM_R_X11Y155_SLICE_X15Y155_D4 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_T1 = 1'b1;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_AO6;
  assign CLBLM_R_X11Y155_SLICE_X15Y155_D5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D1 = CLBLM_R_X3Y152_SLICE_X3Y152_AO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D2 = CLBLM_R_X3Y152_SLICE_X2Y152_AO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D3 = CLBLL_L_X4Y157_SLICE_X4Y157_CO6;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D4 = CLBLL_L_X4Y149_SLICE_X4Y149_AQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D5 = CLBLL_L_X4Y151_SLICE_X4Y151_DQ;
  assign CLBLM_R_X3Y152_SLICE_X3Y152_D6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X11Y155_SLICE_X15Y155_D6 = CLBLM_R_X11Y155_SLICE_X14Y155_BQ;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_D1 = RIOB33_X105Y115_IOB_X1Y116_I;
  assign RIOI3_X105Y177_OLOGIC_X1Y177_T1 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A3 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A5 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y158_T1 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B1 = CLBLL_L_X4Y157_SLICE_X4Y157_CO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B2 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B4 = CLBLL_L_X2Y155_SLICE_X1Y155_CO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B5 = CLBLL_L_X4Y151_SLICE_X4Y151_D5Q;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_B6 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_D1 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C1 = RIOB33_X105Y117_IOB_X1Y117_I;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C2 = CLBLM_R_X3Y158_SLICE_X2Y158_AO5;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C3 = CLBLL_L_X4Y157_SLICE_X4Y157_CO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C4 = CLBLL_L_X2Y155_SLICE_X1Y155_CO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C5 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_C6 = CLBLM_R_X3Y156_SLICE_X3Y156_AO6;
  assign LIOI3_TBYTESRC_X0Y157_OLOGIC_X0Y157_T1 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D1 = CLBLL_L_X4Y153_SLICE_X4Y153_AO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D2 = CLBLL_L_X4Y154_SLICE_X4Y154_BO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D3 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D4 = 1'b1;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D5 = CLBLM_R_X3Y156_SLICE_X2Y156_DO6;
  assign CLBLM_R_X3Y152_SLICE_X2Y152_D6 = CLBLM_R_X3Y155_SLICE_X2Y155_BO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A1 = CLBLM_L_X12Y147_SLICE_X17Y147_DO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A2 = CLBLM_R_X11Y147_SLICE_X15Y147_AO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A3 = CLBLM_L_X12Y148_SLICE_X17Y148_DO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A4 = CLBLM_L_X12Y147_SLICE_X17Y147_BO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A5 = CLBLM_L_X12Y148_SLICE_X16Y148_CO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_A6 = CLBLM_L_X12Y147_SLICE_X17Y147_CO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B1 = CLBLM_R_X7Y146_SLICE_X8Y146_BO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B2 = CLBLM_L_X12Y147_SLICE_X16Y147_BO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B3 = CLBLM_L_X10Y150_SLICE_X13Y150_C5Q;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B4 = CLBLM_R_X7Y148_SLICE_X9Y148_CO5;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B5 = CLBLM_R_X11Y153_SLICE_X15Y153_DQ;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_B6 = CLBLM_R_X7Y146_SLICE_X9Y146_BO6;
  assign CLBLM_R_X13Y153_SLICE_X18Y153_D4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C1 = CLBLM_R_X13Y147_SLICE_X18Y147_AO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C2 = CLBLM_R_X7Y146_SLICE_X8Y146_BO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C3 = CLBLM_L_X12Y147_SLICE_X16Y147_BO5;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C4 = CLBLM_R_X3Y154_SLICE_X2Y154_AO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C5 = CLBLM_L_X12Y149_SLICE_X16Y149_B5Q;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_C6 = CLBLM_L_X10Y149_SLICE_X12Y149_CQ;
  assign CLBLM_R_X13Y153_SLICE_X18Y153_D5 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X13Y153_SLICE_X18Y153_D6 = CLBLM_R_X13Y157_SLICE_X18Y157_AQ;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_C4 = CLBLM_L_X10Y153_SLICE_X12Y153_BQ;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D1 = CLBLM_R_X13Y147_SLICE_X18Y147_BO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D2 = CLBLM_R_X11Y152_SLICE_X14Y152_BQ;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D3 = CLBLM_L_X12Y154_SLICE_X16Y154_A5Q;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D4 = CLBLM_R_X3Y154_SLICE_X2Y154_AO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D5 = CLBLM_R_X7Y146_SLICE_X8Y146_BO6;
  assign CLBLM_L_X12Y147_SLICE_X17Y147_D6 = CLBLM_R_X13Y147_SLICE_X18Y147_DO6;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_C5 = 1'b1;
  assign CLBLM_R_X11Y155_SLICE_X14Y155_B1 = CLBLM_L_X10Y154_SLICE_X13Y154_DQ;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_C6 = CLBLM_R_X5Y152_SLICE_X6Y152_CO5;
  assign CLBLM_R_X11Y155_SLICE_X14Y155_B2 = CLBLM_R_X11Y155_SLICE_X14Y155_BQ;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A1 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A3 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A4 = CLBLM_L_X10Y150_SLICE_X12Y150_A5Q;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A5 = 1'b1;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_A6 = CLBLM_L_X12Y147_SLICE_X16Y147_CO6;
  assign CLBLM_R_X11Y155_SLICE_X14Y155_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y155_SLICE_X14Y155_B4 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B1 = CLBLM_L_X10Y146_SLICE_X12Y146_C5Q;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B2 = CLBLM_L_X10Y145_SLICE_X13Y145_BQ;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B3 = CLBLM_L_X10Y146_SLICE_X12Y146_CQ;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B4 = CLBLM_L_X10Y145_SLICE_X13Y145_CQ;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B5 = CLBLM_R_X11Y150_SLICE_X14Y150_AQ;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_B6 = 1'b1;
  assign CLBLM_R_X11Y155_SLICE_X14Y155_B5 = CLBLM_L_X12Y155_SLICE_X17Y155_BQ;
  assign CLBLM_R_X11Y155_SLICE_X14Y155_B6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C1 = CLBLM_L_X12Y153_SLICE_X17Y153_CQ;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C2 = CLBLM_L_X12Y147_SLICE_X16Y147_AQ;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C3 = CLBLM_R_X13Y147_SLICE_X18Y147_AO5;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C4 = CLBLM_L_X8Y148_SLICE_X11Y148_B5Q;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C5 = CLBLM_R_X13Y147_SLICE_X18Y147_BO5;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_C6 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D1 = CLBLM_R_X11Y150_SLICE_X14Y150_AQ;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D2 = CLBLM_L_X10Y147_SLICE_X12Y147_CQ;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D3 = CLBLM_L_X12Y146_SLICE_X16Y146_DQ;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D4 = CLBLM_R_X13Y153_SLICE_X19Y153_CQ;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D5 = CLBLM_L_X12Y153_SLICE_X17Y153_CQ;
  assign CLBLM_L_X12Y147_SLICE_X16Y147_D6 = CLBLM_L_X10Y145_SLICE_X12Y145_BQ;
  assign CLBLM_R_X11Y155_SLICE_X14Y155_C1 = CLBLM_R_X7Y153_SLICE_X8Y153_AQ;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_D2 = 1'b1;
  assign CLBLM_R_X11Y155_SLICE_X14Y155_C2 = 1'b1;
  assign LIOB33_X0Y107_IOB_X0Y107_O = CLBLM_R_X3Y142_SLICE_X3Y142_CO6;
  assign LIOB33_X0Y107_IOB_X0Y108_O = CLBLM_R_X3Y151_SLICE_X3Y151_BO6;
  assign CLBLM_R_X11Y155_SLICE_X14Y155_C3 = CLBLM_L_X10Y159_SLICE_X12Y159_CO6;
  assign CLBLM_R_X11Y155_SLICE_X14Y155_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_D5 = 1'b1;
  assign CLBLM_R_X11Y155_SLICE_X14Y155_C5 = CLBLM_R_X11Y156_SLICE_X14Y156_DO6;
  assign LIOI3_X0Y73_ILOGIC_X0Y74_D = LIOB33_X0Y73_IOB_X0Y74_I;
  assign CLBLM_R_X7Y157_SLICE_X9Y157_D6 = CLBLM_R_X7Y158_SLICE_X8Y158_BQ;
  assign CLBLM_R_X11Y155_SLICE_X14Y155_C6 = 1'b1;
  assign LIOI3_X0Y73_ILOGIC_X0Y73_D = LIOB33_X0Y73_IOB_X0Y73_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y118_D = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y117_ILOGIC_X1Y117_D = RIOB33_X105Y117_IOB_X1Y117_I;
  assign RIOB33_X105Y193_IOB_X1Y194_O = CLBLM_R_X13Y156_SLICE_X19Y156_AQ;
  assign CLBLM_R_X11Y155_SLICE_X14Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign RIOB33_X105Y193_IOB_X1Y193_O = CLBLM_L_X12Y156_SLICE_X16Y156_AQ;
  assign CLBLM_R_X11Y155_SLICE_X14Y155_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y155_SLICE_X14Y155_D2 = CLBLM_L_X10Y152_SLICE_X12Y152_CO6;
  assign CLBLM_R_X11Y155_SLICE_X14Y155_D3 = CLBLM_R_X11Y155_SLICE_X14Y155_DQ;
  assign CLBLM_R_X11Y155_SLICE_X14Y155_D4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y155_SLICE_X14Y155_D5 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X11Y155_SLICE_X14Y155_D6 = CLBLM_L_X8Y155_SLICE_X11Y155_AQ;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A2 = CLBLL_L_X4Y157_SLICE_X4Y157_CO5;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_A6 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B1 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B2 = CLBLM_R_X3Y155_SLICE_X3Y155_DO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B3 = CLBLL_L_X2Y153_SLICE_X1Y153_BO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B4 = CLBLM_R_X5Y154_SLICE_X6Y154_AQ;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B5 = CLBLM_R_X5Y153_SLICE_X7Y153_AQ;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_B6 = CLBLM_R_X3Y153_SLICE_X3Y153_AO5;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_B6 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C1 = CLBLM_R_X5Y154_SLICE_X6Y154_AQ;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C2 = CLBLL_L_X2Y153_SLICE_X0Y153_AO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C3 = CLBLM_R_X3Y153_SLICE_X2Y153_BO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C4 = CLBLM_R_X3Y153_SLICE_X3Y153_AO5;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_C6 = CLBLM_R_X5Y153_SLICE_X7Y153_AQ;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D1 = CLBLM_R_X3Y153_SLICE_X3Y153_AO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D2 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D3 = CLBLM_R_X11Y152_SLICE_X14Y152_AQ;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D4 = CLBLM_R_X3Y152_SLICE_X3Y152_CO6;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D5 = LIOB33_X0Y61_IOB_X0Y61_I;
  assign CLBLM_R_X3Y153_SLICE_X3Y153_D6 = CLBLL_L_X2Y153_SLICE_X1Y153_AO5;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_D1 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A1 = CLBLL_L_X4Y157_SLICE_X4Y157_CO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A2 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_A6 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B1 = CLBLM_R_X3Y158_SLICE_X2Y158_AO5;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B2 = CLBLM_R_X3Y156_SLICE_X3Y156_AO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B3 = RIOB33_X105Y115_IOB_X1Y115_I;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B4 = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B5 = CLBLL_L_X4Y157_SLICE_X4Y157_CO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_B6 = CLBLM_R_X3Y153_SLICE_X2Y153_AO5;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_C4 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_C5 = CLBLM_R_X7Y159_SLICE_X8Y159_BO5;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C5 = CLBLM_R_X3Y158_SLICE_X2Y158_AO5;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_C6 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_C6 = 1'b1;
  assign LIOI3_X0Y53_ILOGIC_X0Y54_D = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D1 = CLBLM_R_X3Y152_SLICE_X2Y152_BO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D2 = CLBLM_L_X8Y154_SLICE_X11Y154_AQ;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D3 = CLBLM_R_X3Y153_SLICE_X3Y153_AO6;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D4 = CLBLL_L_X4Y152_SLICE_X5Y152_CQ;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D5 = 1'b1;
  assign CLBLM_R_X3Y153_SLICE_X2Y153_D6 = CLBLM_R_X3Y151_SLICE_X2Y151_CO6;
  assign LIOI3_X0Y53_ILOGIC_X0Y53_D = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A1 = CLBLM_R_X13Y149_SLICE_X19Y149_A5Q;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A2 = CLBLM_R_X11Y148_SLICE_X15Y148_CO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A3 = CLBLM_R_X13Y149_SLICE_X18Y149_A5Q;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A4 = CLBLM_L_X12Y148_SLICE_X17Y148_BO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A5 = CLBLM_R_X11Y148_SLICE_X15Y148_DO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_A6 = CLBLM_L_X12Y148_SLICE_X17Y148_CO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B1 = CLBLM_R_X13Y148_SLICE_X18Y148_AO5;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B2 = CLBLM_L_X12Y149_SLICE_X17Y149_CO5;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B3 = CLBLM_R_X3Y154_SLICE_X2Y154_AO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B4 = CLBLM_L_X12Y150_SLICE_X17Y150_BQ;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B5 = CLBLM_R_X7Y146_SLICE_X8Y146_BO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_B6 = CLBLM_L_X12Y157_SLICE_X17Y157_A5Q;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C1 = CLBLM_R_X7Y146_SLICE_X8Y146_BO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C2 = CLBLM_R_X7Y148_SLICE_X9Y148_CO5;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C3 = CLBLM_R_X7Y153_SLICE_X8Y153_DO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C4 = CLBLM_R_X13Y152_SLICE_X18Y152_DO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C5 = CLBLM_R_X7Y146_SLICE_X9Y146_BO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_C6 = CLBLM_L_X12Y146_SLICE_X16Y146_BQ;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D1 = CLBLM_R_X7Y146_SLICE_X8Y146_BO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D2 = CLBLM_L_X12Y149_SLICE_X17Y149_CO5;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D3 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D4 = CLBLM_L_X12Y157_SLICE_X17Y157_A5Q;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D5 = CLBLM_R_X7Y146_SLICE_X9Y146_BO6;
  assign CLBLM_L_X12Y148_SLICE_X17Y148_D6 = CLBLM_R_X7Y148_SLICE_X9Y148_CO5;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_D2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_D3 = CLBLM_R_X7Y157_SLICE_X8Y157_DQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A1 = CLBLM_L_X10Y146_SLICE_X12Y146_C5Q;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A2 = CLBLM_L_X12Y153_SLICE_X17Y153_CQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A3 = CLBLM_L_X10Y145_SLICE_X13Y145_CQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A4 = CLBLM_L_X10Y145_SLICE_X13Y145_BQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A5 = CLBLM_L_X10Y146_SLICE_X12Y146_CQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_A6 = 1'b1;
  assign CLBLM_R_X7Y157_SLICE_X8Y157_D5 = CLBLM_R_X5Y157_SLICE_X7Y157_DQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B1 = CLBLM_L_X12Y149_SLICE_X17Y149_BO5;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B2 = CLBLM_L_X12Y146_SLICE_X16Y146_BQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B3 = CLBLM_L_X12Y149_SLICE_X17Y149_AQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B4 = CLBLM_L_X10Y145_SLICE_X12Y145_CQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B5 = CLBLM_R_X13Y149_SLICE_X18Y149_BQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_B6 = CLBLM_L_X12Y146_SLICE_X16Y146_CQ;
  assign RIOI3_X105Y177_OLOGIC_X1Y178_D1 = CLBLM_R_X103Y177_SLICE_X163Y177_AO5;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C1 = CLBLM_R_X7Y146_SLICE_X8Y146_BO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C2 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C3 = CLBLM_R_X7Y146_SLICE_X9Y146_BO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C4 = CLBLM_L_X12Y148_SLICE_X16Y148_AO5;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C5 = CLBLM_L_X8Y148_SLICE_X11Y148_B5Q;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_C6 = CLBLM_R_X7Y148_SLICE_X9Y148_CO5;
  assign LIOB33_X0Y109_IOB_X0Y109_O = CLBLM_R_X3Y142_SLICE_X3Y142_DO6;
  assign LIOB33_X0Y109_IOB_X0Y110_O = CLBLM_R_X3Y142_SLICE_X3Y142_BO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D1 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D2 = CLBLM_R_X13Y149_SLICE_X19Y149_CQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D3 = CLBLM_R_X13Y149_SLICE_X18Y149_AQ;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D4 = CLBLM_L_X12Y147_SLICE_X16Y147_DO6;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D5 = 1'b1;
  assign CLBLM_L_X12Y148_SLICE_X16Y148_D6 = CLBLM_L_X12Y148_SLICE_X16Y148_BO6;
  assign RIOB33_X105Y195_IOB_X1Y196_O = CLBLM_L_X12Y159_SLICE_X16Y159_AQ;
  assign RIOB33_X105Y195_IOB_X1Y195_O = CLBLM_R_X13Y157_SLICE_X18Y157_AQ;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_A1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_A3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_A4 = CLBLL_L_X4Y157_SLICE_X4Y157_CO5;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_A5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_A6 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_B1 = CLBLL_L_X4Y156_SLICE_X4Y156_BO5;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_B2 = CLBLM_R_X3Y155_SLICE_X2Y155_DO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_B3 = CLBLM_R_X3Y157_SLICE_X2Y157_CO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_B4 = CLBLL_L_X2Y154_SLICE_X1Y154_AO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_B5 = CLBLM_R_X3Y154_SLICE_X3Y154_AO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_B6 = CLBLL_L_X2Y155_SLICE_X1Y155_BO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_C1 = CLBLM_R_X3Y155_SLICE_X2Y155_CO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_C2 = CLBLM_R_X3Y155_SLICE_X2Y155_DO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_C3 = CLBLL_L_X4Y156_SLICE_X4Y156_BO5;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_C4 = CLBLM_R_X3Y153_SLICE_X3Y153_AO5;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_C5 = CLBLL_L_X2Y155_SLICE_X1Y155_BO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_C6 = CLBLL_L_X2Y154_SLICE_X1Y154_AO6;
  assign LIOI3_X0Y155_OLOGIC_X0Y155_T1 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_D1 = CLBLM_R_X3Y154_SLICE_X3Y154_AO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_D2 = CLBLL_L_X2Y155_SLICE_X1Y155_BO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_D3 = CLBLM_R_X3Y157_SLICE_X2Y157_CO6;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_D4 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_D5 = CLBLL_L_X4Y156_SLICE_X4Y156_BO5;
  assign CLBLM_R_X3Y154_SLICE_X3Y154_D6 = CLBLL_L_X2Y154_SLICE_X1Y154_AO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_A1 = CLBLL_L_X4Y154_SLICE_X5Y154_CO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_A2 = CLBLL_L_X4Y154_SLICE_X4Y154_AO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_A3 = CLBLL_L_X4Y154_SLICE_X4Y154_BO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_A4 = CLBLM_R_X3Y156_SLICE_X3Y156_BO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_A5 = CLBLL_L_X4Y153_SLICE_X4Y153_AO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_A6 = CLBLL_L_X4Y154_SLICE_X5Y154_BO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C5 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_B1 = CLBLL_L_X2Y155_SLICE_X1Y155_CO5;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_B2 = CLBLL_L_X2Y155_SLICE_X1Y155_CO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_B3 = CLBLL_L_X4Y152_SLICE_X5Y152_CQ;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_B4 = CLBLM_R_X3Y151_SLICE_X3Y151_BO5;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_B5 = CLBLL_L_X4Y157_SLICE_X4Y157_CO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_B6 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_C1 = CLBLL_L_X4Y157_SLICE_X4Y157_CO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_C2 = CLBLM_R_X3Y156_SLICE_X3Y156_AO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_C3 = CLBLL_L_X2Y155_SLICE_X1Y155_CO5;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_C4 = CLBLM_R_X3Y158_SLICE_X2Y158_AO5;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_C5 = RIOB33_X105Y113_IOB_X1Y114_I;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_C6 = CLBLM_R_X3Y150_SLICE_X2Y150_A5Q;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C6 = 1'b1;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_D1 = CLBLM_R_X3Y152_SLICE_X3Y152_AO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_D2 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_D3 = CLBLL_L_X4Y155_SLICE_X5Y155_AQ;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_D4 = CLBLM_R_X3Y154_SLICE_X2Y154_CO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_D5 = CLBLM_R_X3Y155_SLICE_X2Y155_DO6;
  assign CLBLM_R_X3Y154_SLICE_X2Y154_D6 = CLBLL_L_X2Y153_SLICE_X1Y153_AO5;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_D1 = LIOB33_X0Y73_IOB_X0Y73_I;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A1 = CLBLM_L_X12Y157_SLICE_X17Y157_CQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A2 = CLBLM_L_X12Y146_SLICE_X16Y146_BQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A3 = CLBLM_L_X12Y149_SLICE_X17Y149_AQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A5 = CLBLM_R_X7Y146_SLICE_X8Y146_DO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_A6 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_AX = CLBLM_L_X12Y149_SLICE_X17Y149_BO6;
  assign LIOI3_X0Y197_OLOGIC_X0Y198_T1 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B1 = CLBLM_R_X11Y153_SLICE_X15Y153_DQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B2 = CLBLM_L_X12Y149_SLICE_X17Y149_A5Q;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B3 = CLBLM_R_X7Y150_SLICE_X8Y150_AQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B4 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_B6 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C1 = CLBLM_L_X10Y145_SLICE_X12Y145_BQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C2 = CLBLM_L_X10Y145_SLICE_X13Y145_CQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C3 = CLBLM_L_X10Y146_SLICE_X12Y146_C5Q;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C4 = CLBLM_L_X10Y145_SLICE_X13Y145_BQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C5 = CLBLM_L_X10Y146_SLICE_X12Y146_CQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_C6 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_D1 = LIOB33_X0Y71_IOB_X0Y72_I;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_D1 = CLBLM_R_X13Y154_SLICE_X18Y154_DO6;
  assign LIOI3_X0Y197_OLOGIC_X0Y197_T1 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D1 = CLBLM_L_X12Y146_SLICE_X17Y146_AO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D2 = CLBLM_L_X12Y157_SLICE_X17Y157_A5Q;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D3 = CLBLM_R_X13Y149_SLICE_X19Y149_AQ;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D4 = CLBLM_R_X11Y155_SLICE_X15Y155_BO6;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D5 = CLBLM_L_X12Y149_SLICE_X17Y149_CO5;
  assign CLBLM_L_X12Y149_SLICE_X17Y149_D6 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign LIOB33_X0Y111_IOB_X0Y111_O = 1'b0;
  assign LIOB33_X0Y111_IOB_X0Y112_O = CLBLM_L_X12Y151_SLICE_X16Y151_C5Q;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_D1 = CLBLM_R_X5Y146_SLICE_X6Y146_AQ;
  assign RIOI3_X105Y179_OLOGIC_X1Y180_T1 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A1 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A3 = CLBLM_L_X12Y149_SLICE_X16Y149_AQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A4 = CLBLM_L_X12Y150_SLICE_X16Y150_BQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A5 = CLBLM_L_X12Y147_SLICE_X16Y147_AQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_T1 = 1'b1;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_D1 = CLBLM_L_X12Y159_SLICE_X16Y159_AO5;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B1 = CLBLM_L_X12Y150_SLICE_X16Y150_A5Q;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B2 = CLBLM_R_X13Y149_SLICE_X18Y149_AQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B5 = CLBLM_R_X5Y149_SLICE_X7Y149_BQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_D1 = RIOB33_SING_X105Y149_IOB_X1Y149_I;
  assign RIOI3_X105Y179_OLOGIC_X1Y179_T1 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C2 = CLBLM_L_X12Y151_SLICE_X16Y151_BQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C3 = CLBLM_L_X12Y150_SLICE_X16Y150_BQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C5 = CLBLM_R_X11Y146_SLICE_X14Y146_BQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_C6 = CLBLM_R_X11Y151_SLICE_X15Y151_CO6;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y170_T1 = 1'b1;
  assign RIOB33_X105Y197_IOB_X1Y198_O = CLBLM_L_X16Y156_SLICE_X22Y156_AO5;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOB33_X105Y197_IOB_X1Y197_O = CLBLM_L_X16Y156_SLICE_X22Y156_AO5;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_D1 = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D2 = CLBLM_L_X12Y151_SLICE_X16Y151_BQ;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D3 = 1'b1;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D4 = CLBLM_R_X11Y144_SLICE_X15Y144_A5Q;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y149_SLICE_X16Y149_D6 = CLBLM_R_X11Y151_SLICE_X15Y151_CO6;
  assign LIOI3_TBYTESRC_X0Y169_OLOGIC_X0Y169_T1 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X23Y156_C4 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X23Y156_C5 = 1'b1;
  assign CLBLM_L_X16Y156_SLICE_X23Y156_C6 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_A1 = CLBLM_R_X3Y157_SLICE_X2Y157_CO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_A2 = CLBLL_L_X4Y156_SLICE_X4Y156_BO5;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_A3 = CLBLM_R_X3Y154_SLICE_X3Y154_AO6;
  assign CLBLM_L_X16Y156_SLICE_X23Y156_D5 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_A4 = CLBLL_L_X2Y154_SLICE_X1Y154_AO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_A5 = CLBLL_L_X4Y156_SLICE_X4Y156_CO5;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_A6 = CLBLL_L_X2Y155_SLICE_X1Y155_BO6;
  assign CLBLM_L_X16Y156_SLICE_X23Y156_D6 = 1'b1;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_B1 = CLBLL_L_X2Y155_SLICE_X1Y155_AO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_B2 = CLBLL_L_X2Y154_SLICE_X1Y154_AO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_B3 = CLBLM_R_X3Y155_SLICE_X2Y155_CO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_B4 = CLBLM_R_X3Y155_SLICE_X2Y155_DO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_B5 = CLBLL_L_X4Y156_SLICE_X4Y156_CO5;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_B6 = CLBLL_L_X4Y156_SLICE_X4Y156_BO5;
  assign LIOI3_X0Y75_ILOGIC_X0Y76_D = LIOB33_X0Y75_IOB_X0Y76_I;
  assign LIOI3_X0Y75_ILOGIC_X0Y75_D = LIOB33_X0Y75_IOB_X0Y75_I;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_C1 = CLBLM_R_X3Y154_SLICE_X3Y154_AO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_C2 = CLBLL_L_X4Y157_SLICE_X4Y157_CO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_C3 = CLBLL_L_X4Y157_SLICE_X5Y157_AO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_C4 = CLBLM_R_X3Y152_SLICE_X3Y152_AO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_C5 = CLBLL_L_X4Y156_SLICE_X4Y156_BO5;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_C6 = CLBLL_L_X2Y154_SLICE_X1Y154_AO6;
  assign RIOI3_X105Y121_ILOGIC_X1Y122_D = RIOB33_X105Y121_IOB_X1Y122_I;
  assign RIOI3_X105Y121_ILOGIC_X1Y121_D = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_D1 = CLBLM_R_X3Y157_SLICE_X2Y157_DO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_D2 = CLBLM_R_X3Y155_SLICE_X2Y155_CO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_D3 = CLBLL_L_X4Y156_SLICE_X4Y156_BO5;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_D4 = CLBLL_L_X2Y155_SLICE_X1Y155_BO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_D5 = CLBLM_R_X3Y156_SLICE_X3Y156_DO6;
  assign CLBLM_R_X3Y155_SLICE_X3Y155_D6 = CLBLL_L_X2Y154_SLICE_X1Y154_AO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_A1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_A2 = CLBLL_L_X4Y155_SLICE_X5Y155_AQ;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_A3 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_A4 = CLBLM_R_X3Y156_SLICE_X3Y156_AO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_A5 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_A6 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_B1 = CLBLM_R_X3Y153_SLICE_X2Y153_DO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_B2 = CLBLL_L_X2Y155_SLICE_X1Y155_DO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_B3 = CLBLM_R_X3Y155_SLICE_X3Y155_CO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_B4 = CLBLM_R_X3Y157_SLICE_X3Y157_DO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_B5 = CLBLL_L_X4Y152_SLICE_X5Y152_AQ;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_B6 = CLBLM_R_X3Y157_SLICE_X2Y157_AO5;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_C1 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_C2 = CLBLM_R_X3Y152_SLICE_X3Y152_AO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_C3 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_C4 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_C5 = CLBLL_L_X4Y157_SLICE_X5Y157_AO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_C6 = CLBLL_L_X2Y155_SLICE_X1Y155_CO5;
  assign LIOB33_X0Y143_IOB_X0Y143_O = LIOB33_X0Y55_IOB_X0Y55_I;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_D1 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_D2 = CLBLM_R_X3Y152_SLICE_X3Y152_AO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_D3 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_D4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_D5 = CLBLL_L_X4Y157_SLICE_X5Y157_AO6;
  assign CLBLM_R_X3Y155_SLICE_X2Y155_D6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X12Y158_SLICE_X17Y158_C3 = CLBLM_R_X11Y158_SLICE_X15Y158_CO6;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A1 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A2 = CLBLM_L_X10Y150_SLICE_X12Y150_BO6;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A3 = CLBLM_L_X12Y150_SLICE_X17Y150_AQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A5 = CLBLM_L_X12Y154_SLICE_X17Y154_DQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D3 = 1'b1;
  assign LIOB33_X0Y113_IOB_X0Y113_O = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B1 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B2 = CLBLM_L_X12Y150_SLICE_X17Y150_BQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B3 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B4 = CLBLM_L_X12Y148_SLICE_X17Y148_DO6;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B5 = CLBLM_R_X7Y149_SLICE_X9Y149_BQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOB33_X0Y113_IOB_X0Y114_O = CLBLM_L_X8Y146_SLICE_X10Y146_BQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C1 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C2 = CLBLM_L_X12Y155_SLICE_X17Y155_CQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C3 = CLBLM_L_X12Y154_SLICE_X16Y154_A5Q;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C4 = CLBLM_R_X13Y153_SLICE_X19Y153_CQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C5 = CLBLM_L_X12Y148_SLICE_X16Y148_AO6;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_C6 = CLBLM_L_X10Y146_SLICE_X12Y146_CQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X12Y158_SLICE_X17Y158_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D1 = CLBLM_R_X11Y152_SLICE_X14Y152_BQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D2 = CLBLM_L_X10Y146_SLICE_X12Y146_CQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D3 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D4 = CLBLM_L_X12Y146_SLICE_X16Y146_DQ;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D5 = CLBLM_L_X12Y149_SLICE_X17Y149_CO6;
  assign CLBLM_L_X12Y150_SLICE_X17Y150_D6 = CLBLM_R_X13Y150_SLICE_X18Y150_CQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A2 = CLBLM_R_X13Y149_SLICE_X18Y149_BQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A3 = CLBLM_L_X12Y150_SLICE_X16Y150_AQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A5 = CLBLM_R_X7Y150_SLICE_X9Y150_BO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_A6 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_AX = CLBLM_R_X11Y154_SLICE_X15Y154_CO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B1 = CLBLM_L_X12Y152_SLICE_X16Y152_CQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B2 = CLBLM_L_X12Y150_SLICE_X16Y150_BQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B3 = CLBLM_L_X12Y149_SLICE_X16Y149_CQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_B6 = CLBLM_L_X12Y149_SLICE_X16Y149_DQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C1 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C3 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C4 = CLBLM_L_X8Y153_SLICE_X11Y153_CQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C5 = CLBLM_L_X12Y150_SLICE_X16Y150_DO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_C6 = 1'b1;
  assign CLBLM_L_X12Y158_SLICE_X17Y158_D3 = 1'b1;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X12Y158_SLICE_X17Y158_D4 = CLBLM_R_X11Y159_SLICE_X15Y159_AQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D1 = CLBLM_L_X10Y146_SLICE_X12Y146_CQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D2 = CLBLM_L_X12Y149_SLICE_X17Y149_CO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D3 = CLBLM_L_X8Y155_SLICE_X10Y155_BQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D4 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D5 = CLBLM_L_X12Y150_SLICE_X16Y150_CQ;
  assign CLBLM_L_X12Y150_SLICE_X16Y150_D6 = CLBLM_L_X12Y149_SLICE_X17Y149_A5Q;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A2 = CLBLM_R_X11Y156_SLICE_X15Y156_BQ;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A3 = CLBLM_L_X12Y155_SLICE_X16Y155_AQ;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A5 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_A6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_B6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_C6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X163Y169_D6 = 1'b1;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_A6 = CLBLM_L_X12Y158_SLICE_X16Y158_CO6;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_A6 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_D1 = CLBLL_L_X2Y139_SLICE_X0Y139_BO5;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_B6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_C6 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D1 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D2 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D3 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D4 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D5 = 1'b1;
  assign CLBLM_R_X103Y169_SLICE_X162Y169_D6 = 1'b1;
  assign LIOB33_SING_X0Y100_IOB_X0Y100_O = CLBLL_L_X2Y140_SLICE_X0Y140_AO5;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_A1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_A3 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_A4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_A5 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_A6 = 1'b1;
  assign LIOI3_X0Y103_OLOGIC_X0Y104_T1 = 1'b1;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_B1 = CLBLM_R_X3Y155_SLICE_X3Y155_DO6;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_B2 = CLBLM_R_X3Y155_SLICE_X3Y155_BO6;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_B3 = CLBLM_R_X3Y156_SLICE_X2Y156_AO6;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_B4 = CLBLL_L_X4Y156_SLICE_X5Y156_AO6;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_B5 = CLBLM_R_X3Y156_SLICE_X3Y156_CO6;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_B6 = CLBLM_R_X7Y158_SLICE_X9Y158_DO6;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_C1 = CLBLM_R_X11Y157_SLICE_X15Y157_AQ;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_C1 = CLBLM_R_X3Y157_SLICE_X3Y157_AO6;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_C2 = CLBLL_L_X4Y152_SLICE_X5Y152_AQ;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_C3 = CLBLM_R_X3Y157_SLICE_X2Y157_AO5;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_C4 = CLBLL_L_X4Y156_SLICE_X4Y156_DO6;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_C5 = CLBLM_R_X3Y157_SLICE_X3Y157_BO6;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_C6 = CLBLM_R_X3Y154_SLICE_X2Y154_BO6;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_C2 = CLBLM_L_X12Y158_SLICE_X16Y158_AQ;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_C3 = CLBLM_R_X11Y159_SLICE_X15Y159_AQ;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_D1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_D2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_D3 = CLBLM_L_X16Y156_SLICE_X22Y156_AO6;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_D4 = CLBLM_R_X3Y156_SLICE_X3Y156_AO6;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_D5 = CLBLL_L_X4Y157_SLICE_X4Y157_AO6;
  assign CLBLM_R_X3Y156_SLICE_X3Y156_D6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y78_D = LIOB33_X0Y77_IOB_X0Y78_I;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_A1 = CLBLM_R_X3Y156_SLICE_X2Y156_BO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_A2 = CLBLM_R_X3Y157_SLICE_X2Y157_BO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_A3 = CLBLM_R_X3Y155_SLICE_X2Y155_AO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_A4 = CLBLL_L_X4Y157_SLICE_X5Y157_BO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_A5 = CLBLM_R_X3Y154_SLICE_X2Y154_CO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_A6 = CLBLL_L_X2Y153_SLICE_X1Y153_CO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_B1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_B2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_B3 = CLBLL_L_X4Y157_SLICE_X4Y157_CO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_B4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_B5 = LIOB33_X0Y59_IOB_X0Y59_I;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_B6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOI3_X0Y103_OLOGIC_X0Y103_D1 = CLBLL_L_X2Y139_SLICE_X0Y139_BO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_C1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_C2 = CLBLL_L_X4Y157_SLICE_X4Y157_CO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_C3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_C4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_C5 = LIOB33_X0Y69_IOB_X0Y70_I;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_C6 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign LIOB33_X0Y115_IOB_X0Y115_O = CLBLM_L_X12Y151_SLICE_X16Y151_CQ;
  assign LIOB33_X0Y115_IOB_X0Y116_O = CLBLM_R_X11Y144_SLICE_X15Y144_AQ;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D3 = LIOB33_X0Y57_IOB_X0Y57_I;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D4 = CLBLM_R_X3Y151_SLICE_X2Y151_CO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_D1 = CLBLL_L_X4Y156_SLICE_X5Y156_AO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_D2 = CLBLM_R_X3Y154_SLICE_X2Y154_DO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_D3 = CLBLL_L_X2Y153_SLICE_X1Y153_DO6;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D5 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_D4 = CLBLM_R_X7Y158_SLICE_X9Y158_DO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_D5 = CLBLM_R_X3Y155_SLICE_X3Y155_DO6;
  assign CLBLM_R_X3Y156_SLICE_X2Y156_D6 = CLBLL_L_X4Y157_SLICE_X5Y157_BO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A1 = CLBLM_L_X12Y155_SLICE_X17Y155_CQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A2 = CLBLM_L_X12Y151_SLICE_X17Y151_BQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A3 = CLBLM_R_X5Y152_SLICE_X6Y152_BQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_A6 = 1'b1;
  assign CLBLM_R_X3Y151_SLICE_X2Y151_D6 = CLBLL_L_X2Y153_SLICE_X1Y153_AO5;
  assign CLBLM_R_X13Y154_SLICE_X19Y154_C4 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B1 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B2 = CLBLM_L_X12Y152_SLICE_X16Y152_BQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B4 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_B6 = CLBLM_L_X12Y154_SLICE_X16Y154_A5Q;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_D3 = CLBLM_R_X11Y159_SLICE_X15Y159_AQ;
  assign CLBLM_R_X13Y154_SLICE_X19Y154_C5 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C1 = CLBLM_R_X11Y149_SLICE_X14Y149_BQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C2 = CLBLM_R_X13Y153_SLICE_X19Y153_AQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C3 = CLBLM_R_X13Y151_SLICE_X18Y151_AQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C4 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C5 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_C6 = CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_D4 = CLBLM_L_X12Y159_SLICE_X17Y159_AO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X13Y154_SLICE_X19Y154_C6 = 1'b1;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_O = LIOB33_X0Y61_IOB_X0Y62_I;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_D6 = CLBLM_R_X11Y159_SLICE_X14Y159_AQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D1 = CLBLM_R_X11Y151_SLICE_X15Y151_CO6;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D2 = CLBLM_L_X10Y154_SLICE_X13Y154_BQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D3 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D4 = CLBLM_L_X12Y151_SLICE_X17Y151_BQ;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D5 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X17Y151_D6 = CLBLM_L_X12Y151_SLICE_X16Y151_BQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A1 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A3 = CLBLM_L_X12Y151_SLICE_X16Y151_AQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A5 = CLBLM_L_X12Y149_SLICE_X16Y149_AQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_A6 = CLBLM_R_X11Y157_SLICE_X14Y157_BQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B2 = CLBLM_L_X12Y151_SLICE_X16Y151_BQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B3 = CLBLM_L_X12Y151_SLICE_X17Y151_DO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B4 = CLBLM_L_X12Y152_SLICE_X16Y152_BQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_B6 = CLBLM_L_X10Y154_SLICE_X13Y154_C5Q;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C1 = CLBLM_R_X13Y153_SLICE_X18Y153_BQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C4 = CLBLM_L_X12Y150_SLICE_X17Y150_BQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C5 = CLBLM_R_X11Y151_SLICE_X15Y151_A5Q;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_C6 = 1'b1;
  assign CLBLM_R_X13Y154_SLICE_X19Y154_D2 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D1 = CLBLM_R_X13Y150_SLICE_X19Y150_AQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D2 = CLBLM_L_X12Y153_SLICE_X16Y153_AQ;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D3 = CLBLM_R_X11Y150_SLICE_X15Y150_DO6;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D4 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D5 = 1'b1;
  assign CLBLM_L_X12Y151_SLICE_X16Y151_D6 = CLBLM_R_X11Y151_SLICE_X14Y151_DO6;
  assign CLBLM_R_X13Y154_SLICE_X19Y154_D5 = 1'b1;
  assign CLBLM_R_X13Y154_SLICE_X19Y154_D6 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_D1 = CLBLM_L_X12Y155_SLICE_X17Y155_DO5;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = CLBLM_R_X5Y144_SLICE_X6Y144_AQ;
  assign RIOI3_X105Y183_OLOGIC_X1Y184_T1 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_D1 = CLBLM_L_X12Y155_SLICE_X17Y155_DO6;
  assign LIOB33_SING_X0Y150_IOB_X0Y150_O = LIOB33_X0Y63_IOB_X0Y63_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_D1 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign RIOI3_X105Y183_OLOGIC_X1Y183_T1 = 1'b1;
  assign CLBLM_R_X11Y156_SLICE_X15Y156_C4 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y182_T1 = 1'b1;
  assign CLBLM_R_X11Y156_SLICE_X15Y156_C5 = CLBLM_L_X10Y159_SLICE_X12Y159_DO6;
  assign CLBLM_R_X11Y156_SLICE_X15Y156_C6 = CLBLM_L_X10Y157_SLICE_X12Y157_BQ;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_D1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X11Y156_SLICE_X15Y156_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X13Y154_SLICE_X18Y154_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign LIOI3_TBYTESRC_X0Y181_OLOGIC_X0Y181_T1 = 1'b1;
  assign CLBLM_R_X13Y154_SLICE_X18Y154_B6 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_A1 = CLBLL_L_X2Y155_SLICE_X1Y155_CO6;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_A2 = CLBLM_R_X5Y157_SLICE_X7Y157_BQ;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_A3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_A4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_A5 = CLBLL_L_X2Y155_SLICE_X1Y155_CO5;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_A6 = CLBLM_R_X3Y158_SLICE_X2Y158_AO5;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_B1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_B2 = CLBLL_L_X2Y155_SLICE_X1Y155_CO6;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_B3 = CLBLL_L_X2Y155_SLICE_X1Y155_CO5;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_B4 = CLBLM_R_X3Y158_SLICE_X2Y158_AO5;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_B5 = CLBLM_L_X8Y152_SLICE_X10Y152_CQ;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_B6 = CLBLM_R_X5Y157_SLICE_X7Y157_CQ;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_C1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_C2 = CLBLM_R_X5Y157_SLICE_X7Y157_BQ;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_C3 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_C4 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_C6 = CLBLL_L_X4Y157_SLICE_X4Y157_CO5;
  assign CLBLM_R_X13Y154_SLICE_X18Y154_C1 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X13Y154_SLICE_X18Y154_C2 = CLBLM_R_X13Y154_SLICE_X18Y154_CQ;
  assign CLBLM_R_X13Y154_SLICE_X18Y154_C3 = CLBLM_L_X12Y151_SLICE_X17Y151_AQ;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_D1 = CLBLL_L_X4Y157_SLICE_X4Y157_BO6;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_D2 = CLBLL_L_X4Y157_SLICE_X4Y157_DO6;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_D3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_D4 = CLBLM_R_X3Y157_SLICE_X3Y157_CO6;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_D5 = CLBLM_R_X5Y157_SLICE_X7Y157_CQ;
  assign CLBLM_R_X3Y157_SLICE_X3Y157_D6 = CLBLM_R_X3Y157_SLICE_X2Y157_AO6;
  assign CLBLM_R_X13Y154_SLICE_X18Y154_C4 = CLBLM_R_X7Y152_SLICE_X9Y152_CO6;
  assign LIOB33_X0Y117_IOB_X0Y117_O = CLBLM_R_X5Y147_SLICE_X7Y147_CQ;
  assign CLBLM_R_X11Y156_SLICE_X15Y156_D5 = CLBLM_R_X11Y158_SLICE_X15Y158_BO6;
  assign CLBLM_R_X13Y154_SLICE_X18Y154_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOB33_X0Y117_IOB_X0Y118_O = CLBLM_R_X5Y148_SLICE_X7Y148_BQ;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_A1 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_A3 = CLBLM_R_X3Y158_SLICE_X2Y158_AO6;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_A4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_A5 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_A6 = 1'b1;
  assign CLBLM_R_X11Y156_SLICE_X15Y156_D6 = 1'b1;
  assign CLBLM_R_X13Y154_SLICE_X18Y154_C6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_B1 = CLBLL_L_X4Y157_SLICE_X4Y157_CO6;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_B2 = CLBLL_L_X4Y155_SLICE_X4Y155_AQ;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_B3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_B4 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_B5 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_B6 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_D1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X13Y154_SLICE_X18Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_C1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_C2 = CLBLL_L_X4Y157_SLICE_X4Y157_CO6;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_C3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_C4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_C5 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_C6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_D1 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_D2 = CLBLM_R_X3Y158_SLICE_X2Y158_AO5;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_D3 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_D4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_D5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X3Y157_SLICE_X2Y157_D6 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign LIOB33_SING_X0Y199_IOB_X0Y199_O = LIOB33_X0Y73_IOB_X0Y74_I;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_A1 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_A2 = CLBLM_R_X13Y152_SLICE_X18Y152_AQ;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_A5 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_A6 = CLBLM_R_X7Y151_SLICE_X8Y151_DQ;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_AX = CLBLM_L_X12Y152_SLICE_X17Y152_BO6;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_B1 = CLBLM_L_X12Y151_SLICE_X17Y151_AQ;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_B2 = CLBLL_L_X4Y147_SLICE_X5Y147_AQ;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_B3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_B5 = CLBLM_R_X11Y152_SLICE_X14Y152_CQ;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_B6 = 1'b1;
  assign CLBLM_R_X13Y154_SLICE_X18Y154_D1 = CLBLM_L_X12Y153_SLICE_X17Y153_AQ;
  assign CLBLM_R_X13Y154_SLICE_X18Y154_D2 = 1'b1;
  assign LIOB33_X0Y121_IOB_X0Y122_O = CLBLL_L_X4Y149_SLICE_X5Y149_A5Q;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_C1 = CLBLM_R_X13Y151_SLICE_X18Y151_BQ;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_C2 = CLBLM_R_X11Y153_SLICE_X15Y153_CQ;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_C3 = CLBLM_R_X11Y152_SLICE_X15Y152_CQ;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_C4 = CLBLM_R_X11Y152_SLICE_X15Y152_BQ;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_C5 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_C6 = CLBLM_L_X12Y153_SLICE_X17Y153_BQ;
  assign CLBLM_R_X13Y154_SLICE_X18Y154_D3 = 1'b1;
  assign CLBLM_R_X13Y154_SLICE_X18Y154_D4 = CLBLM_L_X10Y150_SLICE_X13Y150_BQ;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOB33_X0Y121_IOB_X0Y121_O = CLBLM_R_X11Y144_SLICE_X15Y144_A5Q;
  assign LIOI3_X0Y165_OLOGIC_X0Y166_T1 = 1'b1;
  assign CLBLM_R_X13Y154_SLICE_X18Y154_D5 = 1'b1;
  assign CLBLM_R_X7Y158_SLICE_X9Y158_C2 = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_D1 = CLBLM_R_X13Y153_SLICE_X18Y153_AQ;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_D2 = CLBLM_L_X12Y151_SLICE_X17Y151_CO6;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_D3 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_D4 = CLBLM_R_X11Y153_SLICE_X15Y153_CQ;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_D5 = CLBLM_R_X11Y152_SLICE_X15Y152_CQ;
  assign CLBLM_L_X12Y152_SLICE_X17Y152_D6 = CLBLM_L_X10Y153_SLICE_X13Y153_AQ;
  assign CLBLM_R_X7Y158_SLICE_X9Y158_C3 = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X13Y154_SLICE_X18Y154_D6 = CLBLM_R_X11Y152_SLICE_X15Y152_AQ;
  assign CLBLM_R_X7Y158_SLICE_X9Y158_C4 = RIOB33_X105Y133_IOB_X1Y134_I;
  assign LIOI3_X0Y77_ILOGIC_X0Y77_D = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_X105Y123_ILOGIC_X1Y124_D = RIOB33_X105Y123_IOB_X1Y124_I;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_A1 = CLBLM_R_X11Y152_SLICE_X15Y152_CQ;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_A3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_A4 = CLBLM_L_X12Y152_SLICE_X16Y152_CQ;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_A5 = CLBLM_R_X5Y151_SLICE_X6Y151_CQ;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_A6 = 1'b1;
  assign CLBLM_R_X7Y158_SLICE_X9Y158_C5 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X7Y158_SLICE_X9Y158_C6 = CLBLL_L_X4Y157_SLICE_X4Y157_CO5;
  assign RIOI3_X105Y123_ILOGIC_X1Y123_D = RIOB33_X105Y123_IOB_X1Y123_I;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_B2 = CLBLM_L_X10Y150_SLICE_X13Y150_AQ;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_B3 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_B4 = CLBLM_R_X11Y152_SLICE_X15Y152_AQ;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_B5 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_BX = CLBLM_L_X12Y153_SLICE_X17Y153_DO6;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_C1 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_C2 = CLBLM_L_X12Y152_SLICE_X16Y152_CQ;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_C3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_C4 = CLBLM_L_X8Y152_SLICE_X11Y152_CO6;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_C6 = CLBLM_R_X13Y156_SLICE_X18Y156_AQ;
  assign CLBLM_R_X11Y156_SLICE_X14Y156_B5 = CLBLM_R_X11Y152_SLICE_X15Y152_DQ;
  assign CLBLM_R_X11Y156_SLICE_X14Y156_B6 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_D1 = 1'b1;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_D2 = CLBLM_L_X12Y155_SLICE_X16Y155_AO5;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_D3 = CLBLM_L_X12Y152_SLICE_X17Y152_DO6;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_D4 = CLBLM_L_X12Y151_SLICE_X16Y151_DO6;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_D5 = CLBLM_R_X7Y154_SLICE_X9Y154_DO6;
  assign CLBLM_L_X12Y152_SLICE_X16Y152_D6 = CLBLM_R_X13Y152_SLICE_X19Y152_CO6;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_D1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X7Y158_SLICE_X9Y158_D1 = CLBLM_R_X3Y157_SLICE_X2Y157_AO5;
  assign CLBLM_R_X7Y158_SLICE_X9Y158_D2 = CLBLM_R_X5Y151_SLICE_X7Y151_BQ;
  assign LIOB33_X0Y169_IOB_X0Y169_O = RIOB33_X105Y121_IOB_X1Y122_I;
  assign CLBLM_R_X11Y156_SLICE_X14Y156_C4 = CLBLM_L_X12Y157_SLICE_X16Y157_CQ;
  assign CLBLM_R_X7Y158_SLICE_X9Y158_D5 = CLBLL_L_X2Y155_SLICE_X1Y155_BO5;
  assign CLBLM_R_X11Y156_SLICE_X14Y156_C5 = CLBLM_R_X7Y157_SLICE_X9Y157_AQ;
  assign CLBLM_R_X7Y158_SLICE_X9Y158_D6 = CLBLM_R_X7Y156_SLICE_X8Y156_AQ;
  assign CLBLM_R_X11Y156_SLICE_X14Y156_C6 = CLBLM_L_X8Y157_SLICE_X11Y157_DO6;
  assign LIOI3_X0Y165_OLOGIC_X0Y165_T1 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_A1 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_A2 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_A3 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_A4 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_A5 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_A6 = 1'b1;
  assign LIOB33_X0Y119_IOB_X0Y119_O = CLBLM_R_X11Y149_SLICE_X15Y149_AQ;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_B1 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_B2 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_B3 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_B4 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_B5 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_B6 = 1'b1;
  assign LIOB33_X0Y119_IOB_X0Y120_O = CLBLM_L_X12Y149_SLICE_X16Y149_BQ;
  assign CLBLM_R_X7Y158_SLICE_X8Y158_B4 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_C1 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_C2 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_C3 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_C4 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_C5 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_C6 = 1'b1;
  assign CLBLM_R_X7Y158_SLICE_X8Y158_B5 = CLBLM_R_X7Y159_SLICE_X8Y159_AQ;
  assign CLBLM_R_X7Y158_SLICE_X8Y158_B6 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_D1 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_D2 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_D3 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_D4 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_D5 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X3Y158_D6 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_A1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_A2 = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_A3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_A4 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_A5 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_A6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D2 = 1'b1;
  assign CLBLM_R_X7Y158_SLICE_X8Y158_C1 = CLBLM_R_X7Y148_SLICE_X8Y148_BQ;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_B1 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_B2 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_B3 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_B4 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_B5 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_B6 = 1'b1;
  assign CLBLM_R_X7Y158_SLICE_X8Y158_C2 = CLBLM_R_X7Y148_SLICE_X8Y148_AQ;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D5 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_C1 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_C2 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_C3 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_C4 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_C5 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_C6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D6 = 1'b1;
  assign CLBLM_R_X7Y158_SLICE_X8Y158_C6 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_D1 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_D2 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_D3 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_D4 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_D5 = 1'b1;
  assign CLBLM_R_X3Y158_SLICE_X2Y158_D6 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_A1 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_A2 = CLBLM_L_X10Y152_SLICE_X12Y152_DO6;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_A3 = CLBLM_L_X12Y153_SLICE_X17Y153_AQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_A5 = CLBLL_L_X4Y150_SLICE_X5Y150_D5Q;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign RIOI3_X105Y141_ILOGIC_X1Y142_D = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_B1 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_B2 = CLBLM_L_X12Y153_SLICE_X17Y153_BQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_B3 = CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_B4 = CLBLM_L_X10Y157_SLICE_X12Y157_BQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_C1 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_C2 = CLBLM_L_X10Y145_SLICE_X12Y145_CQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_C3 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_C4 = CLBLM_R_X13Y153_SLICE_X18Y153_DQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_C5 = CLBLM_L_X12Y153_SLICE_X17Y153_CQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A2 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign RIOI3_X105Y141_ILOGIC_X1Y141_D = RIOB33_X105Y141_IOB_X1Y141_I;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A3 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_D1 = CLBLM_R_X13Y150_SLICE_X18Y150_CQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_D2 = CLBLM_L_X10Y158_SLICE_X13Y158_BQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_D4 = CLBLM_R_X13Y153_SLICE_X18Y153_DQ;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_D5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y153_SLICE_X17Y153_D6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A5 = 1'b1;
  assign CLBLM_R_X7Y158_SLICE_X8Y158_D1 = CLBLM_L_X8Y157_SLICE_X11Y157_AQ;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_A6 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_A1 = CLBLM_R_X11Y153_SLICE_X15Y153_CQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_A3 = CLBLM_L_X12Y153_SLICE_X16Y153_AQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_A5 = CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_A6 = CLBLL_L_X4Y153_SLICE_X5Y153_AQ;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_A4 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_B2 = CLBLM_R_X7Y151_SLICE_X8Y151_DQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_B3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_B4 = CLBLM_L_X12Y153_SLICE_X17Y153_BQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_B5 = CLBLM_L_X8Y149_SLICE_X11Y149_AQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_B6 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_A5 = 1'b1;
  assign CLBLM_R_X7Y158_SLICE_X8Y158_D5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_A6 = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_C1 = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_C2 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_C3 = RIOB33_X105Y137_IOB_X1Y137_I;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_C4 = CLBLM_L_X8Y153_SLICE_X10Y153_A5Q;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_C5 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_C6 = RIOB33_X105Y127_IOB_X1Y128_I;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_CE = 1'b1;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_D1 = CLBLM_L_X10Y155_SLICE_X12Y155_AQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_D2 = CLBLM_R_X13Y153_SLICE_X18Y153_CQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_D3 = CLBLM_L_X12Y153_SLICE_X17Y153_CQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_D4 = CLBLM_L_X12Y153_SLICE_X16Y153_CO6;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_D5 = CLBLM_R_X7Y152_SLICE_X9Y152_AQ;
  assign CLBLM_L_X12Y153_SLICE_X16Y153_D6 = CLBLM_R_X13Y149_SLICE_X18Y149_A5Q;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B5 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_B1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B6 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_B2 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_B3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A1 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_B4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A3 = CLBLM_R_X13Y156_SLICE_X18Y156_AQ;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A4 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A5 = CLBLM_L_X12Y156_SLICE_X16Y156_BQ;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_B5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_A6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B1 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_B6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_B6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_C6 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_A1 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_A2 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_A3 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_A4 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_A5 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_A6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X163Y172_D1 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_C1 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_B1 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_B2 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_B3 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_B4 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_B5 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_B6 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_C2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C6 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_C3 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_C1 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_C2 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_C3 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_C4 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_C5 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_C6 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_C4 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_C5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_B4 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_C6 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_D1 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_D2 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_D3 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_D4 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_D5 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X19Y147_D6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C3 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_C5 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_A1 = CLBLM_L_X10Y146_SLICE_X12Y146_C5Q;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_A2 = CLBLM_L_X10Y146_SLICE_X12Y146_CQ;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_A3 = CLBLM_L_X10Y145_SLICE_X13Y145_BQ;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_A4 = CLBLM_L_X10Y145_SLICE_X12Y145_CQ;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_A5 = CLBLM_L_X10Y145_SLICE_X13Y145_CQ;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_A6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D1 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D2 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D3 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_B1 = CLBLM_L_X10Y146_SLICE_X12Y146_C5Q;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_B2 = CLBLM_L_X10Y145_SLICE_X13Y145_CQ;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_B3 = CLBLM_L_X10Y145_SLICE_X13Y145_BQ;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_B4 = CLBLM_L_X10Y146_SLICE_X12Y146_CQ;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_B5 = CLBLM_L_X12Y146_SLICE_X16Y146_DQ;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_B6 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D4 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D5 = 1'b1;
  assign CLBLM_R_X103Y172_SLICE_X162Y172_D6 = 1'b1;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_C1 = CLBLM_R_X13Y148_SLICE_X18Y148_BO5;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_C2 = CLBLM_R_X5Y155_SLICE_X6Y155_DO6;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_C3 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_C4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_C5 = CLBLM_R_X13Y155_SLICE_X19Y155_AO6;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_C6 = CLBLM_L_X12Y147_SLICE_X17Y147_AO6;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_D1 = CLBLM_L_X10Y145_SLICE_X13Y145_BQ;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_D2 = CLBLM_L_X10Y145_SLICE_X13Y145_CQ;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_D3 = CLBLM_R_X13Y153_SLICE_X19Y153_CQ;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_D4 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A5 = CLBLM_L_X10Y150_SLICE_X13Y150_B5Q;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_D5 = CLBLM_L_X10Y146_SLICE_X12Y146_C5Q;
  assign CLBLM_R_X13Y147_SLICE_X18Y147_D6 = CLBLM_L_X10Y146_SLICE_X12Y146_CQ;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_D1 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_D2 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_D1 = LIOB33_X0Y53_IOB_X0Y54_I;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_D3 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_D4 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_T1 = 1'b1;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_D5 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_D1 = CLBLM_R_X13Y154_SLICE_X18Y154_AQ;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_D1 = CLBLL_L_X2Y140_SLICE_X0Y140_AO6;
  assign CLBLM_R_X103Y141_SLICE_X162Y141_D6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_D1 = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign RIOI3_X105Y185_OLOGIC_X1Y186_T1 = 1'b1;
  assign LIOI3_X0Y79_OLOGIC_X0Y80_T1 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_T1 = 1'b1;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_D1 = CLBLM_R_X7Y149_SLICE_X9Y149_DO5;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_D1 = LIOB33_X0Y59_IOB_X0Y60_I;
  assign RIOI3_X105Y185_OLOGIC_X1Y185_T1 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B6 = CLBLM_L_X10Y150_SLICE_X13Y150_B5Q;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y194_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_D1 = LIOB33_X0Y55_IOB_X0Y56_I;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_A1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_A2 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_A3 = CLBLL_L_X4Y158_SLICE_X4Y158_AO6;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_A5 = CLBLM_L_X10Y154_SLICE_X13Y154_AQ;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_A6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_AX = CLBLM_L_X12Y154_SLICE_X17Y154_CO6;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_B1 = CLBLM_R_X11Y158_SLICE_X15Y158_BO6;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_B2 = CLBLM_L_X12Y154_SLICE_X17Y154_BQ;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_B3 = CLBLM_L_X12Y154_SLICE_X16Y154_CO5;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_B5 = CLBLM_R_X13Y152_SLICE_X18Y152_CQ;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_B6 = CLBLM_R_X11Y155_SLICE_X15Y155_AQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C1 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C2 = CLBLM_R_X11Y146_SLICE_X14Y146_CQ;
  assign LIOI3_TBYTESRC_X0Y193_OLOGIC_X0Y193_T1 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A1 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A2 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A3 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A4 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A5 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_A6 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_C1 = CLBLM_R_X13Y152_SLICE_X18Y152_A5Q;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_C2 = CLBLM_L_X8Y153_SLICE_X11Y153_BQ;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B1 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B2 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B3 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B4 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B5 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_B6 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_D1 = CLBLM_L_X12Y157_SLICE_X16Y157_AQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C1 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C2 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C3 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C4 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C5 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_C6 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_D3 = CLBLM_L_X12Y154_SLICE_X17Y154_DQ;
  assign CLBLM_L_X12Y154_SLICE_X17Y154_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_A1 = CLBLM_L_X10Y154_SLICE_X12Y154_BO5;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_A2 = CLBLM_R_X13Y154_SLICE_X18Y154_BQ;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_A3 = CLBLM_L_X12Y154_SLICE_X16Y154_AQ;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_A4 = CLBLM_L_X12Y154_SLICE_X16Y154_DO5;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_A6 = CLBLM_L_X12Y154_SLICE_X16Y154_BQ;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D1 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D2 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D3 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D4 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D5 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X13Y144_D6 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_AX = CLBLM_L_X12Y154_SLICE_X16Y154_CO6;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_B1 = CLBLM_L_X10Y154_SLICE_X12Y154_BO5;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_B2 = CLBLM_R_X7Y152_SLICE_X8Y152_A5Q;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_B3 = CLBLM_R_X13Y155_SLICE_X18Y155_AQ;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_B4 = CLBLM_L_X12Y154_SLICE_X16Y154_DO5;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_B5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A1 = CLBLM_L_X8Y153_SLICE_X10Y153_A5Q;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A3 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A4 = CLBLM_L_X10Y147_SLICE_X12Y147_CQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A5 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_A6 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_C1 = CLBLM_L_X12Y152_SLICE_X16Y152_AQ;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_C2 = CLBLM_L_X12Y154_SLICE_X17Y154_A5Q;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_C3 = CLBLM_L_X12Y155_SLICE_X17Y155_AQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B1 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B2 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B3 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B4 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B5 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_B6 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_D1 = CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_D2 = CLBLM_L_X12Y154_SLICE_X16Y154_AQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C1 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C2 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C3 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C4 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C5 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_C6 = 1'b1;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_D3 = CLBLM_R_X11Y154_SLICE_X15Y154_BQ;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_D4 = CLBLM_L_X12Y154_SLICE_X16Y154_BQ;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_D5 = CLBLM_R_X13Y155_SLICE_X18Y155_AQ;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y154_SLICE_X16Y154_D6 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D1 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D2 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D3 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D4 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D5 = 1'b1;
  assign CLBLM_L_X10Y144_SLICE_X12Y144_D6 = 1'b1;
  assign CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_A1 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_A2 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_A3 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_A4 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_A5 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_A6 = 1'b1;
  assign LIOI3_X0Y79_ILOGIC_X0Y79_D = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_B1 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_B2 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_B3 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_B4 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_B5 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_B6 = 1'b1;
  assign RIOI3_X105Y125_ILOGIC_X1Y126_D = RIOB33_X105Y125_IOB_X1Y126_I;
  assign RIOI3_X105Y125_ILOGIC_X1Y125_D = RIOB33_X105Y125_IOB_X1Y125_I;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_C1 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_C2 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_C3 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_C4 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_C5 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_C6 = 1'b1;
  assign LIOB33_X0Y123_IOB_X0Y123_O = CLBLM_L_X8Y146_SLICE_X10Y146_B5Q;
  assign LIOB33_X0Y123_IOB_X0Y124_O = CLBLM_R_X5Y148_SLICE_X7Y148_B5Q;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_D1 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_D2 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_D3 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_D4 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_D5 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X19Y148_D6 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_A1 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_A2 = CLBLM_R_X13Y153_SLICE_X18Y153_CQ;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_A3 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_A4 = CLBLM_R_X13Y148_SLICE_X18Y148_BO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_A6 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_B1 = CLBLM_L_X12Y147_SLICE_X17Y147_AO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_B2 = CLBLM_R_X7Y146_SLICE_X8Y146_DO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_B3 = CLBLM_R_X13Y148_SLICE_X18Y148_AQ;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_B4 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_B5 = CLBLM_R_X13Y148_SLICE_X18Y148_CO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_B6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y119_ILOGIC_X1Y119_D = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_C1 = CLBLM_L_X10Y145_SLICE_X13Y145_BQ;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_C2 = CLBLM_R_X13Y153_SLICE_X18Y153_CQ;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_C3 = CLBLM_L_X10Y145_SLICE_X13Y145_CQ;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_C4 = CLBLM_L_X12Y148_SLICE_X16Y148_DO6;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_C5 = CLBLM_L_X10Y146_SLICE_X12Y146_C5Q;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_C6 = CLBLM_L_X10Y146_SLICE_X12Y146_CQ;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_D1 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_D2 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_D3 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_D4 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_D5 = 1'b1;
  assign CLBLM_R_X13Y148_SLICE_X18Y148_D6 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_A1 = CLBLM_R_X11Y158_SLICE_X15Y158_BO6;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_A3 = CLBLM_L_X12Y155_SLICE_X17Y155_AQ;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_A4 = CLBLM_L_X12Y154_SLICE_X17Y154_CO5;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_A5 = CLBLM_L_X12Y155_SLICE_X16Y155_AQ;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_A6 = CLBLM_L_X12Y155_SLICE_X16Y155_BO5;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_C3 = CLBLM_L_X12Y158_SLICE_X17Y158_AQ;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_B1 = CLBLM_R_X11Y156_SLICE_X14Y156_AQ;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_B2 = CLBLM_L_X12Y155_SLICE_X17Y155_BQ;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_B3 = CLBLM_L_X12Y155_SLICE_X17Y155_CQ;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_B6 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A1 = CLBLM_L_X10Y147_SLICE_X13Y147_CQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A3 = CLBLM_L_X10Y145_SLICE_X13Y145_AQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A5 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_A6 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_C1 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_C2 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_C3 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B1 = CLBLM_L_X10Y145_SLICE_X12Y145_BQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B2 = CLBLM_L_X10Y145_SLICE_X13Y145_BQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B4 = CLBLM_L_X10Y145_SLICE_X13Y145_DO5;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B5 = CLBLM_R_X11Y154_SLICE_X14Y154_DQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_D1 = CLBLM_R_X7Y154_SLICE_X8Y154_AQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C1 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C2 = CLBLM_L_X10Y145_SLICE_X13Y145_CQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C3 = CLBLM_L_X8Y148_SLICE_X11Y148_DO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C4 = CLBLM_R_X11Y146_SLICE_X14Y146_CQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C5 = CLBLM_L_X10Y145_SLICE_X13Y145_DO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_D3 = CLBLM_L_X12Y154_SLICE_X17Y154_DQ;
  assign CLBLM_L_X12Y155_SLICE_X17Y155_D4 = CLBLM_L_X10Y148_SLICE_X13Y148_CQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_A2 = CLBLM_R_X11Y154_SLICE_X15Y154_BQ;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_A3 = CLBLM_R_X13Y155_SLICE_X18Y155_AQ;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_A4 = CLBLM_L_X12Y154_SLICE_X16Y154_AQ;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_A5 = CLBLM_L_X12Y154_SLICE_X16Y154_BQ;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_A6 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D1 = CLBLM_L_X10Y146_SLICE_X12Y146_C5Q;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D2 = CLBLM_L_X10Y145_SLICE_X13Y145_CQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D3 = CLBLM_L_X10Y145_SLICE_X13Y145_BQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D4 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D5 = CLBLM_L_X10Y146_SLICE_X12Y146_CQ;
  assign CLBLM_L_X10Y145_SLICE_X13Y145_D6 = 1'b1;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_AX = CLBLM_L_X12Y151_SLICE_X16Y151_CQ;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_B1 = CLBLM_R_X11Y155_SLICE_X15Y155_AQ;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_B2 = CLBLM_L_X12Y154_SLICE_X17Y154_BQ;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_B3 = CLBLM_L_X12Y154_SLICE_X17Y154_A5Q;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_B4 = CLBLM_L_X8Y153_SLICE_X11Y153_BQ;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_B5 = CLBLM_L_X12Y155_SLICE_X17Y155_AQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A1 = CLBLM_R_X7Y146_SLICE_X9Y146_DO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A3 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A4 = CLBLM_R_X5Y148_SLICE_X7Y148_A5Q;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A5 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_A6 = CLBLM_L_X12Y146_SLICE_X16Y146_AQ;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_C1 = CLBLM_L_X12Y154_SLICE_X16Y154_BQ;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_C2 = CLBLM_R_X11Y154_SLICE_X15Y154_BQ;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_C3 = CLBLM_R_X13Y155_SLICE_X18Y155_AQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B1 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B2 = CLBLM_L_X10Y145_SLICE_X12Y145_BQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B3 = CLBLM_L_X10Y147_SLICE_X12Y147_CQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B5 = CLBLM_R_X11Y144_SLICE_X15Y144_AQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_B6 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_D1 = CLBLM_R_X11Y154_SLICE_X15Y154_BQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C1 = CLBLL_L_X4Y151_SLICE_X5Y151_CQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C2 = CLBLM_L_X10Y145_SLICE_X12Y145_CQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C3 = CLBLM_L_X10Y145_SLICE_X12Y145_BQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C4 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C5 = 1'b1;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_D2 = CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_D3 = CLBLM_R_X13Y155_SLICE_X18Y155_AQ;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_D4 = CLBLM_L_X12Y155_SLICE_X16Y155_AO5;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y155_SLICE_X16Y155_SR = CLBLM_R_X13Y155_SLICE_X18Y155_DO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D1 = CLBLM_L_X10Y146_SLICE_X12Y146_C5Q;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D2 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D3 = CLBLM_L_X10Y146_SLICE_X12Y146_CQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D4 = CLBLM_L_X10Y145_SLICE_X13Y145_CQ;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D5 = CLBLM_L_X8Y148_SLICE_X11Y148_DO6;
  assign CLBLM_L_X10Y145_SLICE_X12Y145_D6 = CLBLM_L_X10Y145_SLICE_X13Y145_BQ;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A2 = CLBLM_R_X13Y153_SLICE_X19Y153_BQ;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A3 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A5 = CLBLM_R_X13Y156_SLICE_X19Y156_AQ;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_A6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_B6 = 1'b1;
  assign LIOI3_X0Y67_ILOGIC_X0Y67_D = LIOB33_X0Y67_IOB_X0Y67_I;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_C6 = 1'b1;
  assign LIOB33_X0Y125_IOB_X0Y125_O = CLBLM_L_X8Y154_SLICE_X10Y154_C5Q;
  assign LIOB33_X0Y125_IOB_X0Y126_O = CLBLL_L_X4Y147_SLICE_X5Y147_AQ;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_A1 = CLBLM_R_X13Y149_SLICE_X18Y149_A5Q;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_A2 = CLBLM_R_X13Y149_SLICE_X19Y149_A5Q;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_A3 = CLBLM_R_X13Y149_SLICE_X19Y149_AQ;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_A4 = CLBLM_R_X13Y149_SLICE_X18Y149_DO6;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_A5 = CLBLM_L_X12Y148_SLICE_X17Y148_AO6;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_A6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D2 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_B1 = CLBLM_R_X13Y149_SLICE_X18Y149_A5Q;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_B2 = CLBLM_R_X13Y149_SLICE_X19Y149_A5Q;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_B3 = CLBLM_R_X13Y149_SLICE_X19Y149_AQ;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_B4 = CLBLM_R_X13Y149_SLICE_X18Y149_DO6;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_B5 = CLBLM_L_X12Y148_SLICE_X17Y148_AO6;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_B6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A2 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_A6 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_C1 = CLBLM_R_X13Y149_SLICE_X18Y149_AQ;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_C2 = CLBLM_R_X13Y149_SLICE_X19Y149_CQ;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_C4 = CLBLM_L_X12Y150_SLICE_X16Y150_A5Q;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_C5 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_C6 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A4 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B2 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_D1 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_D2 = CLBLM_R_X13Y148_SLICE_X18Y148_CO6;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_D3 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_D4 = CLBLM_R_X5Y155_SLICE_X6Y155_DO6;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_D5 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X13Y149_SLICE_X19Y149_D6 = CLBLM_R_X13Y155_SLICE_X19Y155_AO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C1 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C2 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_C5 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_A1 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_B1 = CLBLM_L_X12Y158_SLICE_X16Y158_AQ;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_A2 = CLBLM_R_X13Y149_SLICE_X18Y149_BQ;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_A3 = CLBLM_R_X13Y149_SLICE_X18Y149_AQ;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_A5 = CLBLM_R_X7Y146_SLICE_X8Y146_DO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_A6 = CLBLM_R_X13Y151_SLICE_X18Y151_CQ;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D1 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_AX = CLBLM_R_X13Y149_SLICE_X19Y149_BO6;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D2 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_B1 = CLBLM_L_X10Y153_SLICE_X12Y153_AQ;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_B2 = CLBLM_R_X13Y149_SLICE_X18Y149_BQ;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_B3 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_B4 = CLBLM_L_X12Y149_SLICE_X17Y149_AQ;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_B5 = CLBLM_R_X7Y146_SLICE_X8Y146_DO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D4 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_D6 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_C1 = CLBLM_L_X10Y145_SLICE_X13Y145_BQ;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_C3 = CLBLM_L_X12Y151_SLICE_X17Y151_AQ;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_C5 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_C6 = 1'b1;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_D1 = CLBLM_L_X12Y148_SLICE_X17Y148_AO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_D2 = CLBLM_R_X5Y155_SLICE_X6Y155_BO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_D3 = CLBLM_R_X13Y149_SLICE_X19Y149_DO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_D4 = CLBLM_L_X12Y149_SLICE_X17Y149_DO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_D5 = CLBLM_L_X12Y156_SLICE_X16Y156_AO6;
  assign CLBLM_R_X13Y149_SLICE_X18Y149_D6 = CLBLM_L_X12Y147_SLICE_X17Y147_AO6;
  assign RIOI3_X105Y191_OLOGIC_X1Y192_T1 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_C1 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_C4 = CLBLM_R_X3Y152_SLICE_X3Y152_AO5;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_CE = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign RIOI3_X105Y191_OLOGIC_X1Y191_D1 = CLBLM_L_X12Y156_SLICE_X16Y156_BQ;
  assign CLBLM_L_X12Y156_SLICE_X17Y156_A1 = 1'b1;
  assign CLBLM_L_X12Y156_SLICE_X17Y156_A2 = CLBLM_R_X11Y158_SLICE_X14Y158_DO5;
  assign CLBLM_L_X12Y156_SLICE_X17Y156_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y156_SLICE_X17Y156_A4 = CLBLM_R_X13Y150_SLICE_X18Y150_AQ;
  assign CLBLM_L_X12Y156_SLICE_X17Y156_A5 = CLBLM_R_X11Y159_SLICE_X15Y159_CO5;
  assign CLBLM_L_X12Y156_SLICE_X17Y156_A6 = CLBLM_L_X12Y156_SLICE_X17Y156_CO6;
  assign CLBLM_L_X12Y156_SLICE_X17Y156_B1 = CLBLM_R_X11Y149_SLICE_X14Y149_DQ;
  assign CLBLM_L_X12Y156_SLICE_X17Y156_B2 = CLBLM_L_X12Y156_SLICE_X17Y156_BQ;
  assign CLBLM_L_X12Y156_SLICE_X17Y156_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y156_SLICE_X17Y156_B4 = CLBLM_R_X11Y158_SLICE_X15Y158_AQ;
  assign CLBLM_L_X12Y156_SLICE_X17Y156_B5 = CLBLM_R_X11Y159_SLICE_X15Y159_DO5;
  assign CLBLM_L_X12Y156_SLICE_X17Y156_B6 = CLBLM_R_X11Y158_SLICE_X15Y158_BO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A1 = CLBLM_L_X10Y146_SLICE_X13Y146_BO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A2 = CLBLM_R_X11Y146_SLICE_X15Y146_AQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A3 = CLBLM_L_X8Y146_SLICE_X11Y146_AQ;
  assign CLBLM_L_X12Y156_SLICE_X17Y156_C4 = CLBLM_L_X12Y156_SLICE_X17Y156_AQ;
  assign CLBLM_L_X12Y156_SLICE_X17Y156_C5 = CLBLM_L_X12Y158_SLICE_X16Y158_CO5;
  assign CLBLM_L_X12Y156_SLICE_X17Y156_C6 = CLBLM_R_X11Y158_SLICE_X15Y158_DO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A4 = CLBLM_R_X11Y146_SLICE_X15Y146_BQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A5 = CLBLM_L_X12Y146_SLICE_X16Y146_AQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_A6 = CLBLM_L_X10Y146_SLICE_X13Y146_CO6;
  assign CLBLM_L_X12Y156_SLICE_X17Y156_C1 = CLBLM_L_X8Y154_SLICE_X10Y154_AQ;
  assign CLBLM_L_X12Y156_SLICE_X17Y156_C2 = CLBLM_R_X11Y158_SLICE_X15Y158_AQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B1 = CLBLM_R_X11Y146_SLICE_X15Y146_CQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B2 = CLBLM_L_X10Y147_SLICE_X13Y147_BQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B3 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_L_X12Y156_SLICE_X17Y156_D1 = CLBLM_R_X11Y152_SLICE_X15Y152_BQ;
  assign CLBLM_L_X12Y156_SLICE_X17Y156_D2 = CLBLM_L_X10Y153_SLICE_X12Y153_AQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B4 = CLBLM_L_X10Y146_SLICE_X12Y146_BQ;
  assign CLBLM_L_X12Y156_SLICE_X17Y156_D4 = CLBLM_L_X12Y159_SLICE_X17Y159_CO6;
  assign CLBLM_L_X12Y156_SLICE_X17Y156_D5 = CLBLM_R_X13Y151_SLICE_X19Y151_AO6;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B5 = CLBLM_L_X8Y146_SLICE_X11Y146_BQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_B6 = CLBLM_L_X8Y146_SLICE_X11Y146_CQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C1 = CLBLM_L_X10Y146_SLICE_X12Y146_AQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C2 = CLBLM_L_X10Y147_SLICE_X12Y147_AQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C3 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C4 = CLBLM_L_X8Y147_SLICE_X11Y147_AQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C5 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_C6 = CLBLM_R_X7Y146_SLICE_X9Y146_AQ;
  assign CLBLM_L_X12Y156_SLICE_X16Y156_A1 = CLBLM_R_X11Y158_SLICE_X15Y158_BO6;
  assign CLBLM_L_X12Y156_SLICE_X16Y156_A2 = CLBLM_R_X11Y159_SLICE_X15Y159_DO5;
  assign CLBLM_L_X12Y156_SLICE_X16Y156_A3 = CLBLM_L_X12Y156_SLICE_X16Y156_BO6;
  assign CLBLM_L_X12Y156_SLICE_X16Y156_A4 = CLBLM_R_X11Y158_SLICE_X15Y158_AQ;
  assign CLBLM_L_X12Y156_SLICE_X16Y156_A5 = CLBLM_L_X10Y158_SLICE_X13Y158_AQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D1 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D2 = CLBLM_R_X11Y152_SLICE_X14Y152_BQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D3 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D4 = CLBLM_L_X10Y149_SLICE_X12Y149_CQ;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D5 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X13Y146_D6 = CLBLM_L_X12Y146_SLICE_X16Y146_AQ;
  assign CLBLM_L_X12Y156_SLICE_X16Y156_B4 = CLBLM_L_X12Y157_SLICE_X16Y157_DO5;
  assign CLBLM_L_X12Y156_SLICE_X16Y156_B5 = CLBLM_R_X13Y150_SLICE_X18Y150_AQ;
  assign CLBLM_L_X12Y156_SLICE_X16Y156_B6 = CLBLM_R_X11Y157_SLICE_X15Y157_CO6;
  assign CLBLM_L_X12Y156_SLICE_X16Y156_AX = CLBLM_R_X7Y155_SLICE_X8Y155_AQ;
  assign CLBLM_L_X12Y156_SLICE_X16Y156_B1 = CLBLM_R_X11Y151_SLICE_X15Y151_CO6;
  assign CLBLM_L_X12Y156_SLICE_X16Y156_B2 = CLBLL_L_X4Y156_SLICE_X4Y156_BO6;
  assign CLBLM_L_X12Y156_SLICE_X16Y156_B3 = CLBLM_L_X12Y156_SLICE_X17Y156_DO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A1 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A2 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A3 = CLBLM_L_X10Y146_SLICE_X12Y146_AQ;
  assign CLBLM_L_X12Y156_SLICE_X16Y156_C4 = CLBLM_R_X11Y158_SLICE_X15Y158_DO6;
  assign CLBLM_L_X12Y156_SLICE_X16Y156_C5 = CLBLM_L_X12Y158_SLICE_X16Y158_BO5;
  assign CLBLM_L_X12Y156_SLICE_X16Y156_C6 = CLBLM_R_X11Y158_SLICE_X14Y158_DO5;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A5 = CLBLM_R_X7Y146_SLICE_X9Y146_DO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_A6 = CLBLM_L_X8Y147_SLICE_X11Y147_AQ;
  assign CLBLM_L_X12Y156_SLICE_X16Y156_C1 = CLBLM_L_X10Y158_SLICE_X13Y158_AQ;
  assign CLBLM_L_X12Y156_SLICE_X16Y156_C2 = CLBLM_R_X11Y159_SLICE_X15Y159_CO5;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B1 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B2 = CLBLM_L_X10Y146_SLICE_X12Y146_BQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B3 = CLBLM_L_X10Y145_SLICE_X12Y145_AQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B5 = CLBLM_R_X7Y146_SLICE_X8Y146_DO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_B6 = CLBLM_R_X11Y152_SLICE_X14Y152_BQ;
  assign CLBLM_L_X12Y156_SLICE_X16Y156_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X12Y156_SLICE_X16Y156_D5 = CLBLM_R_X11Y156_SLICE_X14Y156_AQ;
  assign CLBLM_L_X12Y156_SLICE_X16Y156_D1 = CLBLM_R_X11Y159_SLICE_X15Y159_CO5;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C1 = CLBLM_R_X5Y147_SLICE_X7Y147_AQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C2 = CLBLM_R_X11Y158_SLICE_X14Y158_AQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C4 = CLBLM_L_X10Y145_SLICE_X12Y145_DO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C5 = CLBLM_L_X10Y146_SLICE_X12Y146_DO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_C6 = 1'b1;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y156_SLICE_X16Y156_D6 = CLBLM_R_X11Y157_SLICE_X15Y157_BQ;
  assign CLBLM_L_X12Y156_SLICE_X16Y156_SR = CLBLM_R_X13Y155_SLICE_X18Y155_DO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D1 = CLBLM_L_X10Y146_SLICE_X12Y146_C5Q;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D2 = CLBLM_L_X10Y146_SLICE_X12Y146_CQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D3 = CLBLM_L_X8Y148_SLICE_X11Y148_DO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D4 = CLBLM_L_X10Y145_SLICE_X13Y145_CQ;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D5 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_L_X10Y146_SLICE_X12Y146_D6 = CLBLM_L_X10Y145_SLICE_X13Y145_BQ;
  assign LIOB33_X0Y127_IOB_X0Y127_O = CLBLL_L_X4Y152_SLICE_X4Y152_AQ;
  assign LIOB33_X0Y127_IOB_X0Y128_O = CLBLM_R_X3Y151_SLICE_X2Y151_AQ;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_A1 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_A3 = CLBLM_R_X13Y150_SLICE_X19Y150_AQ;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_A4 = CLBLL_L_X4Y149_SLICE_X4Y149_BQ;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_A5 = CLBLM_R_X7Y148_SLICE_X9Y148_BQ;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_B1 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_B2 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_B3 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_B4 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_B5 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_B6 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_C1 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_C2 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_C3 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_C4 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_C5 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_C6 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_D1 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_D2 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_D3 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_D4 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_D5 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X19Y150_D6 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_C4 = CLBLM_L_X8Y157_SLICE_X11Y157_DO6;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_A1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_A2 = CLBLM_L_X12Y146_SLICE_X16Y146_DQ;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_A3 = CLBLM_R_X13Y150_SLICE_X18Y150_AQ;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_C5 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_A5 = CLBLM_L_X12Y149_SLICE_X16Y149_CQ;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_C6 = CLBLM_R_X7Y155_SLICE_X9Y155_BQ;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_B1 = CLBLM_R_X13Y150_SLICE_X18Y150_DO6;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_B2 = CLBLM_R_X13Y150_SLICE_X18Y150_BQ;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_B3 = CLBLM_R_X11Y154_SLICE_X15Y154_DO6;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_B4 = CLBLM_R_X13Y149_SLICE_X18Y149_DO6;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_B5 = CLBLM_R_X13Y149_SLICE_X19Y149_BO5;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_B6 = CLBLM_R_X13Y149_SLICE_X19Y149_AQ;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_C2 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_C3 = CLBLM_R_X13Y151_SLICE_X18Y151_BQ;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_C4 = CLBLM_L_X12Y150_SLICE_X17Y150_DO6;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_C5 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_C6 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X13Y155_SLICE_X18Y155_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_D1 = CLBLM_R_X13Y149_SLICE_X18Y149_A5Q;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_D2 = CLBLM_R_X13Y149_SLICE_X19Y149_A5Q;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_D3 = CLBLM_R_X13Y149_SLICE_X19Y149_AQ;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_D4 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_D5 = 1'b1;
  assign CLBLM_R_X13Y150_SLICE_X18Y150_D6 = 1'b1;
  assign CLBLM_R_X13Y155_SLICE_X18Y155_C1 = CLBLM_R_X11Y154_SLICE_X14Y154_AQ;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_D2 = CLBLM_L_X8Y157_SLICE_X11Y157_DO6;
  assign CLBLM_R_X13Y155_SLICE_X18Y155_C2 = CLBLM_R_X13Y151_SLICE_X18Y151_DQ;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_D3 = 1'b1;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_D5 = CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  assign CLBLM_R_X13Y155_SLICE_X18Y155_C5 = CLBLM_L_X10Y150_SLICE_X13Y150_BQ;
  assign RIOI3_X105Y127_ILOGIC_X1Y128_D = RIOB33_X105Y127_IOB_X1Y128_I;
  assign RIOI3_X105Y127_ILOGIC_X1Y127_D = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLM_R_X11Y157_SLICE_X15Y157_D6 = CLBLM_L_X12Y157_SLICE_X16Y157_CQ;
  assign CLBLM_R_X13Y155_SLICE_X18Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X12Y157_SLICE_X17Y157_A1 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_L_X12Y157_SLICE_X17Y157_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y157_SLICE_X17Y157_A3 = CLBLM_L_X12Y157_SLICE_X16Y157_A5Q;
  assign CLBLM_L_X12Y157_SLICE_X17Y157_A4 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X12Y157_SLICE_X17Y157_A5 = CLBLL_L_X4Y158_SLICE_X4Y158_AO6;
  assign CLBLM_L_X12Y157_SLICE_X17Y157_A6 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_L_X12Y157_SLICE_X17Y157_AX = CLBLM_R_X13Y157_SLICE_X18Y157_AO6;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y132_D = RIOB33_X105Y131_IOB_X1Y132_I;
  assign CLBLM_L_X12Y157_SLICE_X17Y157_B1 = CLBLM_R_X13Y157_SLICE_X18Y157_BO6;
  assign CLBLM_L_X12Y157_SLICE_X17Y157_B2 = CLBLM_L_X12Y157_SLICE_X17Y157_BQ;
  assign CLBLM_L_X12Y157_SLICE_X17Y157_B3 = CLBLM_R_X11Y159_SLICE_X15Y159_CO5;
  assign CLBLM_L_X12Y157_SLICE_X17Y157_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y157_SLICE_X17Y157_B5 = CLBLM_R_X11Y158_SLICE_X14Y158_DO5;
  assign CLBLM_L_X12Y157_SLICE_X17Y157_B6 = CLBLM_L_X12Y157_SLICE_X16Y157_CQ;
  assign RIOI3_TBYTESRC_X105Y131_ILOGIC_X1Y131_D = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A1 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_L_X12Y157_SLICE_X17Y157_C2 = CLBLM_L_X12Y157_SLICE_X17Y157_CQ;
  assign CLBLM_L_X12Y157_SLICE_X17Y157_C3 = CLBLM_R_X11Y158_SLICE_X15Y158_BO6;
  assign CLBLM_L_X12Y157_SLICE_X17Y157_C4 = CLBLM_R_X11Y159_SLICE_X15Y159_DO5;
  assign CLBLM_L_X12Y157_SLICE_X17Y157_C5 = CLBLM_L_X12Y156_SLICE_X17Y156_BQ;
  assign CLBLM_L_X12Y157_SLICE_X17Y157_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A2 = CLBLM_L_X10Y150_SLICE_X13Y150_CQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A3 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A5 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_A6 = CLBLM_R_X11Y147_SLICE_X15Y147_BO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B1 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B2 = CLBLM_L_X10Y147_SLICE_X13Y147_BQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B3 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_L_X12Y157_SLICE_X17Y157_D1 = 1'b1;
  assign CLBLM_L_X12Y157_SLICE_X17Y157_D2 = CLBLM_L_X12Y157_SLICE_X17Y157_CQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B5 = CLBLM_L_X10Y156_SLICE_X12Y156_AQ;
  assign CLBLM_L_X12Y157_SLICE_X17Y157_D5 = CLBLM_L_X12Y158_SLICE_X16Y158_BO5;
  assign CLBLM_L_X12Y157_SLICE_X17Y157_D6 = CLBLM_L_X12Y159_SLICE_X17Y159_BO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_B6 = CLBLM_R_X11Y146_SLICE_X15Y146_CQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C2 = CLBLM_L_X10Y147_SLICE_X13Y147_CQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C3 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C4 = CLBLM_R_X11Y146_SLICE_X15Y146_CQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C5 = CLBLM_L_X8Y147_SLICE_X11Y147_DO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y157_SLICE_X16Y157_A1 = CLBLM_L_X12Y155_SLICE_X16Y155_BO5;
  assign CLBLM_L_X12Y157_SLICE_X16Y157_A2 = CLBLM_L_X12Y158_SLICE_X16Y158_BO6;
  assign CLBLM_L_X12Y157_SLICE_X16Y157_A6 = CLBLL_L_X4Y148_SLICE_X4Y148_AQ;
  assign CLBLM_L_X12Y157_SLICE_X16Y157_A3 = CLBLM_L_X12Y157_SLICE_X16Y157_AQ;
  assign CLBLM_L_X12Y157_SLICE_X16Y157_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y157_SLICE_X16Y157_AX = CLBLM_L_X12Y153_SLICE_X16Y153_BO6;
  assign CLBLM_L_X12Y157_SLICE_X16Y157_A5 = CLBLM_R_X11Y158_SLICE_X15Y158_BO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D1 = CLBLM_L_X10Y146_SLICE_X13Y146_AO6;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D2 = CLBLM_R_X11Y146_SLICE_X15Y146_BQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D3 = CLBLM_L_X8Y147_SLICE_X10Y147_DO5;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D4 = 1'b1;
  assign CLBLM_L_X12Y157_SLICE_X16Y157_B5 = CLBLM_R_X11Y158_SLICE_X15Y158_BO6;
  assign CLBLM_L_X12Y157_SLICE_X16Y157_B6 = CLBLM_L_X12Y157_SLICE_X17Y157_CQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D5 = CLBLM_R_X11Y146_SLICE_X14Y146_DQ;
  assign CLBLM_L_X10Y147_SLICE_X13Y147_D6 = CLBLM_R_X13Y153_SLICE_X18Y153_CQ;
  assign CLBLM_L_X12Y157_SLICE_X16Y157_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y157_SLICE_X16Y157_B2 = CLBLM_L_X12Y157_SLICE_X16Y157_BQ;
  assign CLBLM_L_X12Y157_SLICE_X16Y157_B3 = CLBLM_R_X11Y155_SLICE_X14Y155_DQ;
  assign CLBLM_L_X12Y157_SLICE_X16Y157_C2 = 1'b1;
  assign CLBLM_L_X12Y157_SLICE_X16Y157_C3 = CLBLM_L_X10Y159_SLICE_X12Y159_CO6;
  assign CLBLM_L_X12Y157_SLICE_X16Y157_C4 = CLBLM_R_X11Y157_SLICE_X15Y157_DO6;
  assign CLBLM_L_X12Y157_SLICE_X16Y157_C5 = 1'b1;
  assign CLBLM_L_X12Y157_SLICE_X16Y157_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A1 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A2 = CLBLM_L_X10Y147_SLICE_X13Y147_DO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A3 = CLBLM_L_X10Y147_SLICE_X12Y147_AQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A5 = CLBLM_L_X8Y154_SLICE_X11Y154_AQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_A6 = CLBLM_R_X7Y146_SLICE_X9Y146_DO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B1 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B2 = CLBLM_R_X11Y147_SLICE_X14Y147_BO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B3 = 1'b1;
  assign CLBLM_L_X12Y157_SLICE_X16Y157_D1 = CLBLM_R_X11Y156_SLICE_X14Y156_AQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B5 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_B6 = CLBLM_R_X5Y155_SLICE_X7Y155_AQ;
  assign CLBLM_L_X12Y157_SLICE_X16Y157_D5 = CLBLM_R_X11Y158_SLICE_X15Y158_BO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C1 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C2 = CLBLM_L_X10Y147_SLICE_X12Y147_CQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C3 = CLBLM_L_X12Y148_SLICE_X16Y148_DO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C4 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C5 = CLBLM_R_X7Y148_SLICE_X8Y148_A5Q;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y157_SLICE_X16Y157_D6 = 1'b1;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D1 = CLBLM_L_X8Y147_SLICE_X10Y147_AQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D2 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D3 = CLBLM_L_X10Y147_SLICE_X12Y147_DQ;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D5 = CLBLM_L_X10Y148_SLICE_X12Y148_DO6;
  assign CLBLM_L_X10Y147_SLICE_X12Y147_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_C4 = CLBLM_R_X11Y159_SLICE_X15Y159_DO5;
  assign CLBLM_R_X7Y159_SLICE_X9Y159_D5 = CLBLM_R_X11Y159_SLICE_X14Y159_CQ;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X7Y159_SLICE_X9Y159_D6 = CLBLL_L_X4Y157_SLICE_X4Y157_CO5;
  assign CLBLM_R_X11Y157_SLICE_X14Y157_C6 = CLBLM_R_X11Y158_SLICE_X15Y158_BO6;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_A1 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_A2 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_A3 = CLBLM_R_X13Y150_SLICE_X19Y150_AQ;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_A5 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_A6 = CLBLL_L_X4Y149_SLICE_X4Y149_BQ;
  assign RIOI3_X105Y129_ILOGIC_X1Y130_D = RIOB33_X105Y129_IOB_X1Y130_I;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_B1 = CLBLM_R_X11Y151_SLICE_X14Y151_AQ;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_B2 = CLBLM_R_X13Y153_SLICE_X18Y153_BQ;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_B3 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_B4 = CLBLM_L_X12Y153_SLICE_X16Y153_AQ;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_B5 = CLBLM_R_X13Y153_SLICE_X19Y153_AQ;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_B6 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_C1 = CLBLM_R_X13Y151_SLICE_X18Y151_AQ;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_C2 = CLBLM_R_X13Y152_SLICE_X19Y152_AQ;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_C3 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_C4 = CLBLM_L_X10Y151_SLICE_X12Y151_BQ;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_C5 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_C6 = 1'b1;
  assign RIOI3_X105Y129_ILOGIC_X1Y129_D = RIOB33_X105Y129_IOB_X1Y129_I;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_D1 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_D2 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_D3 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_D4 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_D5 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X19Y151_D6 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_A1 = CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_A2 = CLBLM_R_X11Y156_SLICE_X14Y156_BQ;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_A3 = CLBLM_R_X13Y151_SLICE_X18Y151_AQ;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_A4 = CLBLM_L_X12Y153_SLICE_X16Y153_AQ;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_B1 = CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_B2 = CLBLM_R_X13Y151_SLICE_X18Y151_BQ;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_B4 = CLBLM_L_X10Y151_SLICE_X12Y151_BQ;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_B5 = CLBLM_R_X13Y153_SLICE_X18Y153_AQ;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_C2 = CLBLM_L_X12Y149_SLICE_X16Y149_CQ;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_C3 = CLBLM_R_X13Y155_SLICE_X18Y155_BQ;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_C4 = CLBLM_R_X11Y150_SLICE_X15Y150_AO5;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_C5 = 1'b1;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_C6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_D2 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_D3 = CLBLM_R_X13Y151_SLICE_X18Y151_DQ;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_D4 = CLBLM_R_X11Y151_SLICE_X15Y151_A5Q;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_D5 = CLBLM_L_X10Y152_SLICE_X13Y152_DO6;
  assign CLBLM_R_X13Y151_SLICE_X18Y151_D6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X7Y159_SLICE_X8Y159_B5 = CLBLM_R_X7Y148_SLICE_X8Y148_AQ;
  assign CLBLM_R_X7Y159_SLICE_X8Y159_B6 = 1'b1;
  assign CLBLM_R_X13Y156_SLICE_X18Y156_B2 = CLBLM_L_X12Y157_SLICE_X16Y157_BQ;
  assign CLBLM_R_X7Y159_SLICE_X8Y159_C4 = 1'b1;
  assign CLBLM_R_X7Y159_SLICE_X8Y159_C5 = 1'b1;
  assign CLBLM_L_X12Y158_SLICE_X17Y158_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y158_SLICE_X17Y158_A2 = CLBLM_L_X12Y158_SLICE_X16Y158_DO6;
  assign CLBLM_L_X12Y158_SLICE_X17Y158_A3 = CLBLM_R_X11Y158_SLICE_X15Y158_BO6;
  assign CLBLM_L_X12Y158_SLICE_X17Y158_A4 = CLBLM_L_X12Y158_SLICE_X17Y158_AQ;
  assign CLBLM_L_X12Y158_SLICE_X17Y158_A5 = CLBLM_R_X13Y155_SLICE_X18Y155_AQ;
  assign CLBLM_L_X12Y158_SLICE_X17Y158_A6 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_R_X7Y159_SLICE_X8Y159_C6 = 1'b1;
  assign CLBLM_L_X12Y158_SLICE_X17Y158_B1 = 1'b1;
  assign CLBLM_L_X12Y158_SLICE_X17Y158_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y158_SLICE_X17Y158_B3 = CLBLM_R_X11Y158_SLICE_X15Y158_BO6;
  assign CLBLM_L_X12Y158_SLICE_X17Y158_B4 = CLBLM_R_X5Y148_SLICE_X6Y148_CO6;
  assign CLBLM_L_X12Y158_SLICE_X17Y158_B5 = CLBLM_R_X13Y158_SLICE_X18Y158_AQ;
  assign CLBLM_L_X12Y158_SLICE_X17Y158_B6 = CLBLM_L_X12Y158_SLICE_X17Y158_CO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A1 = CLBLM_L_X10Y148_SLICE_X13Y148_AQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A3 = CLBLM_L_X10Y148_SLICE_X12Y148_CO5;
  assign CLBLM_L_X12Y158_SLICE_X17Y158_C4 = CLBLM_L_X12Y158_SLICE_X17Y158_BQ;
  assign CLBLM_L_X12Y158_SLICE_X17Y158_C5 = CLBLM_L_X12Y158_SLICE_X17Y158_DO6;
  assign CLBLM_L_X12Y158_SLICE_X17Y158_C6 = CLBLM_R_X11Y159_SLICE_X14Y159_AQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A4 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A5 = CLBLM_L_X12Y149_SLICE_X17Y149_AQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_A6 = CLBLM_L_X8Y149_SLICE_X11Y149_DO6;
  assign CLBLM_L_X12Y158_SLICE_X17Y158_C1 = CLBLM_L_X12Y152_SLICE_X17Y152_A5Q;
  assign CLBLM_L_X12Y158_SLICE_X17Y158_C2 = CLBLM_L_X12Y159_SLICE_X17Y159_CO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B2 = CLBLM_L_X10Y148_SLICE_X13Y148_BQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B3 = CLBLM_L_X10Y148_SLICE_X12Y148_CO5;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B4 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_L_X12Y158_SLICE_X17Y158_D2 = CLBLM_L_X12Y158_SLICE_X17Y158_AQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B5 = CLBLM_R_X13Y153_SLICE_X18Y153_C5Q;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_B6 = CLBLM_L_X10Y155_SLICE_X12Y155_BQ;
  assign CLBLM_L_X12Y158_SLICE_X17Y158_D5 = CLBLM_L_X12Y157_SLICE_X16Y157_AQ;
  assign CLBLM_L_X12Y158_SLICE_X17Y158_D6 = CLBLM_R_X11Y159_SLICE_X14Y159_BQ;
  assign CLBLM_L_X12Y158_SLICE_X17Y158_D1 = CLBLM_L_X12Y158_SLICE_X16Y158_AQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C1 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C2 = CLBLM_L_X12Y146_SLICE_X16Y146_CQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C3 = CLBLM_L_X10Y150_SLICE_X13Y150_DO6;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C5 = CLBLM_L_X10Y148_SLICE_X13Y148_CQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_C6 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_A2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_A3 = CLBLM_L_X12Y158_SLICE_X16Y158_AQ;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_A4 = CLBLM_L_X12Y159_SLICE_X17Y159_AO6;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_A5 = CLBLM_L_X12Y157_SLICE_X17Y157_AQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D1 = CLBLM_L_X10Y148_SLICE_X13Y148_BQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D3 = CLBLM_R_X11Y152_SLICE_X15Y152_DQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D4 = CLBLM_L_X10Y155_SLICE_X12Y155_BQ;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D5 = CLBLM_L_X10Y148_SLICE_X13Y148_AQ;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_B5 = CLBLM_L_X12Y158_SLICE_X17Y158_AQ;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_B6 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X13Y148_D6 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_AX = CLBLM_L_X12Y159_SLICE_X16Y159_AO6;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_B1 = CLBLM_L_X12Y157_SLICE_X16Y157_AQ;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_B2 = CLBLM_R_X11Y159_SLICE_X15Y159_AQ;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_B3 = CLBLM_L_X12Y159_SLICE_X16Y159_BO5;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_B4 = CLBLM_L_X12Y155_SLICE_X16Y155_BO5;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A1 = CLBLM_L_X8Y148_SLICE_X11Y148_B5Q;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_C4 = CLBLM_L_X12Y158_SLICE_X17Y158_AQ;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_C5 = CLBLM_R_X11Y159_SLICE_X14Y159_BQ;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_C6 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A2 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A3 = CLBLM_L_X10Y148_SLICE_X12Y148_AQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_A6 = 1'b1;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B3 = CLBLM_L_X10Y151_SLICE_X12Y151_AQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B4 = CLBLM_L_X10Y147_SLICE_X12Y147_DQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B5 = CLBLM_R_X5Y152_SLICE_X6Y152_BQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_B6 = 1'b1;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_D1 = CLBLM_L_X12Y158_SLICE_X17Y158_AQ;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_D2 = CLBLM_L_X12Y158_SLICE_X16Y158_AQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C1 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C3 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C4 = CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_C6 = 1'b1;
  assign CLBLM_L_X12Y158_SLICE_X16Y158_D5 = CLBLM_L_X12Y159_SLICE_X16Y159_BO5;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D1 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D2 = CLBLM_R_X3Y152_SLICE_X3Y152_BO5;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D4 = CLBLM_L_X10Y148_SLICE_X12Y148_CO6;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D5 = CLBLM_L_X8Y150_SLICE_X11Y150_BQ;
  assign CLBLM_L_X10Y148_SLICE_X12Y148_D6 = CLBLM_R_X5Y152_SLICE_X6Y152_BQ;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A1 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A3 = CLBLM_R_X13Y154_SLICE_X18Y154_AQ;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A5 = CLBLM_R_X13Y157_SLICE_X18Y157_AQ;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_A6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_B6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_C6 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_A1 = CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_A3 = CLBLM_R_X13Y152_SLICE_X19Y152_AQ;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_A5 = CLBLM_R_X11Y157_SLICE_X15Y157_BQ;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_A6 = CLBLM_R_X11Y152_SLICE_X15Y152_CQ;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X163Y177_D2 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_B1 = CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_B4 = CLBLM_L_X12Y151_SLICE_X16Y151_BQ;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_B5 = CLBLM_R_X13Y152_SLICE_X18Y152_AQ;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_B6 = CLBLM_R_X13Y152_SLICE_X19Y152_BQ;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A3 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_C1 = CLBLM_R_X13Y152_SLICE_X18Y152_AQ;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_C2 = CLBLM_R_X13Y151_SLICE_X19Y151_CO6;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_C3 = CLBLM_L_X12Y152_SLICE_X17Y152_CO6;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_C4 = CLBLM_R_X13Y152_SLICE_X19Y152_BQ;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_C5 = CLBLM_L_X12Y155_SLICE_X16Y155_AO5;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_C6 = CLBLM_R_X13Y151_SLICE_X19Y151_BO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_A5 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D4 = CLBLM_L_X12Y154_SLICE_X16Y154_A5Q;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_B2 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D5 = CLBLM_L_X10Y146_SLICE_X12Y146_AQ;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_D1 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_D2 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_D3 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_D4 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D6 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_D5 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X19Y152_D6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C1 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C2 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C3 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_C4 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_A1 = CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_A2 = CLBLM_R_X11Y152_SLICE_X14Y152_AQ;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_A3 = CLBLM_R_X13Y152_SLICE_X18Y152_AQ;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_A4 = CLBLM_R_X11Y152_SLICE_X15Y152_BQ;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D1 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_AX = CLBLM_R_X13Y152_SLICE_X18Y152_BO6;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D2 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_B2 = CLBLM_R_X13Y152_SLICE_X18Y152_A5Q;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_B3 = CLBLM_R_X5Y155_SLICE_X6Y155_DO6;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_B5 = CLBLM_L_X10Y151_SLICE_X13Y151_AQ;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_B6 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D4 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D5 = 1'b1;
  assign CLBLM_R_X103Y177_SLICE_X162Y177_D6 = 1'b1;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_C2 = CLBLM_R_X13Y152_SLICE_X18Y152_CQ;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_C3 = CLBLM_L_X12Y150_SLICE_X17Y150_BQ;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_C4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_C5 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_C6 = CLBLM_R_X13Y152_SLICE_X19Y152_BQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A1 = CLBLM_L_X10Y146_SLICE_X12Y146_C5Q;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A2 = CLBLM_L_X10Y146_SLICE_X12Y146_CQ;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_D1 = CLBLM_R_X13Y154_SLICE_X19Y154_AQ;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_D2 = CLBLM_R_X13Y152_SLICE_X19Y152_CO6;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_D3 = CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A3 = CLBLM_L_X12Y149_SLICE_X17Y149_A5Q;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_D4 = CLBLM_R_X5Y155_SLICE_X6Y155_BO6;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_D5 = CLBLM_L_X12Y155_SLICE_X16Y155_AO5;
  assign CLBLM_R_X13Y152_SLICE_X18Y152_D6 = CLBLM_R_X7Y148_SLICE_X9Y148_BQ;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_A1 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_A2 = CLBLM_L_X12Y158_SLICE_X16Y158_BO5;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_A3 = CLBLM_R_X13Y158_SLICE_X18Y158_AQ;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_A4 = CLBLM_R_X13Y159_SLICE_X18Y159_AO6;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_A5 = CLBLM_R_X13Y159_SLICE_X18Y159_BO6;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_A6 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_B1 = CLBLM_L_X12Y158_SLICE_X16Y158_AQ;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_B2 = CLBLM_L_X12Y157_SLICE_X17Y157_BQ;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_B3 = CLBLM_L_X12Y156_SLICE_X17Y156_AQ;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_B4 = CLBLM_L_X12Y158_SLICE_X17Y158_AQ;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_B5 = CLBLM_L_X8Y154_SLICE_X10Y154_AQ;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_B6 = CLBLM_R_X11Y159_SLICE_X15Y159_AQ;
  assign LIOB33_X0Y133_IOB_X0Y133_O = CLBLM_R_X5Y146_SLICE_X6Y146_A5Q;
  assign LIOB33_X0Y133_IOB_X0Y134_O = CLBLM_R_X7Y145_SLICE_X8Y145_AQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A1 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A3 = CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_C4 = CLBLM_R_X11Y159_SLICE_X15Y159_AQ;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_C5 = CLBLM_L_X12Y158_SLICE_X16Y158_AQ;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_C6 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A4 = CLBLM_R_X11Y148_SLICE_X14Y148_BQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_A6 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_C1 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_C2 = CLBLM_R_X11Y159_SLICE_X14Y159_AQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_AX = CLBLM_L_X10Y149_SLICE_X13Y149_BO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B1 = CLBLM_R_X11Y152_SLICE_X14Y152_CQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B2 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B3 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B5 = CLBLM_R_X11Y149_SLICE_X15Y149_BO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_B6 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_D5 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_D6 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_D1 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_BX = CLBLM_R_X11Y150_SLICE_X15Y150_AO6;
  assign CLBLM_L_X12Y159_SLICE_X17Y159_D2 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C1 = CLBLL_L_X4Y153_SLICE_X4Y153_BO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C2 = CLBLM_R_X13Y155_SLICE_X19Y155_AO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C4 = CLBLM_L_X10Y147_SLICE_X13Y147_CQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C5 = CLBLM_L_X10Y149_SLICE_X13Y149_DO6;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_C6 = CLBLM_L_X12Y151_SLICE_X16Y151_BQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_A1 = CLBLM_L_X8Y153_SLICE_X11Y153_CQ;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_A2 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_A3 = CLBLM_L_X12Y159_SLICE_X16Y159_AQ;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D1 = CLBLM_R_X11Y146_SLICE_X14Y146_BQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D2 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D3 = CLBLM_R_X7Y153_SLICE_X9Y153_AQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D4 = CLBLM_L_X10Y145_SLICE_X13Y145_AQ;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D5 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_B5 = CLBLM_R_X11Y157_SLICE_X15Y157_AQ;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_B6 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X13Y149_D6 = CLBLM_L_X8Y149_SLICE_X11Y149_BQ;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_AX = CLBLM_L_X12Y158_SLICE_X17Y158_AQ;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_BX = CLBLM_L_X10Y150_SLICE_X12Y150_CQ;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_B2 = CLBLM_R_X11Y159_SLICE_X14Y159_BQ;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_B3 = CLBLM_L_X12Y159_SLICE_X17Y159_AO6;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_B4 = CLBLM_R_X11Y159_SLICE_X14Y159_AQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A2 = CLBLL_L_X4Y150_SLICE_X5Y150_C5Q;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_C5 = CLBLM_L_X12Y159_SLICE_X16Y159_BQ;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_C6 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A3 = CLBLM_L_X12Y157_SLICE_X17Y157_A5Q;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A5 = CLBLL_L_X4Y151_SLICE_X5Y151_CQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_A6 = CLBLM_L_X8Y148_SLICE_X11Y148_BQ;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_C2 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B1 = CLBLM_L_X10Y151_SLICE_X13Y151_B5Q;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B2 = CLBLM_L_X10Y149_SLICE_X12Y149_BQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B3 = CLBLM_L_X10Y149_SLICE_X12Y149_AQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_B6 = CLBLM_L_X8Y153_SLICE_X10Y153_A5Q;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_D5 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_D1 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C2 = CLBLM_L_X10Y149_SLICE_X13Y149_BQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C3 = CLBLM_L_X10Y152_SLICE_X12Y152_BQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C4 = CLBLM_L_X10Y151_SLICE_X12Y151_BQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_C6 = 1'b1;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_D6 = 1'b1;
  assign CLBLM_L_X12Y159_SLICE_X16Y159_SR = CLBLM_R_X13Y155_SLICE_X18Y155_DO6;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D2 = CLBLL_L_X4Y150_SLICE_X5Y150_DQ;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D3 = CLBLM_L_X10Y151_SLICE_X13Y151_B5Q;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D4 = CLBLM_L_X8Y153_SLICE_X10Y153_A5Q;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y149_SLICE_X12Y149_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y144_D = RIOB33_X105Y143_IOB_X1Y144_I;
  assign RIOI3_TBYTESRC_X105Y143_ILOGIC_X1Y143_D = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X13Y153_SLICE_X19Y153_A1 = CLBLM_R_X13Y153_SLICE_X19Y153_DO6;
  assign CLBLM_R_X13Y153_SLICE_X19Y153_A2 = CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  assign CLBLM_R_X13Y153_SLICE_X19Y153_A3 = CLBLM_R_X13Y153_SLICE_X19Y153_AQ;
  assign CLBLM_R_X13Y153_SLICE_X19Y153_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y153_SLICE_X19Y153_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y153_SLICE_X19Y153_A6 = CLBLM_R_X13Y153_SLICE_X19Y153_BQ;
  assign CLBLM_R_X13Y153_SLICE_X19Y153_B1 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X13Y153_SLICE_X19Y153_B2 = CLBLM_R_X13Y153_SLICE_X19Y153_BQ;
  assign CLBLM_R_X13Y153_SLICE_X19Y153_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y153_SLICE_X19Y153_B4 = CLBLM_L_X12Y149_SLICE_X16Y149_B5Q;
  assign CLBLM_R_X13Y153_SLICE_X19Y153_B5 = 1'b1;
  assign CLBLM_R_X13Y153_SLICE_X19Y153_B6 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_R_X13Y153_SLICE_X19Y153_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y153_SLICE_X19Y153_C2 = CLBLM_R_X13Y153_SLICE_X19Y153_CQ;
  assign CLBLM_R_X13Y153_SLICE_X19Y153_C3 = CLBLM_L_X12Y153_SLICE_X17Y153_CQ;
  assign CLBLM_R_X13Y153_SLICE_X19Y153_C4 = 1'b1;
  assign CLBLM_R_X13Y153_SLICE_X19Y153_C5 = CLBLM_L_X8Y155_SLICE_X11Y155_CQ;
  assign CLBLM_R_X13Y153_SLICE_X19Y153_C6 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_R_X13Y153_SLICE_X19Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X13Y153_SLICE_X19Y153_D1 = CLBLM_R_X13Y155_SLICE_X19Y155_AO6;
  assign CLBLM_R_X13Y153_SLICE_X19Y153_D2 = CLBLM_R_X13Y154_SLICE_X19Y154_AQ;
  assign CLBLM_R_X13Y153_SLICE_X19Y153_D3 = CLBLM_R_X7Y148_SLICE_X9Y148_BQ;
  assign CLBLM_R_X13Y153_SLICE_X19Y153_D4 = CLBLM_R_X13Y152_SLICE_X19Y152_CO6;
  assign CLBLM_R_X13Y153_SLICE_X19Y153_D5 = CLBLM_L_X12Y155_SLICE_X16Y155_AO5;
  assign CLBLM_R_X13Y153_SLICE_X19Y153_D6 = CLBLM_R_X5Y155_SLICE_X6Y155_DO6;
  assign CLBLM_R_X13Y153_SLICE_X18Y153_A1 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X13Y153_SLICE_X18Y153_A2 = CLBLM_R_X13Y152_SLICE_X18Y152_CQ;
  assign CLBLM_R_X13Y153_SLICE_X18Y153_A3 = CLBLM_R_X13Y153_SLICE_X18Y153_AQ;
  assign CLBLM_R_X13Y153_SLICE_X18Y153_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y153_SLICE_X18Y153_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y153_SLICE_X18Y153_A6 = CLBLM_R_X13Y154_SLICE_X18Y154_AQ;
  assign CLBLM_R_X13Y153_SLICE_X18Y153_B1 = CLBLM_R_X13Y151_SLICE_X18Y151_BQ;
  assign CLBLM_R_X13Y153_SLICE_X18Y153_B2 = CLBLM_R_X13Y153_SLICE_X18Y153_BQ;
  assign CLBLM_R_X13Y153_SLICE_X18Y153_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y153_SLICE_X18Y153_B4 = CLBLM_L_X12Y156_SLICE_X17Y156_BQ;
  assign CLBLM_R_X13Y153_SLICE_X18Y153_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y153_SLICE_X18Y153_B6 = CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  assign CLBLM_R_X13Y153_SLICE_X18Y153_C1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y153_SLICE_X18Y153_C2 = CLBLM_L_X10Y145_SLICE_X13Y145_CQ;
  assign CLBLM_R_X13Y153_SLICE_X18Y153_C3 = CLBLM_L_X10Y154_SLICE_X13Y154_AQ;
  assign CLBLM_R_X13Y153_SLICE_X18Y153_C4 = CLBLM_L_X12Y158_SLICE_X17Y158_BQ;
  assign CLBLM_R_X13Y153_SLICE_X18Y153_C5 = CLBLM_R_X13Y148_SLICE_X18Y148_AQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A1 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A2 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A3 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A4 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A5 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_A6 = 1'b1;
  assign CLBLM_R_X13Y153_SLICE_X18Y153_C6 = 1'b1;
  assign CLBLM_R_X13Y153_SLICE_X18Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B1 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B2 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B3 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B4 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B5 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_B6 = 1'b1;
  assign CLBLM_R_X13Y153_SLICE_X18Y153_D1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y153_SLICE_X18Y153_D2 = CLBLM_L_X10Y152_SLICE_X13Y152_DO6;
  assign CLBLM_R_X13Y153_SLICE_X18Y153_D3 = CLBLM_R_X13Y153_SLICE_X18Y153_DQ;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C1 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C2 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C3 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C4 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C5 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_C6 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D1 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D2 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D3 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D4 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D5 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X4Y146_D6 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A1 = CLBLM_R_X5Y149_SLICE_X7Y149_CQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A2 = CLBLM_R_X5Y144_SLICE_X6Y144_CO6;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A3 = CLBLM_R_X5Y146_SLICE_X6Y146_BQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A4 = CLBLM_R_X5Y144_SLICE_X6Y144_AQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_A6 = 1'b1;
  assign LIOB33_X0Y135_IOB_X0Y136_O = CLBLM_R_X7Y144_SLICE_X8Y144_AQ;
  assign LIOB33_X0Y135_IOB_X0Y135_O = CLBLM_R_X5Y146_SLICE_X6Y146_AQ;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B1 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B2 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B3 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B4 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B5 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_B6 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C1 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C2 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C3 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C4 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C5 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_C6 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D1 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D2 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D3 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D4 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D5 = 1'b1;
  assign CLBLL_L_X4Y146_SLICE_X5Y146_D6 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A2 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A4 = CLBLM_L_X12Y151_SLICE_X16Y151_BQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A5 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_A6 = CLBLM_R_X7Y147_SLICE_X9Y147_CQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B1 = CLBLM_R_X7Y149_SLICE_X9Y149_CQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B2 = RIOB33_X105Y119_IOB_X1Y119_I;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B3 = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B5 = CLBLM_L_X10Y150_SLICE_X13Y150_BQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_B6 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C1 = CLBLM_L_X10Y147_SLICE_X13Y147_AQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C2 = CLBLM_L_X10Y150_SLICE_X12Y150_BQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C3 = CLBLM_R_X7Y152_SLICE_X9Y152_BQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C5 = CLBLM_L_X10Y153_SLICE_X12Y153_DO6;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_C6 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D1 = CLBLM_R_X7Y149_SLICE_X8Y149_DO5;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D2 = CLBLM_R_X7Y154_SLICE_X8Y154_AO5;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D3 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D4 = CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y150_SLICE_X13Y150_D6 = CLBLM_R_X7Y150_SLICE_X9Y150_AO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A1 = CLBLM_L_X10Y149_SLICE_X12Y149_AQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A2 = CLBLM_R_X11Y156_SLICE_X15Y156_BQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A4 = CLBLM_L_X10Y150_SLICE_X12Y150_AQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_A6 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B1 = CLBLM_L_X8Y152_SLICE_X10Y152_BQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B2 = CLBLM_L_X8Y150_SLICE_X10Y150_BQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B3 = CLBLM_L_X10Y150_SLICE_X12Y150_AQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B4 = CLBLM_R_X7Y151_SLICE_X8Y151_CQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B5 = CLBLM_L_X8Y147_SLICE_X10Y147_CQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_B6 = 1'b1;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_BX = CLBLM_L_X10Y153_SLICE_X13Y153_BO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C1 = CLBLM_L_X8Y147_SLICE_X10Y147_CQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C2 = CLBLM_L_X8Y150_SLICE_X10Y150_BQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C3 = CLBLM_L_X8Y152_SLICE_X10Y152_BQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C4 = CLBLM_R_X7Y151_SLICE_X8Y151_CQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C5 = CLBLM_R_X13Y152_SLICE_X18Y152_A5Q;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_C6 = CLBLM_R_X5Y147_SLICE_X7Y147_BQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_CX = CLBLM_L_X10Y149_SLICE_X12Y149_DO6;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D1 = CLBLM_L_X10Y148_SLICE_X12Y148_AQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D2 = CLBLM_L_X8Y151_SLICE_X10Y151_BQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D3 = CLBLM_L_X10Y151_SLICE_X12Y151_DQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D4 = CLBLM_R_X11Y148_SLICE_X14Y148_BQ;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D5 = CLBLM_R_X13Y152_SLICE_X18Y152_A5Q;
  assign CLBLM_L_X10Y150_SLICE_X12Y150_D6 = CLBLM_L_X10Y150_SLICE_X12Y150_AQ;
  assign CLBLM_R_X13Y154_SLICE_X19Y154_A1 = CLBLM_R_X13Y154_SLICE_X19Y154_AQ;
  assign CLBLM_R_X13Y154_SLICE_X19Y154_A2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y154_SLICE_X19Y154_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y154_SLICE_X19Y154_A4 = CLBLM_R_X13Y154_SLICE_X18Y154_BQ;
  assign CLBLM_R_X13Y154_SLICE_X19Y154_A5 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X13Y154_SLICE_X19Y154_A6 = CLBLM_L_X10Y155_SLICE_X13Y155_A5Q;
  assign CLBLM_R_X13Y154_SLICE_X19Y154_B1 = 1'b1;
  assign CLBLM_R_X13Y154_SLICE_X19Y154_B2 = 1'b1;
  assign CLBLM_R_X13Y154_SLICE_X19Y154_B3 = 1'b1;
  assign CLBLM_R_X13Y154_SLICE_X19Y154_B4 = 1'b1;
  assign CLBLM_R_X13Y154_SLICE_X19Y154_B5 = 1'b1;
  assign CLBLM_R_X13Y154_SLICE_X19Y154_B6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A2 = CLBLM_L_X12Y157_SLICE_X17Y157_BQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A3 = CLBLM_R_X5Y146_SLICE_X6Y146_AQ;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A4 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A5 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_A6 = 1'b1;
  assign CLBLM_R_X13Y154_SLICE_X19Y154_C1 = 1'b1;
  assign CLBLM_R_X13Y154_SLICE_X19Y154_C2 = 1'b1;
  assign CLBLM_R_X13Y154_SLICE_X19Y154_C3 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B1 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B2 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B3 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B4 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B5 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_B6 = 1'b1;
  assign CLBLM_R_X13Y154_SLICE_X19Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X13Y154_SLICE_X19Y154_D1 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C1 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C2 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C3 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C4 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C5 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_C6 = 1'b1;
  assign CLBLM_R_X13Y154_SLICE_X19Y154_D3 = 1'b1;
  assign CLBLM_R_X13Y154_SLICE_X19Y154_D4 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y154_SLICE_X18Y154_A1 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X13Y154_SLICE_X18Y154_A2 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_R_X13Y154_SLICE_X18Y154_A3 = CLBLM_R_X13Y154_SLICE_X18Y154_AQ;
  assign CLBLM_R_X13Y154_SLICE_X18Y154_A4 = CLBLM_L_X8Y154_SLICE_X11Y154_CQ;
  assign CLBLM_R_X13Y154_SLICE_X18Y154_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D1 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D2 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D3 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D4 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D5 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X15Y144_D6 = 1'b1;
  assign CLBLM_R_X13Y154_SLICE_X18Y154_A6 = 1'b1;
  assign CLBLM_R_X13Y154_SLICE_X18Y154_B1 = CLBLM_R_X13Y148_SLICE_X18Y148_AQ;
  assign CLBLM_R_X13Y154_SLICE_X18Y154_B2 = CLBLM_R_X13Y154_SLICE_X18Y154_BQ;
  assign CLBLM_R_X13Y154_SLICE_X18Y154_B3 = CLBLM_L_X12Y153_SLICE_X17Y153_AQ;
  assign CLBLM_R_X13Y154_SLICE_X18Y154_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A1 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A2 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A1 = CLBLL_L_X4Y154_SLICE_X5Y154_CO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A2 = CLBLL_L_X4Y151_SLICE_X4Y151_C5Q;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A3 = CLBLL_L_X4Y154_SLICE_X5Y154_BO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A5 = CLBLM_R_X3Y151_SLICE_X2Y151_AQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_A6 = CLBLM_R_X5Y149_SLICE_X6Y149_B5Q;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A3 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A4 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_A5 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B2 = CLBLL_L_X4Y151_SLICE_X4Y151_C5Q;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B3 = CLBLM_L_X8Y147_SLICE_X11Y147_CO6;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B4 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B5 = CLBLM_R_X3Y151_SLICE_X2Y151_AQ;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_B6 = CLBLM_R_X5Y149_SLICE_X6Y149_B5Q;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B1 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_B2 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C1 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C2 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C3 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C4 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C5 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_C6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C1 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C2 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C3 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C4 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C5 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_C6 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D1 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D2 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D3 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D4 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D5 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X4Y147_D6 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D1 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D2 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D3 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D4 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D5 = 1'b1;
  assign CLBLM_R_X11Y144_SLICE_X14Y144_D6 = 1'b1;
  assign LIOI3_SING_X0Y50_ILOGIC_X0Y50_D = LIOB33_SING_X0Y50_IOB_X0Y50_I;
  assign LIOB33_X0Y137_IOB_X0Y138_O = CLBLM_R_X5Y146_SLICE_X6Y146_BQ;
  assign LIOB33_X0Y137_IOB_X0Y137_O = CLBLM_R_X5Y144_SLICE_X6Y144_BQ;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_D1 = LIOB33_X0Y65_IOB_X0Y66_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y152_T1 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_D1 = CLBLM_L_X12Y159_SLICE_X16Y159_AQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A2 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A3 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A4 = CLBLM_R_X5Y147_SLICE_X6Y147_AQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A5 = CLBLL_L_X4Y146_SLICE_X5Y146_AO5;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_A6 = CLBLM_L_X10Y148_SLICE_X13Y148_BQ;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_D1 = LIOB33_X0Y65_IOB_X0Y65_I;
  assign RIOI3_X105Y195_OLOGIC_X1Y196_T1 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B2 = CLBLL_L_X4Y147_SLICE_X5Y147_BQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B3 = CLBLM_R_X7Y147_SLICE_X9Y147_AQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B4 = CLBLM_R_X5Y149_SLICE_X6Y149_B5Q;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B5 = CLBLL_L_X4Y146_SLICE_X5Y146_AO5;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign LIOI3_X0Y151_OLOGIC_X0Y151_T1 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C1 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C2 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C3 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C4 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C5 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_C6 = 1'b1;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_D1 = CLBLM_R_X13Y157_SLICE_X18Y157_AQ;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign RIOI3_X105Y195_OLOGIC_X1Y195_T1 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D1 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D2 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D3 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D4 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D5 = 1'b1;
  assign CLBLL_L_X4Y147_SLICE_X5Y147_D6 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A1 = CLBLM_L_X10Y151_SLICE_X13Y151_DO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A2 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A3 = CLBLM_L_X10Y151_SLICE_X13Y151_AQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A5 = CLBLM_R_X11Y149_SLICE_X14Y149_BQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y156_SLICE_X19Y156_C4 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B1 = CLBLM_L_X8Y153_SLICE_X10Y153_A5Q;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B3 = CLBLM_R_X7Y148_SLICE_X8Y148_AQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B5 = CLBLM_R_X11Y151_SLICE_X14Y151_BQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_B6 = 1'b1;
  assign CLBLM_R_X13Y156_SLICE_X19Y156_C5 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_D1 = CLBLL_L_X36Y150_SLICE_X54Y150_AO6;
  assign CLBLM_R_X13Y156_SLICE_X19Y156_C6 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C3 = CLBLM_L_X10Y154_SLICE_X13Y154_CQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C4 = CLBLM_L_X10Y158_SLICE_X13Y158_BQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C5 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y158_SLICE_X18Y158_A2 = CLBLM_R_X11Y158_SLICE_X14Y158_DO5;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y158_T1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D1 = CLBLM_L_X10Y154_SLICE_X13Y154_C5Q;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D2 = CLBLM_L_X8Y152_SLICE_X10Y152_BQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D3 = CLBLM_L_X8Y152_SLICE_X11Y152_BO6;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D4 = CLBLM_L_X10Y158_SLICE_X13Y158_BQ;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D5 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y151_SLICE_X13Y151_D6 = CLBLM_L_X8Y150_SLICE_X10Y150_BQ;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_D1 = RIOB33_X105Y125_IOB_X1Y126_I;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A1 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A2 = CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A3 = CLBLM_L_X10Y151_SLICE_X12Y151_AQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_A6 = CLBLM_L_X8Y153_SLICE_X11Y153_BQ;
  assign CLBLM_R_X13Y158_SLICE_X18Y158_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign RIOI3_TBYTESRC_X105Y157_OLOGIC_X1Y157_T1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B2 = CLBLM_R_X11Y151_SLICE_X14Y151_AQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B3 = CLBLM_L_X8Y147_SLICE_X10Y147_CQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B4 = CLBLM_R_X11Y149_SLICE_X15Y149_DO6;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B5 = CLBLM_L_X10Y151_SLICE_X12Y151_BQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C1 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C2 = CLBLM_L_X10Y151_SLICE_X12Y151_CQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C3 = CLBLM_R_X11Y151_SLICE_X14Y151_AQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C5 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_C6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X13Y156_SLICE_X19Y156_D2 = 1'b1;
  assign CLBLM_R_X13Y158_SLICE_X18Y158_A4 = CLBLM_L_X12Y158_SLICE_X16Y158_AQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D1 = CLBLM_R_X5Y150_SLICE_X6Y150_AQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D2 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D3 = CLBLM_L_X10Y151_SLICE_X12Y151_DQ;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D5 = 1'b1;
  assign CLBLM_L_X10Y151_SLICE_X12Y151_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y156_SLICE_X19Y156_D5 = 1'b1;
  assign CLBLM_R_X13Y156_SLICE_X19Y156_D6 = 1'b1;
  assign CLBLM_R_X13Y158_SLICE_X18Y158_A5 = CLBLM_R_X11Y159_SLICE_X15Y159_CO5;
  assign LIOB33_X0Y173_IOB_X0Y174_O = CLBLM_L_X10Y163_SLICE_X13Y163_AO6;
  assign CLBLM_R_X13Y155_SLICE_X19Y155_A1 = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLM_R_X13Y155_SLICE_X19Y155_A2 = 1'b1;
  assign CLBLM_R_X13Y155_SLICE_X19Y155_A3 = RIOB33_X105Y131_IOB_X1Y131_I;
  assign CLBLM_R_X13Y155_SLICE_X19Y155_A4 = 1'b1;
  assign CLBLM_R_X13Y155_SLICE_X19Y155_A5 = CLBLL_L_X4Y158_SLICE_X4Y158_AO6;
  assign CLBLM_R_X13Y155_SLICE_X19Y155_A6 = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X13Y158_SLICE_X18Y158_A6 = CLBLM_R_X13Y158_SLICE_X18Y158_CO6;
  assign CLBLM_R_X13Y155_SLICE_X19Y155_B1 = 1'b1;
  assign CLBLM_R_X13Y155_SLICE_X19Y155_B2 = 1'b1;
  assign CLBLM_R_X13Y155_SLICE_X19Y155_B3 = 1'b1;
  assign CLBLM_R_X13Y155_SLICE_X19Y155_B4 = 1'b1;
  assign CLBLM_R_X13Y155_SLICE_X19Y155_B5 = 1'b1;
  assign CLBLM_R_X13Y155_SLICE_X19Y155_B6 = 1'b1;
  assign CLBLM_R_X13Y155_SLICE_X19Y155_C1 = 1'b1;
  assign CLBLM_R_X13Y155_SLICE_X19Y155_C2 = 1'b1;
  assign CLBLM_R_X13Y155_SLICE_X19Y155_C3 = 1'b1;
  assign CLBLM_R_X13Y155_SLICE_X19Y155_C4 = 1'b1;
  assign CLBLM_R_X13Y155_SLICE_X19Y155_C5 = 1'b1;
  assign CLBLM_R_X13Y155_SLICE_X19Y155_C6 = 1'b1;
  assign CLBLM_R_X13Y156_SLICE_X18Y156_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y155_SLICE_X19Y155_D1 = 1'b1;
  assign CLBLM_R_X13Y155_SLICE_X19Y155_D2 = 1'b1;
  assign CLBLM_R_X13Y155_SLICE_X19Y155_D3 = 1'b1;
  assign CLBLM_R_X13Y155_SLICE_X19Y155_D4 = 1'b1;
  assign CLBLM_R_X13Y155_SLICE_X19Y155_D5 = 1'b1;
  assign CLBLM_R_X13Y155_SLICE_X19Y155_D6 = 1'b1;
  assign RIOI3_X105Y133_ILOGIC_X1Y134_D = RIOB33_X105Y133_IOB_X1Y134_I;
  assign CLBLM_R_X11Y160_SLICE_X15Y160_C4 = 1'b1;
  assign RIOI3_X105Y133_ILOGIC_X1Y133_D = RIOB33_X105Y133_IOB_X1Y133_I;
  assign CLBLM_R_X13Y155_SLICE_X18Y155_A1 = CLBLM_R_X13Y155_SLICE_X18Y155_AQ;
  assign CLBLM_R_X13Y155_SLICE_X18Y155_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y155_SLICE_X18Y155_A3 = CLBLM_R_X7Y153_SLICE_X8Y153_AQ;
  assign CLBLM_R_X13Y155_SLICE_X18Y155_A4 = CLBLM_L_X12Y158_SLICE_X17Y158_BQ;
  assign CLBLM_R_X13Y155_SLICE_X18Y155_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y155_SLICE_X18Y155_A6 = CLBLM_L_X12Y155_SLICE_X16Y155_AO6;
  assign CLBLM_R_X11Y158_SLICE_X15Y158_C4 = CLBLM_R_X11Y159_SLICE_X14Y159_BQ;
  assign CLBLM_R_X13Y155_SLICE_X18Y155_B1 = CLBLM_L_X12Y152_SLICE_X17Y152_BO5;
  assign CLBLM_R_X13Y155_SLICE_X18Y155_B2 = CLBLM_L_X12Y156_SLICE_X17Y156_AQ;
  assign CLBLM_R_X13Y155_SLICE_X18Y155_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y155_SLICE_X18Y155_B4 = 1'b1;
  assign CLBLM_R_X11Y158_SLICE_X15Y158_C5 = CLBLM_L_X12Y158_SLICE_X16Y158_AQ;
  assign CLBLM_R_X13Y155_SLICE_X18Y155_B5 = CLBLM_L_X8Y155_SLICE_X11Y155_CQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A3 = CLBLL_L_X4Y152_SLICE_X4Y152_AQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A4 = CLBLM_R_X11Y148_SLICE_X15Y148_AQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A5 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_A6 = CLBLL_L_X4Y151_SLICE_X4Y151_CQ;
  assign CLBLM_R_X11Y158_SLICE_X15Y158_C6 = CLBLM_L_X12Y158_SLICE_X17Y158_AQ;
  assign CLBLM_R_X11Y160_SLICE_X15Y160_C5 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B3 = CLBLL_L_X4Y151_SLICE_X4Y151_BQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B4 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B5 = CLBLM_L_X10Y151_SLICE_X12Y151_CQ;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_B6 = 1'b1;
  assign CLBLM_R_X13Y155_SLICE_X18Y155_C3 = CLBLM_R_X13Y154_SLICE_X18Y154_CQ;
  assign CLBLM_R_X13Y155_SLICE_X18Y155_C4 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
  assign CLBLM_R_X13Y155_SLICE_X18Y155_C6 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C1 = CLBLL_L_X4Y150_SLICE_X5Y150_C5Q;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C2 = CLBLM_R_X5Y155_SLICE_X6Y155_DO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C4 = CLBLL_L_X4Y154_SLICE_X5Y154_BO6;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C5 = CLBLL_L_X4Y148_SLICE_X4Y148_BO5;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_C6 = CLBLL_L_X4Y149_SLICE_X5Y149_DO6;
  assign CLBLM_R_X13Y155_SLICE_X18Y155_D1 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y160_SLICE_X15Y160_C6 = 1'b1;
  assign CLBLM_R_X13Y155_SLICE_X18Y155_D2 = 1'b1;
  assign CLBLM_R_X13Y155_SLICE_X18Y155_D3 = 1'b1;
  assign CLBLM_R_X13Y155_SLICE_X18Y155_D4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X13Y155_SLICE_X18Y155_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D1 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D2 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D3 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D4 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D5 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X4Y148_D6 = 1'b1;
  assign CLBLM_R_X13Y156_SLICE_X18Y156_C1 = CLBLM_L_X12Y157_SLICE_X17Y157_BQ;
  assign CLBLM_R_X11Y158_SLICE_X15Y158_D2 = CLBLM_R_X11Y159_SLICE_X15Y159_AQ;
  assign CLBLM_R_X13Y156_SLICE_X18Y156_C2 = CLBLM_R_X11Y157_SLICE_X14Y157_AQ;
  assign CLBLM_R_X11Y158_SLICE_X15Y158_D3 = CLBLM_L_X12Y158_SLICE_X17Y158_AQ;
  assign CLBLM_R_X13Y156_SLICE_X18Y156_C3 = CLBLM_R_X11Y158_SLICE_X14Y158_AQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A1 = CLBLL_L_X4Y148_SLICE_X5Y148_AQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A2 = CLBLL_L_X4Y151_SLICE_X4Y151_BQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A3 = CLBLM_L_X10Y151_SLICE_X12Y151_CQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A5 = CLBLM_R_X11Y152_SLICE_X15Y152_DQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_A6 = CLBLL_L_X4Y150_SLICE_X5Y150_BQ;
  assign CLBLM_R_X11Y158_SLICE_X15Y158_D5 = CLBLM_L_X12Y155_SLICE_X16Y155_BO5;
  assign CLBLM_R_X13Y156_SLICE_X18Y156_C4 = CLBLM_L_X8Y154_SLICE_X10Y154_AQ;
  assign CLBLM_R_X11Y158_SLICE_X15Y158_D6 = CLBLM_L_X12Y158_SLICE_X16Y158_AQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B1 = CLBLL_L_X4Y150_SLICE_X5Y150_DQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B2 = CLBLL_L_X4Y148_SLICE_X5Y148_BQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B3 = CLBLM_L_X8Y147_SLICE_X10Y147_BQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B5 = CLBLM_R_X5Y152_SLICE_X6Y152_CO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_B6 = 1'b1;
  assign CLBLM_R_X13Y156_SLICE_X18Y156_C6 = CLBLM_L_X12Y158_SLICE_X16Y158_CO5;
  assign CLBLM_R_X13Y158_SLICE_X18Y158_B1 = CLBLM_R_X13Y158_SLICE_X18Y158_DO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C1 = CLBLM_R_X5Y148_SLICE_X7Y148_BQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C2 = CLBLL_L_X4Y148_SLICE_X5Y148_CQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C3 = 1'b1;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C5 = CLBLM_R_X5Y152_SLICE_X6Y152_CO6;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_C6 = CLBLM_L_X10Y150_SLICE_X13Y150_CQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y156_SLICE_X18Y156_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D1 = CLBLM_L_X10Y149_SLICE_X12Y149_BQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D2 = CLBLM_L_X10Y149_SLICE_X12Y149_DO5;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D3 = CLBLL_L_X4Y148_SLICE_X5Y148_DQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D5 = CLBLL_L_X4Y148_SLICE_X5Y148_AQ;
  assign CLBLL_L_X4Y148_SLICE_X5Y148_D6 = CLBLM_R_X7Y148_SLICE_X8Y148_A5Q;
  assign CLBLM_R_X13Y158_SLICE_X18Y158_B2 = CLBLM_R_X13Y158_SLICE_X18Y158_BQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A1 = CLBLM_L_X8Y152_SLICE_X11Y152_DO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A2 = CLBLM_L_X10Y149_SLICE_X13Y149_BO5;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A3 = CLBLM_L_X10Y152_SLICE_X13Y152_AQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A5 = CLBLM_L_X10Y149_SLICE_X13Y149_CO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_A6 = CLBLM_L_X10Y153_SLICE_X13Y153_CQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B1 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B3 = CLBLM_L_X10Y152_SLICE_X13Y152_AQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B4 = CLBLM_R_X5Y147_SLICE_X7Y147_BQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B5 = CLBLM_L_X12Y151_SLICE_X17Y151_AQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_B6 = 1'b1;
  assign CLBLM_R_X13Y156_SLICE_X18Y156_D1 = CLBLM_L_X12Y157_SLICE_X17Y157_BQ;
  assign CLBLM_R_X13Y156_SLICE_X18Y156_D2 = CLBLM_R_X11Y157_SLICE_X14Y157_AQ;
  assign CLBLM_R_X13Y158_SLICE_X18Y158_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C1 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C2 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C3 = CLBLM_L_X10Y148_SLICE_X13Y148_AQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C4 = CLBLM_L_X10Y155_SLICE_X12Y155_BQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C5 = CLBLM_L_X10Y148_SLICE_X13Y148_BQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_C6 = 1'b1;
  assign CLBLM_R_X13Y156_SLICE_X18Y156_D3 = CLBLM_L_X12Y156_SLICE_X17Y156_AQ;
  assign CLBLM_R_X13Y156_SLICE_X18Y156_D4 = CLBLM_L_X8Y154_SLICE_X10Y154_AQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X13Y156_SLICE_X18Y156_D5 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D2 = CLBLM_R_X11Y152_SLICE_X14Y152_DO5;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D3 = CLBLM_L_X10Y149_SLICE_X13Y149_BO5;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D4 = CLBLL_L_X4Y154_SLICE_X4Y154_BO6;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D5 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X10Y152_SLICE_X13Y152_D6 = CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  assign CLBLM_R_X13Y156_SLICE_X18Y156_D6 = CLBLM_L_X12Y158_SLICE_X16Y158_CO5;
  assign CLBLM_R_X13Y158_SLICE_X18Y158_B4 = CLBLM_R_X11Y158_SLICE_X14Y158_DO5;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A2 = CLBLM_L_X10Y153_SLICE_X12Y153_BQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A4 = CLBLM_L_X10Y149_SLICE_X12Y149_C5Q;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A5 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_A6 = CLBLM_L_X10Y152_SLICE_X13Y152_BO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B2 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B4 = CLBLM_R_X7Y153_SLICE_X9Y153_BQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B5 = 1'b1;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_B6 = CLBLM_R_X11Y149_SLICE_X15Y149_A5Q;
  assign CLBLM_R_X13Y158_SLICE_X18Y158_B5 = CLBLM_R_X11Y159_SLICE_X15Y159_CO5;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C1 = CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C2 = CLBLL_L_X4Y154_SLICE_X4Y154_BO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C3 = CLBLM_L_X10Y152_SLICE_X13Y152_BO5;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C5 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_C6 = 1'b1;
  assign CLBLM_R_X11Y158_SLICE_X14Y158_B5 = CLBLM_R_X11Y158_SLICE_X14Y158_BQ;
  assign CLBLM_R_X11Y158_SLICE_X14Y158_B6 = CLBLM_R_X7Y154_SLICE_X9Y154_CQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D1 = CLBLM_L_X10Y149_SLICE_X13Y149_AQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D2 = CLBLM_R_X3Y156_SLICE_X2Y156_DO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D3 = CLBLM_R_X7Y146_SLICE_X8Y146_AQ;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D4 = CLBLM_L_X10Y152_SLICE_X13Y152_BO6;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D5 = CLBLM_L_X10Y149_SLICE_X13Y149_BO5;
  assign CLBLM_L_X10Y152_SLICE_X12Y152_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y158_SLICE_X18Y158_B6 = CLBLM_L_X10Y158_SLICE_X13Y158_BQ;
  assign CLBLM_R_X11Y158_SLICE_X14Y158_C4 = CLBLM_R_X11Y159_SLICE_X15Y159_AQ;
  assign CLBLM_R_X11Y158_SLICE_X14Y158_C5 = CLBLM_L_X12Y158_SLICE_X17Y158_AQ;
  assign CLBLM_R_X13Y156_SLICE_X19Y156_A1 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_R_X13Y156_SLICE_X19Y156_A3 = CLBLM_R_X13Y156_SLICE_X19Y156_AQ;
  assign CLBLM_R_X13Y156_SLICE_X19Y156_A4 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X13Y156_SLICE_X19Y156_A5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y158_SLICE_X14Y158_C6 = CLBLM_R_X11Y159_SLICE_X14Y159_BQ;
  assign CLBLM_R_X13Y156_SLICE_X19Y156_A6 = 1'b1;
  assign CLBLM_R_X13Y156_SLICE_X19Y156_A2 = CLBLM_R_X7Y154_SLICE_X8Y154_BQ;
  assign CLBLM_R_X13Y156_SLICE_X19Y156_B1 = 1'b1;
  assign CLBLM_R_X13Y156_SLICE_X19Y156_B2 = 1'b1;
  assign CLBLM_R_X13Y156_SLICE_X19Y156_B3 = 1'b1;
  assign CLBLM_R_X13Y156_SLICE_X19Y156_B4 = 1'b1;
  assign CLBLM_R_X13Y156_SLICE_X19Y156_B5 = 1'b1;
  assign CLBLM_R_X13Y156_SLICE_X19Y156_B6 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A2 = CLBLM_L_X10Y147_SLICE_X12Y147_AQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A3 = CLBLM_R_X11Y146_SLICE_X15Y146_AQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A4 = CLBLM_R_X7Y146_SLICE_X9Y146_DO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A5 = CLBLM_L_X12Y147_SLICE_X16Y147_AQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_A6 = 1'b1;
  assign CLBLM_R_X13Y156_SLICE_X19Y156_C1 = 1'b1;
  assign CLBLM_R_X13Y156_SLICE_X19Y156_C2 = 1'b1;
  assign CLBLM_R_X13Y156_SLICE_X19Y156_C3 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B2 = CLBLM_R_X11Y146_SLICE_X15Y146_BQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B3 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B4 = CLBLM_R_X7Y146_SLICE_X8Y146_DO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B5 = CLBLM_L_X8Y146_SLICE_X11Y146_CQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_B6 = CLBLM_R_X11Y153_SLICE_X15Y153_BQ;
  assign CLBLM_R_X13Y156_SLICE_X19Y156_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X13Y156_SLICE_X19Y156_D1 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C1 = CLBLM_R_X11Y154_SLICE_X15Y154_BQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C2 = CLBLM_R_X11Y146_SLICE_X15Y146_CQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C4 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C5 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_C6 = CLBLM_L_X8Y146_SLICE_X11Y146_AQ;
  assign CLBLM_R_X13Y156_SLICE_X19Y156_D3 = 1'b1;
  assign CLBLM_R_X13Y156_SLICE_X19Y156_D4 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y156_SLICE_X18Y156_A1 = 1'b1;
  assign CLBLM_R_X13Y156_SLICE_X18Y156_A2 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X13Y156_SLICE_X18Y156_A3 = CLBLM_R_X13Y156_SLICE_X18Y156_AQ;
  assign CLBLM_R_X13Y156_SLICE_X18Y156_A4 = CLBLM_R_X13Y157_SLICE_X19Y157_AQ;
  assign CLBLM_R_X13Y156_SLICE_X18Y156_A5 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D1 = CLBLM_L_X10Y145_SLICE_X13Y145_CQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D2 = CLBLM_L_X10Y145_SLICE_X13Y145_BQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D3 = CLBLM_L_X10Y146_SLICE_X12Y146_C5Q;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D4 = CLBLM_L_X10Y147_SLICE_X12Y147_CQ;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D5 = CLBLM_L_X10Y146_SLICE_X12Y146_CQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A1 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A3 = CLBLL_L_X4Y149_SLICE_X4Y149_AQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A4 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A5 = CLBLM_L_X10Y146_SLICE_X12Y146_CQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_A6 = CLBLL_L_X4Y149_SLICE_X4Y149_CO6;
  assign CLBLM_R_X11Y146_SLICE_X15Y146_D6 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_AX = CLBLL_L_X4Y148_SLICE_X4Y148_BO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A1 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B1 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B2 = CLBLL_L_X4Y149_SLICE_X4Y149_BQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B3 = CLBLL_L_X4Y151_SLICE_X4Y151_C5Q;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B5 = CLBLM_R_X11Y148_SLICE_X15Y148_AQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A2 = CLBLM_R_X11Y148_SLICE_X14Y148_AQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A3 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C1 = CLBLL_L_X4Y152_SLICE_X4Y152_AQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C3 = LIOB33_X0Y53_IOB_X0Y53_I;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C4 = CLBLL_L_X4Y151_SLICE_X4Y151_CQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_C6 = CLBLM_R_X5Y149_SLICE_X6Y149_A5Q;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B1 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B2 = CLBLM_R_X11Y146_SLICE_X14Y146_BQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_B5 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D1 = CLBLL_L_X4Y151_SLICE_X4Y151_C5Q;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D2 = CLBLM_R_X3Y151_SLICE_X2Y151_AQ;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D4 = CLBLM_R_X5Y149_SLICE_X6Y149_B5Q;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D5 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X4Y149_D6 = CLBLM_L_X10Y154_SLICE_X13Y154_CQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C3 = CLBLM_R_X13Y147_SLICE_X18Y147_CO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_C6 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D1 = 1'b1;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D2 = CLBLM_L_X10Y147_SLICE_X13Y147_BQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D3 = CLBLM_R_X11Y146_SLICE_X14Y146_DQ;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D4 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y146_SLICE_X14Y146_D6 = CLBLM_R_X11Y146_SLICE_X15Y146_BQ;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_D1 = CLBLL_L_X2Y140_SLICE_X0Y140_AO5;
  assign LIOI3_SING_X0Y100_OLOGIC_X0Y100_T1 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A1 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A2 = CLBLM_R_X7Y153_SLICE_X8Y153_AQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A3 = CLBLL_L_X4Y149_SLICE_X5Y149_AQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A5 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_A6 = LIOB33_X0Y79_IOB_X0Y79_I;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_AX = CLBLL_L_X4Y149_SLICE_X5Y149_BO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B2 = CLBLL_L_X4Y150_SLICE_X5Y150_AQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B3 = RIOB33_X105Y127_IOB_X1Y127_I;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B4 = CLBLM_R_X5Y149_SLICE_X6Y149_DO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B5 = CLBLL_L_X4Y150_SLICE_X5Y150_BQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_B6 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C1 = CLBLM_R_X7Y153_SLICE_X8Y153_AQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C2 = CLBLM_L_X8Y148_SLICE_X11Y148_BQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C3 = CLBLL_L_X4Y150_SLICE_X5Y150_C5Q;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C4 = CLBLL_L_X4Y151_SLICE_X5Y151_CQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_C6 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D3 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D4 = 1'b1;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D1 = CLBLL_L_X4Y149_SLICE_X5Y149_CO5;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D2 = CLBLM_R_X3Y155_SLICE_X2Y155_BO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D3 = CLBLL_L_X4Y154_SLICE_X5Y154_CO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D4 = CLBLL_L_X4Y147_SLICE_X5Y147_AQ;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D5 = CLBLL_L_X4Y153_SLICE_X4Y153_BO6;
  assign CLBLL_L_X4Y149_SLICE_X5Y149_D6 = CLBLM_L_X10Y149_SLICE_X13Y149_A5Q;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D5 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X163Y174_D6 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A2 = CLBLM_R_X5Y153_SLICE_X6Y153_AQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A3 = CLBLM_L_X10Y153_SLICE_X13Y153_AQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A5 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_A6 = CLBLM_R_X11Y157_SLICE_X14Y157_CQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B3 = CLBLM_R_X11Y153_SLICE_X14Y153_AQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B4 = CLBLL_L_X4Y155_SLICE_X4Y155_AQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B5 = CLBLM_L_X10Y151_SLICE_X13Y151_BQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_B6 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C2 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C4 = CLBLM_R_X11Y154_SLICE_X14Y154_CQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C5 = CLBLM_L_X10Y153_SLICE_X13Y153_BO5;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_C6 = CLBLM_R_X7Y153_SLICE_X9Y153_AQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D1 = CLBLM_L_X10Y156_SLICE_X12Y156_AQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D2 = CLBLM_L_X10Y151_SLICE_X13Y151_CQ;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D3 = CLBLM_L_X12Y153_SLICE_X16Y153_BO5;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D4 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y153_SLICE_X13Y153_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_A5 = 1'b1;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_D1 = LIOB33_X0Y67_IOB_X0Y68_I;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A2 = CLBLM_L_X10Y155_SLICE_X12Y155_AQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A3 = CLBLM_L_X10Y153_SLICE_X12Y153_AQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A4 = CLBLM_R_X7Y155_SLICE_X8Y155_CO6;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A5 = CLBLM_L_X10Y147_SLICE_X12Y147_DQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_A6 = CLBLM_R_X7Y158_SLICE_X8Y158_CO5;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B2 = CLBLM_R_X11Y152_SLICE_X14Y152_DO5;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B4 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B5 = CLBLM_R_X5Y150_SLICE_X6Y150_AQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_B6 = CLBLM_L_X12Y154_SLICE_X17Y154_A5Q;
  assign LIOI3_X0Y153_OLOGIC_X0Y154_T1 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_D1 = CLBLM_L_X16Y156_SLICE_X22Y156_AO5;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C1 = CLBLM_R_X13Y149_SLICE_X18Y149_A5Q;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C2 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C3 = CLBLM_L_X10Y154_SLICE_X12Y154_DQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C4 = CLBLM_R_X11Y149_SLICE_X15Y149_A5Q;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C5 = CLBLM_R_X11Y153_SLICE_X15Y153_AQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_C6 = CLBLM_R_X7Y154_SLICE_X8Y154_AO5;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_D1 = LIOB33_X0Y67_IOB_X0Y67_I;
  assign RIOI3_X105Y197_OLOGIC_X1Y198_T1 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign LIOI3_X0Y153_OLOGIC_X0Y153_T1 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D1 = CLBLM_L_X10Y152_SLICE_X12Y152_AQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D2 = CLBLL_L_X4Y153_SLICE_X5Y153_AQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D4 = CLBLM_L_X10Y153_SLICE_X12Y153_BQ;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D5 = 1'b1;
  assign CLBLM_L_X10Y153_SLICE_X12Y153_D6 = CLBLM_L_X10Y150_SLICE_X13Y150_CQ;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B3 = 1'b1;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B4 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_D1 = CLBLM_L_X16Y156_SLICE_X22Y156_AO5;
  assign CLBLM_R_X103Y174_SLICE_X162Y174_B5 = 1'b1;
  assign RIOI3_X105Y197_OLOGIC_X1Y197_T1 = 1'b1;
  assign CLBLM_R_X13Y157_SLICE_X19Y157_A1 = CLBLM_R_X13Y154_SLICE_X18Y154_CQ;
  assign CLBLM_R_X13Y157_SLICE_X19Y157_A2 = CLBLM_R_X11Y158_SLICE_X14Y158_DO5;
  assign CLBLM_R_X13Y157_SLICE_X19Y157_A3 = CLBLM_R_X13Y157_SLICE_X18Y157_CO6;
  assign CLBLM_R_X13Y157_SLICE_X19Y157_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y157_SLICE_X19Y157_A5 = CLBLM_R_X11Y159_SLICE_X15Y159_CO5;
  assign CLBLM_R_X13Y157_SLICE_X19Y157_A6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_D1 = CLBLM_R_X103Y169_SLICE_X163Y169_AO5;
  assign CLBLM_R_X13Y157_SLICE_X19Y157_B1 = CLBLM_R_X13Y159_SLICE_X18Y159_CO6;
  assign CLBLM_R_X13Y157_SLICE_X19Y157_B2 = CLBLM_R_X11Y157_SLICE_X15Y157_BQ;
  assign CLBLM_R_X13Y157_SLICE_X19Y157_B3 = CLBLM_R_X11Y157_SLICE_X14Y157_AQ;
  assign CLBLM_R_X13Y157_SLICE_X19Y157_B4 = 1'b1;
  assign CLBLM_R_X13Y157_SLICE_X19Y157_B5 = CLBLM_R_X11Y158_SLICE_X14Y158_AQ;
  assign CLBLM_R_X13Y157_SLICE_X19Y157_B6 = CLBLM_R_X13Y158_SLICE_X18Y158_BQ;
  assign RIOI3_TBYTESRC_X105Y169_OLOGIC_X1Y170_T1 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A1 = CLBLM_R_X11Y152_SLICE_X14Y152_B5Q;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A2 = CLBLM_R_X11Y146_SLICE_X15Y146_DO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A3 = CLBLM_R_X11Y147_SLICE_X14Y147_AO5;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A4 = CLBLM_R_X7Y146_SLICE_X8Y146_BO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A5 = CLBLM_L_X8Y155_SLICE_X10Y155_BQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_A6 = CLBLM_R_X3Y154_SLICE_X2Y154_AO6;
  assign CLBLM_R_X13Y157_SLICE_X19Y157_C1 = 1'b1;
  assign CLBLM_R_X13Y157_SLICE_X19Y157_C2 = 1'b1;
  assign CLBLM_R_X13Y157_SLICE_X19Y157_C3 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B1 = CLBLM_L_X10Y150_SLICE_X13Y150_C5Q;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B2 = CLBLM_L_X10Y147_SLICE_X13Y147_AQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B3 = CLBLM_R_X11Y153_SLICE_X15Y153_DQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B4 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B5 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_B6 = CLBLM_L_X12Y147_SLICE_X16Y147_BO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D3 = CLBLM_R_X11Y157_SLICE_X14Y157_DO6;
  assign CLBLM_R_X13Y157_SLICE_X19Y157_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C1 = CLBLM_R_X11Y146_SLICE_X15Y146_CQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C2 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C3 = CLBLM_L_X10Y150_SLICE_X13Y150_C5Q;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C4 = CLBLM_L_X10Y147_SLICE_X13Y147_BQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C5 = CLBLM_R_X11Y147_SLICE_X15Y147_DO6;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_C6 = CLBLM_L_X8Y155_SLICE_X10Y155_BQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D5 = CLBLM_R_X7Y146_SLICE_X9Y146_BO6;
  assign CLBLM_R_X13Y157_SLICE_X19Y157_D4 = 1'b1;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_A1 = CLBLM_L_X12Y157_SLICE_X16Y157_A5Q;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D6 = CLBLM_R_X7Y146_SLICE_X8Y146_BO6;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_A2 = 1'b1;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y157_SLICE_X18Y157_A4 = RIOB33_X105Y143_IOB_X1Y143_I;
  assign CLBLM_R_X13Y156_SLICE_X18Y156_B1 = CLBLM_R_X13Y156_SLICE_X18Y156_DO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A1 = CLBLM_R_X11Y149_SLICE_X14Y149_CQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A2 = CLBLL_L_X4Y150_SLICE_X4Y150_BQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A3 = CLBLL_L_X4Y150_SLICE_X4Y150_AQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A4 = CLBLL_L_X4Y151_SLICE_X4Y151_BQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A5 = CLBLM_L_X10Y151_SLICE_X12Y151_CQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D1 = CLBLM_L_X8Y146_SLICE_X11Y146_AQ;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D2 = CLBLM_L_X8Y148_SLICE_X11Y148_B5Q;
  assign CLBLM_R_X11Y147_SLICE_X15Y147_D3 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B1 = CLBLM_L_X8Y150_SLICE_X10Y150_DO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B2 = CLBLL_L_X4Y150_SLICE_X4Y150_BQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B3 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B4 = CLBLM_R_X3Y150_SLICE_X3Y150_AQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A4 = CLBLM_L_X10Y145_SLICE_X13Y145_BQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A5 = CLBLM_L_X10Y145_SLICE_X13Y145_CQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_A6 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C1 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C2 = CLBLM_R_X7Y151_SLICE_X9Y151_BQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C3 = CLBLM_R_X5Y148_SLICE_X7Y148_B5Q;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C5 = CLBLM_L_X8Y150_SLICE_X10Y150_DO6;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B1 = CLBLM_R_X13Y147_SLICE_X18Y147_AO5;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B2 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B3 = CLBLM_L_X10Y147_SLICE_X12Y147_BQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B4 = CLBLM_R_X11Y150_SLICE_X14Y150_AQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B5 = CLBLM_R_X11Y147_SLICE_X14Y147_AO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_B6 = CLBLM_L_X10Y149_SLICE_X12Y149_CQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D1 = CLBLM_L_X8Y148_SLICE_X11Y148_BQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D2 = CLBLL_L_X4Y150_SLICE_X5Y150_C5Q;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D3 = CLBLL_L_X4Y151_SLICE_X5Y151_CQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D5 = CLBLM_R_X7Y153_SLICE_X8Y153_AQ;
  assign CLBLL_L_X4Y150_SLICE_X4Y150_D6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C1 = CLBLM_L_X12Y149_SLICE_X16Y149_B5Q;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C2 = CLBLM_R_X11Y147_SLICE_X15Y147_CO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C3 = CLBLM_R_X13Y153_SLICE_X18Y153_CQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C4 = CLBLM_L_X8Y147_SLICE_X11Y147_AQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C5 = CLBLM_R_X11Y147_SLICE_X14Y147_DO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_C6 = CLBLM_L_X10Y147_SLICE_X13Y147_DO6;
  assign CLBLM_R_X13Y156_SLICE_X18Y156_B3 = CLBLM_R_X11Y159_SLICE_X15Y159_CO5;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D1 = CLBLM_R_X11Y146_SLICE_X15Y146_AQ;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D2 = CLBLM_L_X10Y146_SLICE_X13Y146_DO6;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D3 = CLBLM_R_X11Y152_SLICE_X14Y152_B5Q;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D4 = CLBLM_L_X12Y157_SLICE_X17Y157_A5Q;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D5 = 1'b1;
  assign CLBLM_R_X11Y147_SLICE_X14Y147_D6 = CLBLM_L_X10Y147_SLICE_X12Y147_AQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A1 = CLBLM_R_X5Y152_SLICE_X7Y152_CQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A2 = CLBLL_L_X4Y150_SLICE_X5Y150_BQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A3 = CLBLL_L_X4Y150_SLICE_X5Y150_AQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A4 = CLBLM_L_X10Y149_SLICE_X12Y149_DO5;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A5 = CLBLM_R_X5Y149_SLICE_X6Y149_DO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y156_SLICE_X18Y156_B4 = CLBLM_L_X12Y158_SLICE_X16Y158_BO5;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B1 = 1'b1;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B2 = CLBLL_L_X4Y150_SLICE_X5Y150_BQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B3 = CLBLM_R_X5Y149_SLICE_X6Y149_DO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B4 = CLBLM_L_X10Y149_SLICE_X12Y149_DO5;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B5 = CLBLM_R_X5Y157_SLICE_X6Y157_AQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C1 = CLBLM_L_X12Y155_SLICE_X16Y155_CO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C2 = CLBLM_R_X13Y151_SLICE_X18Y151_AQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C3 = CLBLM_R_X5Y155_SLICE_X6Y155_DO6;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C5 = CLBLL_L_X4Y149_SLICE_X4Y149_A5Q;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_C6 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B2 = CLBLM_R_X11Y148_SLICE_X14Y148_BQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X13Y156_SLICE_X18Y156_B5 = CLBLM_R_X11Y158_SLICE_X15Y158_DO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B3 = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1 = LIOB33_X0Y61_IOB_X0Y62_I;
  assign RIOI3_X105Y135_ILOGIC_X1Y136_D = RIOB33_X105Y135_IOB_X1Y136_I;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D1 = CLBLL_L_X4Y155_SLICE_X5Y155_AQ;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D4 = CLBLL_L_X4Y149_SLICE_X4Y149_A5Q;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D5 = CLBLM_R_X5Y148_SLICE_X6Y148_A5Q;
  assign CLBLL_L_X4Y150_SLICE_X5Y150_D6 = 1'b1;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1 = 1'b1;
  assign RIOI3_X105Y135_ILOGIC_X1Y135_D = RIOB33_X105Y135_IOB_X1Y135_I;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y156_SLICE_X18Y156_B6 = CLBLM_R_X11Y158_SLICE_X14Y158_AQ;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_A1 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_A2 = CLBLM_L_X10Y154_SLICE_X13Y154_BQ;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_A3 = CLBLM_R_X11Y153_SLICE_X15Y153_AQ;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_A5 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_A6 = 1'b1;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_B1 = 1'b1;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_B3 = CLBLM_L_X8Y150_SLICE_X10Y150_A5Q;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_B5 = CLBLM_L_X8Y154_SLICE_X10Y154_AQ;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_B6 = 1'b1;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_C1 = CLBLM_L_X12Y154_SLICE_X17Y154_AQ;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_C3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_C4 = CLBLM_L_X8Y154_SLICE_X10Y154_C5Q;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_C5 = CLBLM_L_X10Y154_SLICE_X13Y154_C5Q;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_C6 = 1'b1;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_D1 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_D2 = CLBLM_R_X7Y152_SLICE_X9Y152_CO6;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_D3 = CLBLM_L_X10Y154_SLICE_X13Y154_DQ;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_D5 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y154_SLICE_X13Y154_D6 = CLBLM_R_X5Y152_SLICE_X6Y152_AQ;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_A1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_A2 = CLBLM_R_X11Y154_SLICE_X14Y154_AQ;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_A3 = CLBLM_L_X10Y154_SLICE_X12Y154_AQ;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_A4 = 1'b1;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_A5 = CLBLM_L_X10Y156_SLICE_X12Y156_AQ;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_A6 = CLBLM_R_X7Y153_SLICE_X9Y153_CO6;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_AX = CLBLM_L_X10Y154_SLICE_X12Y154_BO6;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_B1 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_B2 = CLBLM_L_X10Y154_SLICE_X12Y154_A5Q;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_B3 = CLBLM_R_X7Y153_SLICE_X8Y153_AQ;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_B4 = CLBLM_R_X11Y153_SLICE_X14Y153_AQ;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_B6 = 1'b1;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_C1 = CLBLM_R_X11Y159_SLICE_X15Y159_CO6;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_C2 = 1'b1;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_C3 = 1'b1;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_C4 = CLBLL_L_X4Y150_SLICE_X5Y150_C5Q;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_C6 = CLBLM_L_X8Y153_SLICE_X11Y153_BQ;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_D2 = CLBLM_L_X10Y154_SLICE_X13Y154_AO5;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_D3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_D4 = CLBLM_L_X8Y155_SLICE_X11Y155_BQ;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_D5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y154_SLICE_X12Y154_D6 = CLBLM_L_X10Y154_SLICE_X12Y154_CQ;
  assign LIOB33_X0Y145_IOB_X0Y146_O = LIOB33_X0Y59_IOB_X0Y59_I;
  assign LIOB33_X0Y145_IOB_X0Y145_O = LIOB33_X0Y57_IOB_X0Y58_I;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X13Y158_SLICE_X19Y158_A1 = CLBLM_L_X12Y156_SLICE_X17Y156_AQ;
  assign CLBLM_R_X13Y158_SLICE_X19Y158_A2 = CLBLM_L_X12Y158_SLICE_X16Y158_CO5;
  assign CLBLM_R_X13Y158_SLICE_X19Y158_A3 = CLBLM_L_X12Y157_SLICE_X17Y157_BQ;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_C5 = CLBLM_R_X5Y157_SLICE_X7Y157_DQ;
  assign CLBLM_R_X13Y158_SLICE_X19Y158_A4 = CLBLM_L_X8Y154_SLICE_X10Y154_AQ;
  assign CLBLM_R_X13Y158_SLICE_X19Y158_A5 = CLBLM_R_X11Y158_SLICE_X14Y158_AQ;
  assign CLBLM_R_X13Y158_SLICE_X19Y158_A6 = CLBLM_R_X11Y157_SLICE_X14Y157_AQ;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X13Y158_SLICE_X19Y158_B1 = CLBLM_L_X12Y156_SLICE_X17Y156_AQ;
  assign CLBLM_R_X13Y158_SLICE_X19Y158_B2 = CLBLM_L_X12Y158_SLICE_X16Y158_CO5;
  assign CLBLM_R_X13Y158_SLICE_X19Y158_B3 = CLBLM_L_X12Y157_SLICE_X17Y157_BQ;
  assign CLBLM_R_X13Y158_SLICE_X19Y158_B4 = CLBLM_L_X8Y154_SLICE_X10Y154_AQ;
  assign CLBLM_R_X13Y158_SLICE_X19Y158_B5 = CLBLM_R_X11Y158_SLICE_X14Y158_AQ;
  assign CLBLM_R_X13Y158_SLICE_X19Y158_B6 = CLBLM_R_X11Y157_SLICE_X14Y157_AQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A1 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A3 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A4 = CLBLM_R_X11Y148_SLICE_X15Y148_BO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A5 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_A6 = CLBLM_R_X13Y151_SLICE_X18Y151_DQ;
  assign CLBLM_R_X13Y158_SLICE_X19Y158_C1 = 1'b1;
  assign CLBLM_R_X13Y158_SLICE_X19Y158_C2 = 1'b1;
  assign CLBLM_R_X13Y158_SLICE_X19Y158_C3 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B1 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B2 = CLBLM_L_X12Y148_SLICE_X16Y148_AO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B3 = CLBLM_R_X11Y148_SLICE_X15Y148_AQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B4 = CLBLM_L_X10Y146_SLICE_X12Y146_CQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B5 = CLBLM_L_X12Y149_SLICE_X16Y149_B5Q;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_B6 = CLBLM_L_X10Y145_SLICE_X12Y145_CQ;
  assign CLBLM_R_X13Y158_SLICE_X19Y158_D1 = 1'b1;
  assign CLBLM_R_X13Y158_SLICE_X19Y158_D2 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C1 = CLBLM_R_X7Y148_SLICE_X9Y148_CO5;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C2 = CLBLM_L_X12Y156_SLICE_X16Y156_CO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C3 = CLBLM_R_X7Y146_SLICE_X9Y146_BO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C4 = CLBLM_L_X8Y148_SLICE_X11Y148_B5Q;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C5 = CLBLM_R_X11Y156_SLICE_X15Y156_CO6;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_C6 = CLBLM_R_X7Y146_SLICE_X8Y146_BO6;
  assign CLBLM_R_X13Y158_SLICE_X19Y158_D3 = 1'b1;
  assign CLBLM_R_X13Y158_SLICE_X19Y158_D4 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X13Y158_SLICE_X18Y158_A1 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A1 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A3 = CLBLL_L_X4Y151_SLICE_X4Y151_AQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A4 = CLBLM_R_X13Y150_SLICE_X18Y150_CQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A5 = CLBLL_L_X4Y152_SLICE_X4Y152_AQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_A6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D1 = CLBLM_R_X11Y150_SLICE_X14Y150_AQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D2 = CLBLM_R_X7Y148_SLICE_X9Y148_CO5;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B1 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B3 = CLBLM_L_X10Y151_SLICE_X12Y151_CQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B4 = CLBLL_L_X4Y151_SLICE_X4Y151_D5Q;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B5 = CLBLL_L_X4Y150_SLICE_X5Y150_D5Q;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_B6 = 1'b1;
  assign CLBLM_R_X5Y152_SLICE_X7Y152_D2 = CLBLM_L_X10Y152_SLICE_X12Y152_AQ;
  assign CLBLM_R_X11Y148_SLICE_X15Y148_D4 = CLBLM_L_X12Y152_SLICE_X16Y152_DO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A1 = CLBLM_R_X11Y148_SLICE_X14Y148_CQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C1 = CLBLL_L_X4Y152_SLICE_X4Y152_AQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C2 = CLBLM_R_X5Y151_SLICE_X7Y151_BQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C3 = CLBLM_R_X3Y151_SLICE_X2Y151_AQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C4 = CLBLL_L_X4Y158_SLICE_X5Y158_AQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C5 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_C6 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A3 = CLBLM_R_X11Y148_SLICE_X14Y148_AQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A5 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_A6 = CLBLM_L_X8Y150_SLICE_X11Y150_AQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B1 = CLBLM_L_X10Y150_SLICE_X13Y150_C5Q;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D1 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D2 = CLBLM_R_X3Y155_SLICE_X2Y155_BO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D3 = CLBLM_L_X10Y149_SLICE_X12Y149_BQ;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D5 = CLBLL_L_X4Y154_SLICE_X5Y154_BO6;
  assign CLBLL_L_X4Y151_SLICE_X4Y151_D6 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_B5 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C1 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C2 = CLBLM_L_X10Y144_SLICE_X12Y144_AQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C3 = RIOB33_X105Y141_IOB_X1Y142_I;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C4 = CLBLM_L_X10Y151_SLICE_X12Y151_DQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C5 = CLBLM_R_X11Y148_SLICE_X14Y148_DO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_C6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D1 = CLBLM_R_X11Y152_SLICE_X14Y152_B5Q;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D2 = CLBLM_R_X11Y148_SLICE_X14Y148_CQ;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D3 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D4 = CLBLM_R_X11Y146_SLICE_X15Y146_DO6;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D5 = 1'b1;
  assign CLBLM_R_X11Y148_SLICE_X14Y148_D6 = CLBLM_R_X7Y146_SLICE_X8Y146_CO6;
  assign CLBLM_R_X13Y156_SLICE_X18Y156_C5 = CLBLM_L_X12Y156_SLICE_X17Y156_AQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A1 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A2 = CLBLM_R_X7Y151_SLICE_X9Y151_BQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A3 = CLBLL_L_X4Y151_SLICE_X5Y151_AQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A5 = CLBLM_L_X12Y151_SLICE_X16Y151_C5Q;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_A6 = CLBLM_R_X5Y152_SLICE_X6Y152_CO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B1 = CLBLM_L_X12Y149_SLICE_X16Y149_DQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B2 = CLBLL_L_X4Y151_SLICE_X5Y151_BQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B3 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B4 = CLBLM_L_X8Y150_SLICE_X11Y150_AQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B5 = CLBLM_R_X5Y152_SLICE_X6Y152_CO5;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_A3 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_A4 = CLBLM_R_X5Y152_SLICE_X7Y152_BQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C1 = CLBLM_R_X7Y151_SLICE_X9Y151_C5Q;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C3 = CLBLL_L_X4Y156_SLICE_X4Y156_AQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C4 = CLBLM_R_X3Y150_SLICE_X3Y150_AQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C5 = CLBLM_R_X3Y151_SLICE_X3Y151_AQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_C6 = CLBLM_R_X3Y150_SLICE_X3Y150_BQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_A5 = 1'b1;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D1 = CLBLM_R_X5Y147_SLICE_X6Y147_BQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D2 = CLBLL_L_X2Y153_SLICE_X1Y153_AO5;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D3 = CLBLL_L_X4Y157_SLICE_X4Y157_BO6;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D4 = CLBLL_L_X4Y152_SLICE_X5Y152_BQ;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D5 = LIOB33_X0Y65_IOB_X0Y65_I;
  assign CLBLL_L_X4Y151_SLICE_X5Y151_D6 = CLBLM_R_X3Y151_SLICE_X2Y151_CO5;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_A1 = CLBLM_L_X10Y155_SLICE_X13Y155_AQ;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_A2 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_A3 = CLBLM_R_X11Y149_SLICE_X14Y149_AQ;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_A4 = CLBLM_L_X8Y150_SLICE_X10Y150_AQ;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_A6 = 1'b1;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_B1 = CLBLM_R_X5Y157_SLICE_X7Y157_AQ;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_B2 = CLBLM_L_X10Y155_SLICE_X13Y155_BQ;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_B3 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_B4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_B5 = CLBLM_L_X10Y150_SLICE_X13Y150_DO6;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_B6 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_D1 = LIOB33_X0Y63_IOB_X0Y63_I;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_C1 = CLBLM_L_X8Y152_SLICE_X11Y152_AO6;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_C2 = CLBLM_R_X7Y153_SLICE_X9Y153_CO6;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_C3 = CLBLM_R_X11Y152_SLICE_X14Y152_AQ;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_C4 = CLBLM_L_X8Y156_SLICE_X11Y156_DO6;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_C5 = CLBLM_L_X8Y153_SLICE_X11Y153_CQ;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_C6 = CLBLM_L_X10Y155_SLICE_X13Y155_DO6;
  assign LIOI3_SING_X0Y150_OLOGIC_X0Y150_T1 = 1'b1;
  assign LIOI3_SING_X0Y199_OLOGIC_X0Y199_D1 = LIOB33_X0Y73_IOB_X0Y74_I;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_CLK = CLK_HROW_TOP_R_X139Y182_BUFHCE_X0Y44_O;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_D1 = CLBLM_L_X10Y155_SLICE_X13Y155_BQ;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_D2 = CLBLM_R_X7Y154_SLICE_X8Y154_AO5;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_D3 = CLBLM_L_X10Y156_SLICE_X13Y156_AO5;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_D4 = CLBLM_L_X10Y156_SLICE_X13Y156_CO6;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_D5 = CLBLM_R_X11Y153_SLICE_X14Y153_DO6;
  assign CLBLM_L_X10Y155_SLICE_X13Y155_D6 = CLBLM_L_X10Y152_SLICE_X13Y152_CO5;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_A1 = CLBLM_R_X11Y146_SLICE_X14Y146_DQ;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_A2 = CLBLM_R_X7Y155_SLICE_X8Y155_CO6;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_A3 = CLBLM_L_X10Y155_SLICE_X12Y155_AQ;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_A4 = CLBLM_R_X7Y157_SLICE_X9Y157_AQ;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_A5 = CLBLM_R_X7Y158_SLICE_X8Y158_CO5;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_A6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_C3 = RIOB33_X105Y121_IOB_X1Y121_I;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_B1 = CLBLM_L_X10Y155_SLICE_X12Y155_CQ;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_B2 = CLBLM_L_X10Y155_SLICE_X12Y155_BQ;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_B3 = CLBLM_R_X11Y146_SLICE_X14Y146_AQ;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_B4 = RIOB33_X105Y117_IOB_X1Y118_I;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_B5 = CLBLM_R_X7Y149_SLICE_X9Y149_AQ;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_B6 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_C4 = CLBLM_R_X5Y154_SLICE_X6Y154_AQ;
  assign CLBLM_R_X5Y152_SLICE_X6Y152_C5 = CLBLM_L_X12Y149_SLICE_X16Y149_CQ;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_C2 = 1'b1;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_C3 = CLBLM_L_X10Y148_SLICE_X12Y148_BO5;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_C4 = LIOB33_X0Y77_IOB_X0Y77_I;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_C5 = CLBLM_L_X10Y156_SLICE_X13Y156_BQ;
  assign CLBLM_L_X10Y155_SLICE_X12Y155_C6 = CLBLM_R_X7Y149_SLICE_X8Y149_AQ;
endmodule
