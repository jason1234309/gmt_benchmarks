module top(
  input LIOB33_SING_X0Y100_IOB_X0Y100_IPAD,
  input LIOB33_X0Y101_IOB_X0Y101_IPAD,
  input LIOB33_X0Y101_IOB_X0Y102_IPAD,
  input LIOB33_X0Y103_IOB_X0Y103_IPAD,
  input LIOB33_X0Y103_IOB_X0Y104_IPAD,
  input LIOB33_X0Y105_IOB_X0Y105_IPAD,
  input LIOB33_X0Y105_IOB_X0Y106_IPAD,
  input LIOB33_X0Y107_IOB_X0Y107_IPAD,
  input LIOB33_X0Y107_IOB_X0Y108_IPAD,
  input LIOB33_X0Y109_IOB_X0Y109_IPAD,
  input LIOB33_X0Y109_IOB_X0Y110_IPAD,
  input LIOB33_X0Y111_IOB_X0Y111_IPAD,
  input LIOB33_X0Y111_IOB_X0Y112_IPAD,
  input LIOB33_X0Y113_IOB_X0Y113_IPAD,
  input LIOB33_X0Y113_IOB_X0Y114_IPAD,
  input LIOB33_X0Y115_IOB_X0Y115_IPAD,
  input LIOB33_X0Y115_IOB_X0Y116_IPAD,
  input LIOB33_X0Y117_IOB_X0Y117_IPAD,
  input RIOB33_SING_X105Y100_IOB_X1Y100_IPAD,
  input RIOB33_X105Y101_IOB_X1Y101_IPAD,
  input RIOB33_X105Y101_IOB_X1Y102_IPAD,
  input RIOB33_X105Y103_IOB_X1Y103_IPAD,
  input RIOB33_X105Y103_IOB_X1Y104_IPAD,
  input RIOB33_X105Y105_IOB_X1Y105_IPAD,
  input RIOB33_X105Y105_IOB_X1Y106_IPAD,
  input RIOB33_X105Y107_IOB_X1Y107_IPAD,
  input RIOB33_X105Y107_IOB_X1Y108_IPAD,
  input RIOB33_X105Y109_IOB_X1Y109_IPAD,
  input RIOB33_X105Y109_IOB_X1Y110_IPAD,
  input RIOB33_X105Y111_IOB_X1Y111_IPAD,
  input RIOB33_X105Y111_IOB_X1Y112_IPAD,
  input RIOB33_X105Y113_IOB_X1Y113_IPAD,
  output LIOB33_SING_X0Y149_IOB_X0Y149_OPAD,
  output LIOB33_X0Y117_IOB_X0Y118_OPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD,
  output LIOB33_X0Y125_IOB_X0Y125_OPAD,
  output LIOB33_X0Y125_IOB_X0Y126_OPAD,
  output LIOB33_X0Y127_IOB_X0Y127_OPAD,
  output LIOB33_X0Y127_IOB_X0Y128_OPAD,
  output LIOB33_X0Y129_IOB_X0Y129_OPAD,
  output LIOB33_X0Y129_IOB_X0Y130_OPAD,
  output LIOB33_X0Y131_IOB_X0Y131_OPAD,
  output LIOB33_X0Y131_IOB_X0Y132_OPAD,
  output LIOB33_X0Y133_IOB_X0Y133_OPAD,
  output LIOB33_X0Y133_IOB_X0Y134_OPAD,
  output LIOB33_X0Y135_IOB_X0Y135_OPAD,
  output LIOB33_X0Y135_IOB_X0Y136_OPAD,
  output LIOB33_X0Y137_IOB_X0Y137_OPAD,
  output LIOB33_X0Y137_IOB_X0Y138_OPAD,
  output LIOB33_X0Y139_IOB_X0Y139_OPAD,
  output LIOB33_X0Y139_IOB_X0Y140_OPAD,
  output LIOB33_X0Y141_IOB_X0Y141_OPAD,
  output LIOB33_X0Y141_IOB_X0Y142_OPAD,
  output LIOB33_X0Y143_IOB_X0Y143_OPAD,
  output LIOB33_X0Y145_IOB_X0Y145_OPAD,
  output LIOB33_X0Y145_IOB_X0Y146_OPAD,
  output LIOB33_X0Y147_IOB_X0Y147_OPAD,
  output LIOB33_X0Y147_IOB_X0Y148_OPAD
  );
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A1;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A2;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A3;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A4;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_AMUX;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_AO5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_AO6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A_CY;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A_XOR;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B1;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B2;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B3;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B4;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_BO5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_BO6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B_CY;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B_XOR;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C1;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C2;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C3;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C4;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_CO5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_CO6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C_CY;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C_XOR;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D1;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D2;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D3;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D4;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_DO5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_DO6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D_CY;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D_XOR;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A1;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A2;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A3;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A4;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_AO5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_AO6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A_CY;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A_XOR;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B1;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B2;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B3;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B4;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_BO5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_BO6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B_CY;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B_XOR;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C1;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C2;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C3;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C4;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_CMUX;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_CO5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_CO6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C_CY;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C_XOR;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D1;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D2;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D3;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D4;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_DO5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_DO6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D_CY;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_AO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_AO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_BO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_BO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_CO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_CO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_DO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_DO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_AO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_AO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_BO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_BO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_CO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_CO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_DO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_DO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_AO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_AO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_BO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_BO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_CO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_CO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_DO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_DO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_AO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_AO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_BO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_BO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_CO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_CO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_DO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_DO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_AMUX;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_AO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_BO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_CO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_DO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_DO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_AO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_BO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_CO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_CO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_DO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_DO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_AO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_BO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_BO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_CO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_CO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_DO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_DO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_AO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_AO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_BO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_BO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_CO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_CO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_DO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_AMUX;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_AO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_A_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_BO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_B_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_CMUX;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_CO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_CO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_C_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_DO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_DO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X0Y111_D_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_AMUX;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_AO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_A_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_BMUX;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_BO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_B_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_CO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_CO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_C_XOR;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D1;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D2;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D3;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D4;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_DO5;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D_CY;
  wire [0:0] CLBLL_L_X2Y111_SLICE_X1Y111_D_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_AMUX;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_A_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_BMUX;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_BO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_BO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_B_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_CMUX;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_CO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_CO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_C_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_DO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X0Y112_D_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_AMUX;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_AO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_AO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_A_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_BO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_BO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_B_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_CO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_CO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_C_XOR;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D1;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D2;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D3;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D4;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_DO5;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_DO6;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D_CY;
  wire [0:0] CLBLL_L_X2Y112_SLICE_X1Y112_D_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_AMUX;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_AO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_A_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_BO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_BO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_B_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_CO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_CO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_C_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_DO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_DO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X0Y113_D_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_AO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_A_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_BO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_BO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_B_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_CO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_CO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_C_XOR;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D1;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D2;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D3;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D4;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_DO5;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_DO6;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D_CY;
  wire [0:0] CLBLL_L_X2Y113_SLICE_X1Y113_D_XOR;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_A;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_A1;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_A2;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_A3;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_A4;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_A5;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_A6;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_AMUX;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_AO5;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_AO6;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_A_CY;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_A_XOR;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_B;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_B1;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_B2;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_B3;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_B4;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_B5;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_B6;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_BO5;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_BO6;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_B_CY;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_B_XOR;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_C;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_C1;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_C2;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_C3;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_C4;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_C5;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_C6;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_CO5;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_CO6;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_C_CY;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_C_XOR;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_D;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_D1;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_D2;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_D3;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_D4;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_D5;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_D6;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_DO5;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_DO6;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_D_CY;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X4Y101_D_XOR;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_A;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_A1;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_A2;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_A3;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_A4;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_A5;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_A6;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_AO5;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_AO6;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_A_CY;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_A_XOR;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_B;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_B1;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_B2;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_B3;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_B4;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_B5;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_B6;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_BO5;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_BO6;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_B_CY;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_B_XOR;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_C;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_C1;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_C2;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_C3;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_C4;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_C5;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_C6;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_CO5;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_CO6;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_C_CY;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_C_XOR;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_D;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_D1;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_D2;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_D3;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_D4;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_D5;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_D6;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_DO5;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_DO6;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_D_CY;
  wire [0:0] CLBLL_L_X4Y101_SLICE_X5Y101_D_XOR;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_A;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_A1;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_A2;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_A3;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_A4;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_A5;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_A6;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_AMUX;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_AO5;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_AO6;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_A_CY;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_A_XOR;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_B;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_B1;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_B2;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_B3;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_B4;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_B5;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_B6;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_BO5;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_BO6;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_B_CY;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_B_XOR;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_C;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_C1;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_C2;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_C3;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_C4;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_C5;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_C6;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_CO5;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_CO6;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_C_CY;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_C_XOR;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_D;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_D1;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_D2;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_D3;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_D4;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_D5;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_D6;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_DO5;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_DO6;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_D_CY;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X4Y102_D_XOR;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_A;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_A1;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_A2;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_A3;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_A4;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_A5;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_A6;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_AO5;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_AO6;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_A_CY;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_A_XOR;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_B;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_B1;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_B2;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_B3;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_B4;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_B5;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_B6;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_BO5;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_BO6;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_B_CY;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_B_XOR;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_C;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_C1;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_C2;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_C3;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_C4;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_C5;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_C6;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_CO5;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_CO6;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_C_CY;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_C_XOR;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_D;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_D1;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_D2;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_D3;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_D4;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_D5;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_D6;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_DO5;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_DO6;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_D_CY;
  wire [0:0] CLBLL_L_X4Y102_SLICE_X5Y102_D_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_AMUX;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_AO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_AO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_BMUX;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_BO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_BO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_CO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_CO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_DO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_DO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_AMUX;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_AO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_AO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_BMUX;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_BO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_BO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_CO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_CO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_DO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_DO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_AMUX;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_AO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_AO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_BMUX;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_BO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_BO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_CMUX;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_CO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_DMUX;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_DO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_DO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_AMUX;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_AO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_AO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_BO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_BO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_CO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_CO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_DO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_DO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_AO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_AO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_BO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_BO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_CO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_DO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_DO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_AMUX;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_AO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_AO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_BMUX;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_BO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_CO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_CO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_DO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_DO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_AMUX;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_AO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_AO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_BMUX;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_BO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_BO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_CO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_DO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_DO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_AMUX;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_AO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_AO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_BO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_BO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_CO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_CO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_DO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_DO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_AMUX;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_AO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_BMUX;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_BO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_CO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_DO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_DO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_AMUX;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_AO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_AO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_BO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_CO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_DO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AMUX;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_BO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_CMUX;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_CO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_DO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_AO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_BO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_CO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_DO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_DO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_DMUX;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_DO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_BO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_DO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AMUX;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_A_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_BMUX;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_BO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_B_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_C_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_DO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X4Y111_D_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AMUX;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_A_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_BO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_B_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_CO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_C_XOR;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D1;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D2;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D3;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D4;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_DO5;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D_CY;
  wire [0:0] CLBLL_L_X4Y111_SLICE_X5Y111_D_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AMUX;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_A_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_BMUX;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_BO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_B_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_C_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_DO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X4Y112_D_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AMUX;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_A_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_BMUX;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_BO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_B_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_C_XOR;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D1;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D2;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D3;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D4;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_DO5;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D_CY;
  wire [0:0] CLBLL_L_X4Y112_SLICE_X5Y112_D_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_A_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_B_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_C_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_DO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X4Y113_D_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_A_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_B_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_C_XOR;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D1;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D2;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D3;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D4;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DO5;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D_CY;
  wire [0:0] CLBLL_L_X4Y113_SLICE_X5Y113_D_XOR;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_A;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_A1;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_A2;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_A3;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_A4;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_A5;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_A6;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_AO5;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_AO6;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_A_CY;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_A_XOR;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_B;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_B1;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_B2;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_B3;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_B4;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_B5;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_B6;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_BO5;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_BO6;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_B_CY;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_B_XOR;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_C;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_C1;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_C2;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_C3;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_C4;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_C5;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_C6;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_CO5;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_CO6;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_C_CY;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_C_XOR;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_D;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_D1;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_D2;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_D3;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_D4;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_D5;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_D6;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_DO5;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_DO6;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_D_CY;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X12Y101_D_XOR;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_A;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_A1;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_A2;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_A3;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_A4;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_A5;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_A6;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_AO5;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_AO6;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_A_CY;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_A_XOR;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_B;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_B1;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_B2;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_B3;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_B4;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_B5;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_B6;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_BO5;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_BO6;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_B_CY;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_B_XOR;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_C;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_C1;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_C2;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_C3;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_C4;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_C5;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_C6;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_CO5;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_CO6;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_C_CY;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_C_XOR;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_D;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_D1;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_D2;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_D3;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_D4;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_D5;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_D6;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_DO5;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_DO6;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_D_CY;
  wire [0:0] CLBLM_L_X10Y101_SLICE_X13Y101_D_XOR;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A1;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A2;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A3;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A4;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_AO5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_AO6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A_CY;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_A_XOR;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B1;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B2;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B3;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B4;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_BO5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_BO6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B_CY;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_B_XOR;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C1;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C2;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C3;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C4;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_CO5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_CO6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C_CY;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_C_XOR;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D1;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D2;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D3;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D4;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_DO5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_DO6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D_CY;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X12Y102_D_XOR;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A1;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A2;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A3;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A4;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_AMUX;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_AO5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_AO6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A_CY;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_A_XOR;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B1;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B2;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B3;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B4;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_BMUX;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_BO5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_BO6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B_CY;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_B_XOR;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C1;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C2;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C3;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C4;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_CMUX;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_CO5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_CO6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C_CY;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_C_XOR;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D1;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D2;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D3;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D4;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_DO5;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_DO6;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D_CY;
  wire [0:0] CLBLM_L_X10Y102_SLICE_X13Y102_D_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_AO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_AO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_A_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_BO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_BO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_B_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_CO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_CO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_C_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_DO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_DO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X12Y103_D_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_AMUX;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_AO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_AO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_A_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_BO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_BO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_B_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_CO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_CO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_C_XOR;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D1;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D2;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D3;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D4;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_DO5;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_DO6;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D_CY;
  wire [0:0] CLBLM_L_X10Y103_SLICE_X13Y103_D_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_AO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_AO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_A_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_BO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_B_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_CO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_CO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_C_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_DO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_DO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X12Y104_D_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_AO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_AO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_A_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_BMUX;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_BO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_BO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_B_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_CO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_CO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_C_XOR;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D1;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D2;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D3;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D4;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_DO5;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_DO6;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D_CY;
  wire [0:0] CLBLM_L_X10Y104_SLICE_X13Y104_D_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_AMUX;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_AO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_AO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_A_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_BMUX;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_BO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_BO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_B_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_CO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_CO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_C_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_DO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_DO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X12Y105_D_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_AMUX;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_AO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_AO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_A_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_BO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_BO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_B_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_CO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_CO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_C_XOR;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D1;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D2;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D3;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D4;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_DO5;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_DO6;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D_CY;
  wire [0:0] CLBLM_L_X10Y105_SLICE_X13Y105_D_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_AMUX;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_AO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_AO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_A_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_BO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_B_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_CMUX;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_CO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_CO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_C_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_DMUX;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_DO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_DO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X12Y106_D_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_AO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_A_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_BO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_BO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_B_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_CO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_C_XOR;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D1;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D2;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D3;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D4;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_DO5;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_DO6;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D_CY;
  wire [0:0] CLBLM_L_X10Y106_SLICE_X13Y106_D_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_AMUX;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_AO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_AO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_A_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_BO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_B_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_CO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_CO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_C_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_DO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_DO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X12Y107_D_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_AMUX;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_AO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_A_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_BO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_B_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_CO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_C_XOR;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D1;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D2;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D3;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D4;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_DO5;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D_CY;
  wire [0:0] CLBLM_L_X10Y107_SLICE_X13Y107_D_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_AO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_A_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_BO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_B_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_CO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_C_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_DO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X12Y108_D_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_AO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_A_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_BO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_B_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_CO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_C_XOR;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D1;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D2;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D3;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D4;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_DO5;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D_CY;
  wire [0:0] CLBLM_L_X10Y108_SLICE_X13Y108_D_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_AMUX;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_AO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_A_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_BO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_B_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_CO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_C_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_DO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X12Y109_D_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_AMUX;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_AO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_AO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_A_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_BMUX;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_BO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_B_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_CO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_C_XOR;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D1;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D2;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D3;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D4;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_DO5;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D_CY;
  wire [0:0] CLBLM_L_X10Y109_SLICE_X13Y109_D_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_AO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_AO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_A_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_BO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_BO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_B_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_CO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_C_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_DMUX;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_DO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_DO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X12Y110_D_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_AMUX;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_AO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_AO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_A_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_BMUX;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_BO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_B_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_CO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_CO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_C_XOR;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D1;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D2;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D3;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D4;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_DO5;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D_CY;
  wire [0:0] CLBLM_L_X10Y110_SLICE_X13Y110_D_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_AMUX;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_AO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_AO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_A_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_BO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_BO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_B_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_CO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_CO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_C_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_DO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X12Y111_D_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_AO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_AO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_A_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_BO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_B_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_CO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_C_XOR;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D1;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D2;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D3;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D4;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_DO5;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_DO6;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D_CY;
  wire [0:0] CLBLM_L_X10Y111_SLICE_X13Y111_D_XOR;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_A;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_A1;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_A2;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_A3;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_A4;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_A5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_A6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_AO5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_AO6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_A_CY;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_A_XOR;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_B;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_B1;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_B2;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_B3;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_B4;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_B5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_B6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_BO5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_BO6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_B_CY;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_B_XOR;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_C;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_C1;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_C2;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_C3;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_C4;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_C5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_C6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_CO5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_CO6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_C_CY;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_C_XOR;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_D;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_D1;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_D2;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_D3;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_D4;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_D5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_D6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_DO5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_DO6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_D_CY;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X16Y104_D_XOR;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_A;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_A1;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_A2;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_A3;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_A4;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_A5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_A6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_AO5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_AO6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_A_CY;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_A_XOR;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_B;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_B1;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_B2;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_B3;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_B4;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_B5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_B6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_BO5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_BO6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_B_CY;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_B_XOR;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_C;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_C1;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_C2;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_C3;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_C4;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_C5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_C6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_CO5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_CO6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_C_CY;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_C_XOR;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_D;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_D1;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_D2;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_D3;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_D4;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_D5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_D6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_DO5;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_DO6;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_D_CY;
  wire [0:0] CLBLM_L_X12Y104_SLICE_X17Y104_D_XOR;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_A;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_A1;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_A2;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_A3;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_A4;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_A5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_A6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_AO5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_AO6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_A_CY;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_A_XOR;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_B;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_B1;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_B2;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_B3;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_B4;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_B5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_B6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_BO5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_BO6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_B_CY;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_B_XOR;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_C;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_C1;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_C2;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_C3;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_C4;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_C5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_C6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_CO5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_CO6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_C_CY;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_C_XOR;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_D;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_D1;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_D2;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_D3;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_D4;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_D5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_D6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_DO5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_DO6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_D_CY;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X10Y101_D_XOR;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_A;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_A1;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_A2;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_A3;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_A4;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_A5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_A6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_AO5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_AO6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_A_CY;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_A_XOR;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_B;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_B1;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_B2;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_B3;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_B4;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_B5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_B6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_BO5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_BO6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_B_CY;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_B_XOR;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_C;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_C1;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_C2;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_C3;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_C4;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_C5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_C6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_CO5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_CO6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_C_CY;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_C_XOR;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_D;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_D1;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_D2;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_D3;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_D4;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_D5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_D6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_DO5;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_DO6;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_D_CY;
  wire [0:0] CLBLM_L_X8Y101_SLICE_X11Y101_D_XOR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A1;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A2;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A3;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A4;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_AMUX;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_AO5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_AO6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A_CY;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_A_XOR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B1;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B2;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B3;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B4;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_BO5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_BO6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B_CY;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_B_XOR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C1;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C2;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C3;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C4;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_CO5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_CO6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C_CY;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_C_XOR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D1;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D2;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D3;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D4;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_DO5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_DO6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D_CY;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X10Y102_D_XOR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A1;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A2;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A3;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A4;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_AMUX;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_AO5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_AO6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A_CY;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_A_XOR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B1;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B2;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B3;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B4;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_BO5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_BO6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B_CY;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_B_XOR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C1;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C2;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C3;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C4;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_CO5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_CO6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C_CY;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_C_XOR;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D1;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D2;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D3;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D4;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_DO5;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_DO6;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D_CY;
  wire [0:0] CLBLM_L_X8Y102_SLICE_X11Y102_D_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_AO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_AO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_A_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_BO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_BO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_B_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_CO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_CO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_C_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_DO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_DO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X10Y103_D_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_AO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_AO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_A_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_BO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_BO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_B_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_CO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_CO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_C_XOR;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D1;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D2;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D3;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D4;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_DO5;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_DO6;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D_CY;
  wire [0:0] CLBLM_L_X8Y103_SLICE_X11Y103_D_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_AO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_A_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_BO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_BO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_B_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_CO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_CO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_C_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_DO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_DO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X10Y104_D_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_AO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_AO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_A_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_BO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_BO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_B_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_CO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_CO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_C_XOR;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D1;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D2;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D3;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D4;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_DO5;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_DO6;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D_CY;
  wire [0:0] CLBLM_L_X8Y104_SLICE_X11Y104_D_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_AMUX;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_AO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_AO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_A_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_BO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_BO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_B_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_CO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_CO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_C_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_DO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_DO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X10Y105_D_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_AO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_AO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_A_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_BO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_BO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_B_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_CO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_CO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_C_XOR;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D1;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D2;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D3;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D4;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_DO5;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_DO6;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D_CY;
  wire [0:0] CLBLM_L_X8Y105_SLICE_X11Y105_D_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_AO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_AO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_A_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_BO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_BO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_B_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_CO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_CO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_C_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_DO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_DO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X10Y106_D_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_AO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_A_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_BO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_BO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_B_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_CO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_CO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_C_XOR;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D1;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D2;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D3;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D4;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_DO5;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_DO6;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D_CY;
  wire [0:0] CLBLM_L_X8Y106_SLICE_X11Y106_D_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_AMUX;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_AO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_AO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_A_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_BO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_B_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_CO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_CO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_C_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_DO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_DO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X10Y107_D_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_AMUX;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_AO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_A_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_BO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_BO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_B_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_CO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_CO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_C_XOR;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D1;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D2;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D3;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D4;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_DO5;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_DO6;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D_CY;
  wire [0:0] CLBLM_L_X8Y107_SLICE_X11Y107_D_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_AO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_A_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_BO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_B_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_CO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_CO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_C_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_DO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_DO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X10Y108_D_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_AO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_A_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_BO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_BO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_B_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_CO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_CO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_C_XOR;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D1;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D2;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D3;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D4;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_DO5;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_DO6;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D_CY;
  wire [0:0] CLBLM_L_X8Y108_SLICE_X11Y108_D_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_AO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_AO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_A_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_BO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_B_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_CO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_C_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_DO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_DO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X10Y109_D_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_AMUX;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_AO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_A_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_BO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_BO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_B_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_CO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_CO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_C_XOR;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D1;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D2;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D3;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D4;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_DO5;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_DO6;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D_CY;
  wire [0:0] CLBLM_L_X8Y109_SLICE_X11Y109_D_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_AO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_A_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_BO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_B_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_CO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_C_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_DO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X10Y110_D_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_AO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_A_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_BO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_B_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_CO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_C_XOR;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D1;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D2;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D3;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D4;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_DO5;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D_CY;
  wire [0:0] CLBLM_L_X8Y110_SLICE_X11Y110_D_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_AMUX;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_AO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_A_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_BMUX;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_BO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_B_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_CMUX;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_CO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_C_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_DO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X10Y111_D_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_AO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_A_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_BO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_B_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_CO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_C_XOR;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D1;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D2;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D3;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D4;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_DO5;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_DO6;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D_CY;
  wire [0:0] CLBLM_L_X8Y111_SLICE_X11Y111_D_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_AO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_A_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_BO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_B_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_CO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_C_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_DO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X10Y112_D_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_AMUX;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_AO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_A_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_BO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_B_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_CMUX;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_CO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_C_XOR;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D1;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D2;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D3;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D4;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_DO5;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_DO6;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D_CY;
  wire [0:0] CLBLM_L_X8Y112_SLICE_X11Y112_D_XOR;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_A;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_A1;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_A2;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_A3;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_A4;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_A5;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_A6;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_AMUX;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_AO5;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_AO6;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_A_CY;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_A_XOR;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_B;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_B1;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_B2;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_B3;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_B4;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_B5;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_B6;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_BO5;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_BO6;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_B_CY;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_B_XOR;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_C;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_C1;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_C2;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_C3;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_C4;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_C5;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_C6;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_CO5;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_CO6;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_C_CY;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_C_XOR;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_D;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_D1;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_D2;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_D3;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_D4;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_D5;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_D6;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_DO5;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_DO6;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_D_CY;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X14Y103_D_XOR;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_A;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_A1;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_A2;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_A3;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_A4;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_A5;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_A6;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_AO5;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_AO6;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_A_CY;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_A_XOR;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_B;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_B1;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_B2;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_B3;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_B4;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_B5;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_B6;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_BO5;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_BO6;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_B_CY;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_B_XOR;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_C;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_C1;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_C2;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_C3;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_C4;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_C5;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_C6;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_CO5;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_CO6;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_C_CY;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_C_XOR;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_D;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_D1;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_D2;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_D3;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_D4;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_D5;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_D6;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_DO5;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_DO6;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_D_CY;
  wire [0:0] CLBLM_R_X11Y103_SLICE_X15Y103_D_XOR;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A1;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A2;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A3;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A4;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_AMUX;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_AO5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_AO6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A_CY;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_A_XOR;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B1;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B2;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B3;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B4;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_BO5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_BO6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B_CY;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_B_XOR;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C1;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C2;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C3;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C4;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_CO5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_CO6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C_CY;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_C_XOR;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D1;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D2;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D3;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D4;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_DO5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_DO6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D_CY;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X14Y104_D_XOR;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A1;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A2;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A3;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A4;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_AMUX;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_AO5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_AO6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A_CY;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_A_XOR;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B1;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B2;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B3;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B4;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_BMUX;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_BO5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_BO6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B_CY;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_B_XOR;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C1;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C2;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C3;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C4;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_CO5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_CO6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C_CY;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_C_XOR;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D1;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D2;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D3;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D4;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_DO5;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_DO6;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D_CY;
  wire [0:0] CLBLM_R_X11Y104_SLICE_X15Y104_D_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_AMUX;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_AO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_AO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_A_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_BO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_BO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_B_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_CO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_CO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_C_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_DO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_DO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X14Y105_D_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_AO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_AO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_A_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_BO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_BO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_B_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_CMUX;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_CO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_CO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_C_XOR;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D1;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D2;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D3;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D4;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_DO5;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_DO6;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D_CY;
  wire [0:0] CLBLM_R_X11Y105_SLICE_X15Y105_D_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_AO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_A_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_BO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_B_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_CO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_C_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_DO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_DO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X14Y106_D_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_AMUX;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_AO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_AO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_A_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_BMUX;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_BO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_B_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_CO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_CO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_C_XOR;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D1;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D2;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D3;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D4;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_DO5;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_DO6;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D_CY;
  wire [0:0] CLBLM_R_X11Y106_SLICE_X15Y106_D_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_AMUX;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_AO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_AO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_A_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_BO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_BO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_B_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_CO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_CO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_C_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_DO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_DO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X14Y107_D_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_AMUX;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_AO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_AO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_A_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_BO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_BO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_B_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_CMUX;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_CO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_CO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_C_XOR;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D1;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D2;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D3;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D4;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_DO5;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_DO6;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D_CY;
  wire [0:0] CLBLM_R_X11Y107_SLICE_X15Y107_D_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_AO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_AO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_A_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_BO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_B_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_CO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_CO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_C_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_DO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_DO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X14Y108_D_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_AMUX;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_AO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_AO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_A_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_BO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_BO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_B_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_CMUX;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_CO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_C_XOR;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D1;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D2;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D3;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D4;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_DO5;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_DO6;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D_CY;
  wire [0:0] CLBLM_R_X11Y108_SLICE_X15Y108_D_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_AMUX;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_AO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_AO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_A_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_BO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_B_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_CO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_CO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_C_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_DO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_DO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X14Y109_D_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_AO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_A_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_BO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_BO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_B_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_CO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_CO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_C_XOR;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D1;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D2;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D3;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D4;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_DO5;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_DO6;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D_CY;
  wire [0:0] CLBLM_R_X11Y109_SLICE_X15Y109_D_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_AMUX;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_AO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_AO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_A_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_BO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_BO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_B_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_CO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_CO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_C_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_DO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_DO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X14Y110_D_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_AO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_AO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_A_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_BO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_BO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_B_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_CO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_CO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_C_XOR;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D1;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D2;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D3;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D4;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_DO5;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_DO6;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D_CY;
  wire [0:0] CLBLM_R_X11Y110_SLICE_X15Y110_D_XOR;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_A;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_A1;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_A2;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_A3;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_A4;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_A5;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_A6;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_AMUX;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_AO5;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_AO6;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_A_CY;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_A_XOR;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_B;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_B1;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_B2;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_B3;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_B4;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_B5;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_B6;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_BMUX;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_BO5;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_BO6;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_B_CY;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_B_XOR;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_C;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_C1;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_C2;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_C3;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_C4;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_C5;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_C6;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_CO5;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_CO6;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_C_CY;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_C_XOR;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_D;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_D1;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_D2;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_D3;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_D4;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_D5;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_D6;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_DO5;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_DO6;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_D_CY;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X2Y102_D_XOR;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_A;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_A1;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_A2;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_A3;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_A4;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_A5;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_A6;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_AMUX;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_AO5;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_AO6;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_A_CY;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_A_XOR;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_B;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_B1;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_B2;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_B3;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_B4;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_B5;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_B6;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_BO5;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_BO6;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_B_CY;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_B_XOR;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_C;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_C1;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_C2;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_C3;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_C4;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_C5;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_C6;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_CO5;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_CO6;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_C_CY;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_C_XOR;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_D;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_D1;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_D2;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_D3;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_D4;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_D5;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_D6;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_DO5;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_DO6;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_D_CY;
  wire [0:0] CLBLM_R_X3Y102_SLICE_X3Y102_D_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_AO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_AO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_BO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_BO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_CO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_CO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_DO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_DO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_AMUX;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_AO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_AO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_BO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_BO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_CMUX;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_CO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_CO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_DO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_DO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_AMUX;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_AO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_AO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_BO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_BO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_CO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_CO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_DO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_DO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_AMUX;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_AO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_AO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_BMUX;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_BO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_CO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_CO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_DO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_DO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_AO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_BO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_BO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_CO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_CO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_DO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_DO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_AMUX;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_AO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_AO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_BMUX;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_BO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_CMUX;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_CO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_DO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_DO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_AO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_AO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_BO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_BO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_CO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_DO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_DO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_AMUX;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_AO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_AO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_BO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_CO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_CO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_DO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_DO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_AMUX;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_AO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_BO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_BO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_CMUX;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_CO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_DO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_DO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_AO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_AO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_BO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_BO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_CO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_DMUX;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_DO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_DO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_AO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_AO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_BO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_BO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_CO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_CO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_DO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_AO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_BO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_CO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_DO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AMUX;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_BMUX;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_BO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_BO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_DO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_DO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AMUX;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_BO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_DO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AMUX;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_BO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_CO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_DO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AMUX;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_BO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_CO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_DO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_AMUX;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_A_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_BO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_B_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_CO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_C_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_DO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_DO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X2Y111_D_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AMUX;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_A_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_BMUX;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_BO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_B_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_CMUX;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_CO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_C_XOR;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D1;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D2;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D3;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D4;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_DO5;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D_CY;
  wire [0:0] CLBLM_R_X3Y111_SLICE_X3Y111_D_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_A_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_BO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_B_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_CO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_C_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_DO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X2Y112_D_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AMUX;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_A_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_B_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_C_XOR;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D1;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D2;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D3;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D4;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_DO5;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D_CY;
  wire [0:0] CLBLM_R_X3Y112_SLICE_X3Y112_D_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AMUX;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_A_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_BMUX;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_BO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_BO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_B_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_CMUX;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_CO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_C_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_DO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X2Y113_D_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_A_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_BMUX;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_BO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_B_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_CO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_C_XOR;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D1;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D2;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D3;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D4;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_DO5;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D_CY;
  wire [0:0] CLBLM_R_X3Y113_SLICE_X3Y113_D_XOR;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_A;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_A1;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_A2;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_A3;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_A4;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_A5;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_A6;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_AO5;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_AO6;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_A_CY;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_A_XOR;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_B;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_B1;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_B2;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_B3;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_B4;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_B5;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_B6;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_BO5;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_BO6;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_B_CY;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_B_XOR;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_C;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_C1;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_C2;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_C3;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_C4;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_C5;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_C6;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_CO5;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_CO6;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_C_CY;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_C_XOR;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_D;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_D1;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_D2;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_D3;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_D4;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_D5;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_D6;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_DO5;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_DO6;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_D_CY;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X6Y100_D_XOR;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_A;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_A1;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_A2;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_A3;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_A4;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_A5;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_A6;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_AO5;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_AO6;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_A_CY;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_A_XOR;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_B;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_B1;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_B2;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_B3;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_B4;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_B5;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_B6;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_BO5;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_BO6;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_B_CY;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_B_XOR;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_C;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_C1;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_C2;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_C3;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_C4;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_C5;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_C6;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_CO5;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_CO6;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_C_CY;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_C_XOR;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_D;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_D1;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_D2;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_D3;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_D4;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_D5;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_D6;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_DO5;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_DO6;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_D_CY;
  wire [0:0] CLBLM_R_X5Y100_SLICE_X7Y100_D_XOR;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_A;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_A1;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_A2;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_A3;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_A4;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_A5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_A6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_AMUX;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_AO5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_AO6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_A_CY;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_A_XOR;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_B;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_B1;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_B2;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_B3;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_B4;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_B5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_B6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_BO5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_BO6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_B_CY;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_B_XOR;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_C;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_C1;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_C2;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_C3;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_C4;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_C5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_C6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_CO5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_CO6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_C_CY;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_C_XOR;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_D;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_D1;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_D2;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_D3;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_D4;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_D5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_D6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_DO5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_DO6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_D_CY;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X6Y101_D_XOR;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_A;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_A1;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_A2;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_A3;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_A4;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_A5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_A6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_AMUX;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_AO5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_AO6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_A_CY;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_A_XOR;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_B;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_B1;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_B2;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_B3;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_B4;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_B5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_B6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_BO5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_BO6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_B_CY;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_B_XOR;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_C;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_C1;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_C2;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_C3;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_C4;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_C5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_C6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_CO5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_CO6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_C_CY;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_C_XOR;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_D;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_D1;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_D2;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_D3;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_D4;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_D5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_D6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_DO5;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_DO6;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_D_CY;
  wire [0:0] CLBLM_R_X5Y101_SLICE_X7Y101_D_XOR;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_A;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_A1;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_A2;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_A3;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_A4;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_A5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_A6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_AO5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_AO6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_A_CY;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_A_XOR;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_B;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_B1;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_B2;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_B3;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_B4;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_B5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_B6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_BO5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_BO6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_B_CY;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_B_XOR;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_C;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_C1;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_C2;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_C3;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_C4;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_C5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_C6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_CMUX;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_CO5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_CO6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_C_CY;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_C_XOR;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_D;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_D1;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_D2;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_D3;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_D4;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_D5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_D6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_DO5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_DO6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_D_CY;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X6Y102_D_XOR;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_A;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_A1;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_A2;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_A3;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_A4;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_A5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_A6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_AMUX;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_AO5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_AO6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_A_CY;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_A_XOR;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_B;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_B1;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_B2;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_B3;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_B4;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_B5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_B6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_BMUX;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_BO5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_BO6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_B_CY;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_B_XOR;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_C;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_C1;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_C2;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_C3;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_C4;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_C5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_C6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_CO5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_CO6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_C_CY;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_C_XOR;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_D;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_D1;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_D2;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_D3;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_D4;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_D5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_D6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_DO5;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_DO6;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_D_CY;
  wire [0:0] CLBLM_R_X5Y102_SLICE_X7Y102_D_XOR;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A1;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A2;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A3;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A4;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_AMUX;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_AO5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_AO6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A_CY;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A_XOR;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B1;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B2;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B3;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B4;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_BO5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_BO6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B_CY;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B_XOR;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C1;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C2;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C3;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C4;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_CO5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_CO6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C_CY;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C_XOR;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D1;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D2;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D3;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D4;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_DO5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_DO6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D_CY;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D_XOR;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A1;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A2;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A3;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A4;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_AO5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_AO6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A_CY;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A_XOR;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B1;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B2;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B3;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B4;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_BO5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_BO6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B_CY;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B_XOR;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C1;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C2;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C3;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C4;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_CO5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_CO6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C_CY;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C_XOR;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D1;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D2;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D3;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D4;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_DO5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_DO6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D_CY;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_AMUX;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_AO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_AO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_BO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_BO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_CO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_CO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_DO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_DO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_AMUX;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_AO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_AO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_BO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_BO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_CO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_CO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_DO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_DO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_AMUX;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_AO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_BO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_BO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_CO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_CO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_DO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_DO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_AMUX;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_AO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_AO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_BMUX;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_BO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_BO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_CO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_DO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_DO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_AMUX;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_AO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_BO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_CO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_DO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_AMUX;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_AO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_AO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_BMUX;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_BO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_CO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_CO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_DO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_DO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_AO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_BO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_CO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_CO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_DMUX;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_DO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_AMUX;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_AO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_AO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_BO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_CO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_CO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_DO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_DO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_AO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_A_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_BO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_B_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_CO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_C_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_DO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X6Y108_D_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_AO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_AO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_A_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_BO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_B_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_CMUX;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_CO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_C_XOR;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D1;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D2;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D3;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D4;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_DO5;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_DO6;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D_CY;
  wire [0:0] CLBLM_R_X5Y108_SLICE_X7Y108_D_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_AMUX;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_AO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_A_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_BO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_B_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_CO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_C_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_DO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X6Y109_D_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AMUX;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_A_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_BO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_B_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_CO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_C_XOR;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D1;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D2;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D3;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D4;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_DO5;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_DO6;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D_CY;
  wire [0:0] CLBLM_R_X5Y109_SLICE_X7Y109_D_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_AO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_A_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_BO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_B_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_CO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_C_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_DO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X6Y110_D_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_AMUX;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_AO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_A_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_BO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_B_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_CO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_C_XOR;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D1;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D2;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D3;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D4;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_DO5;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D_CY;
  wire [0:0] CLBLM_R_X5Y110_SLICE_X7Y110_D_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_AMUX;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_AO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_A_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_BO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_B_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_CO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_C_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_DO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X6Y111_D_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_AMUX;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_AO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_A_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_BMUX;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_BO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_B_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_CO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_C_XOR;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D1;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D2;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D3;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D4;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_DO5;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D_CY;
  wire [0:0] CLBLM_R_X5Y111_SLICE_X7Y111_D_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AMUX;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_A_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_BO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_B_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_CO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_C_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_DO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X6Y112_D_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_A_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_BO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_BO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_B_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_CO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_CO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_C_XOR;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D1;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D2;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D3;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D4;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_DO5;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D_CY;
  wire [0:0] CLBLM_R_X5Y112_SLICE_X7Y112_D_XOR;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_A;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_A1;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_A2;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_A3;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_A4;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_A5;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_A6;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_AMUX;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_AO5;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_AO6;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_A_CY;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_A_XOR;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_B;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_B1;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_B2;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_B3;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_B4;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_B5;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_B6;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_BMUX;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_BO5;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_BO6;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_B_CY;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_B_XOR;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_C;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_C1;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_C2;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_C3;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_C4;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_C5;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_C6;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_CO5;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_CO6;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_C_CY;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_C_XOR;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_D;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_D1;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_D2;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_D3;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_D4;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_D5;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_D6;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_DO5;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_DO6;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_D_CY;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X8Y100_D_XOR;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_A;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_A1;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_A2;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_A3;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_A4;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_A5;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_A6;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_AO5;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_AO6;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_A_CY;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_A_XOR;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_B;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_B1;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_B2;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_B3;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_B4;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_B5;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_B6;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_BO5;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_BO6;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_B_CY;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_B_XOR;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_C;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_C1;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_C2;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_C3;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_C4;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_C5;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_C6;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_CO5;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_CO6;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_C_CY;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_C_XOR;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_D;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_D1;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_D2;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_D3;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_D4;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_D5;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_D6;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_DO5;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_DO6;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_D_CY;
  wire [0:0] CLBLM_R_X7Y100_SLICE_X9Y100_D_XOR;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_A;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_A1;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_A2;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_A3;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_A4;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_A5;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_A6;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_AMUX;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_AO5;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_AO6;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_A_CY;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_A_XOR;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_B;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_B1;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_B2;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_B3;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_B4;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_B5;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_B6;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_BMUX;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_BO5;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_BO6;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_B_CY;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_B_XOR;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_C;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_C1;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_C2;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_C3;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_C4;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_C5;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_C6;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_CMUX;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_CO5;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_CO6;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_C_CY;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_C_XOR;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_D;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_D1;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_D2;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_D3;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_D4;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_D5;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_D6;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_DO5;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_DO6;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_D_CY;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X8Y101_D_XOR;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_A;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_A1;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_A2;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_A3;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_A4;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_A5;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_A6;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_AO5;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_AO6;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_A_CY;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_A_XOR;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_B;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_B1;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_B2;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_B3;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_B4;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_B5;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_B6;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_BO5;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_BO6;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_B_CY;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_B_XOR;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_C;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_C1;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_C2;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_C3;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_C4;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_C5;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_C6;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_CO5;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_CO6;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_C_CY;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_C_XOR;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_D;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_D1;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_D2;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_D3;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_D4;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_D5;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_D6;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_DO5;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_DO6;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_D_CY;
  wire [0:0] CLBLM_R_X7Y101_SLICE_X9Y101_D_XOR;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A1;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A2;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A3;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A4;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_AMUX;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_AO5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_AO6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A_CY;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_A_XOR;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B1;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B2;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B3;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B4;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_BO5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_BO6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B_CY;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_B_XOR;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C1;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C2;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C3;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C4;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_CO5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_CO6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C_CY;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_C_XOR;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D1;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D2;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D3;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D4;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_DO5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_DO6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D_CY;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X8Y102_D_XOR;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A1;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A2;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A3;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A4;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_AO5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_AO6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A_CY;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_A_XOR;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B1;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B2;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B3;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B4;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_BO5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_BO6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B_CY;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_B_XOR;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C1;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C2;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C3;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C4;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_CO5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_CO6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C_CY;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_C_XOR;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D1;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D2;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D3;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D4;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_DO5;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_DO6;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D_CY;
  wire [0:0] CLBLM_R_X7Y102_SLICE_X9Y102_D_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_AMUX;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_AO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_AO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_A_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_BO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_BO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_B_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_CO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_CO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_C_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_DO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_DO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X8Y103_D_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_AMUX;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_AO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_AO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_A_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_BO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_BO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_B_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_CMUX;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_CO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_CO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_C_XOR;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D1;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D2;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D3;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D4;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_DO5;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_DO6;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D_CY;
  wire [0:0] CLBLM_R_X7Y103_SLICE_X9Y103_D_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_AMUX;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_AO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_AO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_A_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_BMUX;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_BO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_BO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_B_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_CO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_CO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_C_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_DMUX;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_DO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_DO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X8Y104_D_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_AMUX;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_AO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_AO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_A_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_BO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_BO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_B_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_CO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_CO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_C_XOR;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D1;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D2;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D3;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D4;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_DO5;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_DO6;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D_CY;
  wire [0:0] CLBLM_R_X7Y104_SLICE_X9Y104_D_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_AO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_AO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_A_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_BO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_BO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_B_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_CO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_CO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_C_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_DO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_DO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X8Y105_D_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_AO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_AO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_A_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_BO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_BO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_B_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_CO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_CO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_C_XOR;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D1;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D2;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D3;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D4;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_DO5;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_DO6;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D_CY;
  wire [0:0] CLBLM_R_X7Y105_SLICE_X9Y105_D_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_AO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_A_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_BO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_BO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_B_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_CO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_C_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_DO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_DO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X8Y106_D_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_AMUX;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_AO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_AO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_A_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_BO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_BO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_B_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_CO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_CO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_C_XOR;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D1;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D2;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D3;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D4;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_DO5;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_DO6;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D_CY;
  wire [0:0] CLBLM_R_X7Y106_SLICE_X9Y106_D_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_AO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_A_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_BO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_BO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_B_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_CO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_CO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_C_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_DO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_DO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X8Y107_D_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_AMUX;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_AO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_AO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_A_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_BMUX;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_BO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_B_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_CMUX;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_CO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_CO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_C_XOR;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D1;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D2;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D3;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D4;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_DO5;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_DO6;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D_CY;
  wire [0:0] CLBLM_R_X7Y107_SLICE_X9Y107_D_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_AO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_A_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_BO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_B_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_CO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_CO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_C_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_DO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_DO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X8Y108_D_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_AMUX;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_AO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_A_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_BMUX;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_BO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_B_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_CO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_C_XOR;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D1;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D2;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D3;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D4;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_DO5;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_DO6;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D_CY;
  wire [0:0] CLBLM_R_X7Y108_SLICE_X9Y108_D_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_AO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_A_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_BO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_B_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_CO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_C_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_DO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X8Y109_D_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_AMUX;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_AO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_A_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_BO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_BO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_B_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_CO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_C_XOR;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D1;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D2;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D3;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D4;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_DO5;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D_CY;
  wire [0:0] CLBLM_R_X7Y109_SLICE_X9Y109_D_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_AMUX;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_AO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_AO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_A_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_BO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_B_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_CO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_C_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_DO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X8Y110_D_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_AMUX;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_A_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_BO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_B_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_CO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_C_XOR;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D1;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D2;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D3;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D4;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_DO5;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D_CY;
  wire [0:0] CLBLM_R_X7Y110_SLICE_X9Y110_D_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_AMUX;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_AO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_A_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_BO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_B_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_CO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_C_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_DO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X8Y111_D_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_AO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_A_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_BO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_B_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_CO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_C_XOR;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D1;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D2;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D3;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D4;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_DO5;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_DO6;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D_CY;
  wire [0:0] CLBLM_R_X7Y111_SLICE_X9Y111_D_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_AO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_A_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_BO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_B_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_CO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_C_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_DO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X8Y112_D_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_AMUX;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_A_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_BO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_B_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_CO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_C_XOR;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D1;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D2;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D3;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D4;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_DO5;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D_CY;
  wire [0:0] CLBLM_R_X7Y112_SLICE_X9Y112_D_XOR;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_I;
  wire [0:0] LIOB33_SING_X0Y149_IOB_X0Y149_O;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y125_O;
  wire [0:0] LIOB33_X0Y125_IOB_X0Y126_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y127_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y129_O;
  wire [0:0] LIOB33_X0Y129_IOB_X0Y130_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y131_O;
  wire [0:0] LIOB33_X0Y131_IOB_X0Y132_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y133_O;
  wire [0:0] LIOB33_X0Y133_IOB_X0Y134_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y135_O;
  wire [0:0] LIOB33_X0Y135_IOB_X0Y136_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y137_O;
  wire [0:0] LIOB33_X0Y137_IOB_X0Y138_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y139_O;
  wire [0:0] LIOB33_X0Y139_IOB_X0Y140_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y141_O;
  wire [0:0] LIOB33_X0Y141_IOB_X0Y142_O;
  wire [0:0] LIOB33_X0Y143_IOB_X0Y143_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y145_O;
  wire [0:0] LIOB33_X0Y145_IOB_X0Y146_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y147_O;
  wire [0:0] LIOB33_X0Y147_IOB_X0Y148_O;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_D;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_O;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1;
  wire [0:0] LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_O;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_O;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_D1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_OQ;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_T1;
  wire [0:0] LIOI3_X0Y117_OLOGIC_X0Y118_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y125_TQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_D1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_OQ;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_T1;
  wire [0:0] LIOI3_X0Y125_OLOGIC_X0Y126_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y127_TQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_D1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_OQ;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_T1;
  wire [0:0] LIOI3_X0Y127_OLOGIC_X0Y128_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y129_TQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_D1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_OQ;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_T1;
  wire [0:0] LIOI3_X0Y129_OLOGIC_X0Y130_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y133_TQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_D1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_OQ;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_T1;
  wire [0:0] LIOI3_X0Y133_OLOGIC_X0Y134_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y135_TQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_D1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_OQ;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_T1;
  wire [0:0] LIOI3_X0Y135_OLOGIC_X0Y136_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y139_TQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_D1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_OQ;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_T1;
  wire [0:0] LIOI3_X0Y139_OLOGIC_X0Y140_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y141_TQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_D1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_OQ;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_T1;
  wire [0:0] LIOI3_X0Y141_OLOGIC_X0Y142_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y145_TQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_D1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_OQ;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_T1;
  wire [0:0] LIOI3_X0Y145_OLOGIC_X0Y146_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y147_TQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_D1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_OQ;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_T1;
  wire [0:0] LIOI3_X0Y147_OLOGIC_X0Y148_TQ;
  wire [0:0] RIOB33_SING_X105Y100_IOB_X1Y100_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y101_I;
  wire [0:0] RIOB33_X105Y101_IOB_X1Y102_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y103_I;
  wire [0:0] RIOB33_X105Y103_IOB_X1Y104_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y105_I;
  wire [0:0] RIOB33_X105Y105_IOB_X1Y106_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y107_I;
  wire [0:0] RIOB33_X105Y107_IOB_X1Y108_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y109_I;
  wire [0:0] RIOB33_X105Y109_IOB_X1Y110_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y111_I;
  wire [0:0] RIOB33_X105Y111_IOB_X1Y112_I;
  wire [0:0] RIOB33_X105Y113_IOB_X1Y113_I;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_D;
  wire [0:0] RIOI3_SING_X105Y100_ILOGIC_X1Y100_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D;
  wire [0:0] RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D;
  wire [0:0] RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y101_O;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_D;
  wire [0:0] RIOI3_X105Y101_ILOGIC_X1Y102_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y103_O;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_D;
  wire [0:0] RIOI3_X105Y103_ILOGIC_X1Y104_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y105_O;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_D;
  wire [0:0] RIOI3_X105Y105_ILOGIC_X1Y106_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y109_O;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_D;
  wire [0:0] RIOI3_X105Y109_ILOGIC_X1Y110_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y111_O;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_D;
  wire [0:0] RIOI3_X105Y111_ILOGIC_X1Y112_O;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f13ff5fb320ffa0)
  ) CLBLL_L_X2Y103_SLICE_X0Y103_DLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(CLBLL_L_X2Y103_SLICE_X0Y103_AO5),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLL_L_X2Y104_SLICE_X0Y104_AO6),
.O5(CLBLL_L_X2Y103_SLICE_X0Y103_DO5),
.O6(CLBLL_L_X2Y103_SLICE_X0Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93a05f936c5fa0)
  ) CLBLL_L_X2Y103_SLICE_X0Y103_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(CLBLL_L_X2Y103_SLICE_X0Y103_AO5),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLL_L_X2Y104_SLICE_X0Y104_AO6),
.O5(CLBLL_L_X2Y103_SLICE_X0Y103_CO5),
.O6(CLBLL_L_X2Y103_SLICE_X0Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he7dd18229a009a00)
  ) CLBLL_L_X2Y103_SLICE_X0Y103_BLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(CLBLL_L_X2Y103_SLICE_X1Y103_DO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(RIOB33_X105Y109_IOB_X1Y110_I),
.O5(CLBLL_L_X2Y103_SLICE_X0Y103_BO5),
.O6(CLBLL_L_X2Y103_SLICE_X0Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3f00f30f3f0ff)
  ) CLBLL_L_X2Y103_SLICE_X0Y103_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(CLBLL_L_X2Y103_SLICE_X1Y103_AO6),
.I3(CLBLL_L_X2Y103_SLICE_X0Y103_BO6),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y103_SLICE_X0Y103_AO5),
.O6(CLBLL_L_X2Y103_SLICE_X0Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f07ff7f7f3fff7f)
  ) CLBLL_L_X2Y103_SLICE_X1Y103_DLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(RIOB33_X105Y111_IOB_X1Y111_I),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(CLBLM_R_X3Y102_SLICE_X2Y102_AO6),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLL_L_X2Y103_SLICE_X1Y103_DO5),
.O6(CLBLL_L_X2Y103_SLICE_X1Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3cb33b37f3fff7f)
  ) CLBLL_L_X2Y103_SLICE_X1Y103_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(RIOB33_X105Y111_IOB_X1Y111_I),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(CLBLM_R_X3Y102_SLICE_X2Y102_AO6),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLL_L_X2Y103_SLICE_X1Y103_CO5),
.O6(CLBLL_L_X2Y103_SLICE_X1Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ca0935f935f6ca0)
  ) CLBLL_L_X2Y103_SLICE_X1Y103_BLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(CLBLL_L_X2Y103_SLICE_X1Y103_CO6),
.I5(CLBLL_L_X4Y102_SLICE_X4Y102_BO6),
.O5(CLBLL_L_X2Y103_SLICE_X1Y103_BO5),
.O6(CLBLL_L_X2Y103_SLICE_X1Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffdf5f135f4c00)
  ) CLBLL_L_X2Y103_SLICE_X1Y103_ALUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(CLBLL_L_X2Y103_SLICE_X1Y103_CO6),
.I5(CLBLL_L_X4Y102_SLICE_X4Y102_BO6),
.O5(CLBLL_L_X2Y103_SLICE_X1Y103_AO5),
.O6(CLBLL_L_X2Y103_SLICE_X1Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y104_SLICE_X0Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y104_SLICE_X0Y104_DO5),
.O6(CLBLL_L_X2Y104_SLICE_X0Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y104_SLICE_X0Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y104_SLICE_X0Y104_CO5),
.O6(CLBLL_L_X2Y104_SLICE_X0Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y104_SLICE_X0Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y104_SLICE_X0Y104_BO5),
.O6(CLBLL_L_X2Y104_SLICE_X0Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa2f4fbf4fff0fff)
  ) CLBLL_L_X2Y104_SLICE_X0Y104_ALUT (
.I0(CLBLL_L_X2Y103_SLICE_X1Y103_DO6),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLL_L_X2Y104_SLICE_X0Y104_AO5),
.O6(CLBLL_L_X2Y104_SLICE_X0Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y104_SLICE_X1Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y104_SLICE_X1Y104_DO5),
.O6(CLBLL_L_X2Y104_SLICE_X1Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y104_SLICE_X1Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y104_SLICE_X1Y104_CO5),
.O6(CLBLL_L_X2Y104_SLICE_X1Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y104_SLICE_X1Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y104_SLICE_X1Y104_BO5),
.O6(CLBLL_L_X2Y104_SLICE_X1Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y104_SLICE_X1Y104_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y104_SLICE_X1Y104_AO5),
.O6(CLBLL_L_X2Y104_SLICE_X1Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y105_SLICE_X0Y105_DO5),
.O6(CLBLL_L_X2Y105_SLICE_X0Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y105_SLICE_X0Y105_CO5),
.O6(CLBLL_L_X2Y105_SLICE_X0Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd7dfb5975f5fdf5f)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_BLUT (
.I0(RIOB33_X105Y111_IOB_X1Y111_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(CLBLL_L_X2Y105_SLICE_X0Y105_AO6),
.I5(LIOB33_X0Y113_IOB_X0Y113_I),
.O5(CLBLL_L_X2Y105_SLICE_X0Y105_BO5),
.O6(CLBLL_L_X2Y105_SLICE_X0Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2bbf3bff2fffbfff)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_ALUT (
.I0(CLBLL_L_X2Y103_SLICE_X1Y103_DO6),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLL_L_X2Y105_SLICE_X0Y105_AO5),
.O6(CLBLL_L_X2Y105_SLICE_X0Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y105_SLICE_X1Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y105_SLICE_X1Y105_DO5),
.O6(CLBLL_L_X2Y105_SLICE_X1Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y105_SLICE_X1Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y105_SLICE_X1Y105_CO5),
.O6(CLBLL_L_X2Y105_SLICE_X1Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y105_SLICE_X1Y105_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y105_SLICE_X1Y105_BO5),
.O6(CLBLL_L_X2Y105_SLICE_X1Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y105_SLICE_X1Y105_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y105_SLICE_X1Y105_AO5),
.O6(CLBLL_L_X2Y105_SLICE_X1Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f137f1fff7fffff)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_DLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(RIOB33_X105Y111_IOB_X1Y111_I),
.I3(CLBLL_L_X2Y105_SLICE_X0Y105_AO6),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(LIOB33_X0Y113_IOB_X0Y113_I),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_DO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h08888fff0008888f)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_CLUT (
.I0(RIOB33_X105Y111_IOB_X1Y111_I),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(CLBLL_L_X2Y103_SLICE_X0Y103_DO6),
.I3(CLBLM_R_X3Y103_SLICE_X2Y103_CO6),
.I4(CLBLL_L_X2Y106_SLICE_X0Y106_DO6),
.I5(CLBLL_L_X2Y106_SLICE_X0Y106_BO6),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_CO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha6aacc00996a0cc0)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(RIOB33_X105Y111_IOB_X1Y111_I),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(CLBLL_L_X2Y105_SLICE_X0Y105_AO6),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_BO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha55aa55a63c663c6)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_ALUT (
.I0(CLBLL_L_X2Y103_SLICE_X0Y103_DO6),
.I1(CLBLL_L_X2Y105_SLICE_X0Y105_BO6),
.I2(CLBLL_L_X2Y106_SLICE_X0Y106_BO6),
.I3(CLBLM_R_X3Y103_SLICE_X2Y103_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_AO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_DO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_CO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_BO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_AO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_DO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_CO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_BO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h500010005ca09ca0)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_ALUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_AO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_DO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_CO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_BO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_AO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb4783cf0d21e965a)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_DLUT (
.I0(CLBLL_L_X2Y111_SLICE_X0Y111_AO6),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(CLBLL_L_X2Y111_SLICE_X1Y111_BO6),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(CLBLL_L_X2Y112_SLICE_X0Y112_AO6),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_DO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h460f0aa075f00aa0)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_CLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_CO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h072588aa5af00aa0)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_BLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_BO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88887777ff00ff77)
  ) CLBLL_L_X2Y111_SLICE_X0Y111_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(1'b1),
.I3(CLBLL_L_X2Y110_SLICE_X0Y110_AO6),
.I4(CLBLL_L_X2Y111_SLICE_X0Y111_CO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X0Y111_AO5),
.O6(CLBLL_L_X2Y111_SLICE_X0Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbaba00ba00ffba)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_DLUT (
.I0(CLBLL_L_X2Y110_SLICE_X0Y110_AO6),
.I1(CLBLL_L_X2Y111_SLICE_X0Y111_CO6),
.I2(CLBLL_L_X2Y112_SLICE_X1Y112_AO5),
.I3(CLBLL_L_X2Y111_SLICE_X1Y111_AO5),
.I4(CLBLM_R_X3Y110_SLICE_X2Y110_AO6),
.I5(CLBLM_R_X3Y111_SLICE_X3Y111_AO5),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_DO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha6599a9a659a9a9a)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_CLUT (
.I0(CLBLM_R_X3Y111_SLICE_X2Y111_BO6),
.I1(CLBLL_L_X2Y111_SLICE_X0Y111_AO5),
.I2(CLBLM_R_X3Y111_SLICE_X2Y111_AO6),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_CO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h66669996aaaa5a5a)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_BLUT (
.I0(CLBLM_R_X3Y110_SLICE_X2Y110_AO6),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(CLBLL_L_X2Y111_SLICE_X0Y111_CO6),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(CLBLL_L_X2Y110_SLICE_X0Y110_AO6),
.I5(LIOB33_X0Y101_IOB_X0Y101_I),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_BO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777777755ff55ff)
  ) CLBLL_L_X2Y111_SLICE_X1Y111_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y111_SLICE_X1Y111_AO5),
.O6(CLBLL_L_X2Y111_SLICE_X1Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h007a0050808aa0a0)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_DLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_DO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c6c93936c6cc66c)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_CLUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(CLBLL_L_X2Y111_SLICE_X0Y111_CO6),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(CLBLL_L_X2Y112_SLICE_X0Y112_DO6),
.I5(CLBLL_L_X2Y111_SLICE_X0Y111_BO6),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_CO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ffcc0033ff)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_BLUT (
.I0(1'b1),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(1'b1),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(CLBLL_L_X2Y112_SLICE_X0Y112_CO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_BO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haabbaaffcc3300ff)
  ) CLBLL_L_X2Y112_SLICE_X0Y112_ALUT (
.I0(CLBLL_L_X2Y112_SLICE_X0Y112_DO6),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(1'b1),
.I3(CLBLL_L_X2Y111_SLICE_X0Y111_BO6),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.O6(CLBLL_L_X2Y112_SLICE_X0Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcf3c030fefbc832)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_DLUT (
.I0(CLBLL_L_X2Y112_SLICE_X1Y112_AO6),
.I1(CLBLL_L_X2Y111_SLICE_X0Y111_CO6),
.I2(CLBLL_L_X2Y112_SLICE_X0Y112_DO6),
.I3(CLBLL_L_X2Y112_SLICE_X1Y112_AO5),
.I4(CLBLL_L_X2Y112_SLICE_X0Y112_BO6),
.I5(CLBLL_L_X2Y111_SLICE_X0Y111_BO6),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_DO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fdf134cdfdf4c4c)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_CLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(CLBLL_L_X2Y111_SLICE_X1Y111_BO6),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(CLBLL_L_X2Y112_SLICE_X1Y112_DO6),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_CO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a95c03f956a3fc0)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(CLBLL_L_X2Y111_SLICE_X1Y111_CO6),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(CLBLL_L_X2Y112_SLICE_X1Y112_CO6),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_BO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff0f0fffff)
  ) CLBLL_L_X2Y112_SLICE_X1Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y112_SLICE_X1Y112_AO5),
.O6(CLBLL_L_X2Y112_SLICE_X1Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_DO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_CO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_BO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f0003f3f3f3f)
  ) CLBLL_L_X2Y113_SLICE_X0Y113_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X0Y113_AO5),
.O6(CLBLL_L_X2Y113_SLICE_X0Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_DO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_CO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_BO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y113_SLICE_X1Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y113_SLICE_X1Y113_AO5),
.O6(CLBLL_L_X2Y113_SLICE_X1Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y101_SLICE_X4Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y101_SLICE_X4Y101_DO5),
.O6(CLBLL_L_X4Y101_SLICE_X4Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0445ddff5ddfddff)
  ) CLBLL_L_X4Y101_SLICE_X4Y101_CLUT (
.I0(CLBLL_L_X4Y101_SLICE_X5Y101_BO6),
.I1(CLBLM_R_X5Y101_SLICE_X7Y101_CO6),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(CLBLL_L_X4Y101_SLICE_X4Y101_AO5),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLL_L_X4Y101_SLICE_X4Y101_CO5),
.O6(CLBLL_L_X4Y101_SLICE_X4Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he62a19d573bf8c40)
  ) CLBLL_L_X4Y101_SLICE_X4Y101_BLUT (
.I0(CLBLM_R_X5Y101_SLICE_X7Y101_CO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(CLBLL_L_X4Y101_SLICE_X5Y101_BO6),
.I5(CLBLL_L_X4Y101_SLICE_X4Y101_AO5),
.O5(CLBLL_L_X4Y101_SLICE_X4Y101_BO5),
.O6(CLBLL_L_X4Y101_SLICE_X4Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h956a6a953fc0c03f)
  ) CLBLL_L_X4Y101_SLICE_X4Y101_ALUT (
.I0(CLBLM_R_X5Y101_SLICE_X7Y101_CO6),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(CLBLM_R_X5Y101_SLICE_X7Y101_AO5),
.I4(CLBLM_R_X5Y100_SLICE_X6Y100_AO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y101_SLICE_X4Y101_AO5),
.O6(CLBLL_L_X4Y101_SLICE_X4Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f037f1f7f13ffff)
  ) CLBLL_L_X4Y101_SLICE_X5Y101_DLUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(CLBLM_R_X5Y101_SLICE_X6Y101_BO6),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(CLBLM_R_X5Y101_SLICE_X7Y101_DO6),
.I4(CLBLM_R_X5Y101_SLICE_X6Y101_CO6),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLL_L_X4Y101_SLICE_X5Y101_DO5),
.O6(CLBLL_L_X4Y101_SLICE_X5Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8fe3701c7f1380ec)
  ) CLBLL_L_X4Y101_SLICE_X5Y101_CLUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(CLBLM_R_X5Y101_SLICE_X6Y101_BO6),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(CLBLM_R_X5Y101_SLICE_X7Y101_DO6),
.I4(CLBLM_R_X5Y101_SLICE_X6Y101_CO6),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLL_L_X4Y101_SLICE_X5Y101_CO5),
.O6(CLBLL_L_X4Y101_SLICE_X5Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb87b787747848788)
  ) CLBLL_L_X4Y101_SLICE_X5Y101_BLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(CLBLM_R_X5Y100_SLICE_X6Y100_AO6),
.I3(CLBLM_R_X5Y101_SLICE_X7Y101_AO5),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLL_L_X4Y101_SLICE_X5Y101_CO6),
.O5(CLBLL_L_X4Y101_SLICE_X5Y101_BO5),
.O6(CLBLL_L_X4Y101_SLICE_X5Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1051f3f375f7ffff)
  ) CLBLL_L_X4Y101_SLICE_X5Y101_ALUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(CLBLM_R_X5Y101_SLICE_X7Y101_AO5),
.I2(CLBLM_R_X5Y100_SLICE_X6Y100_AO6),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(CLBLL_L_X4Y101_SLICE_X5Y101_CO6),
.O5(CLBLL_L_X4Y101_SLICE_X5Y101_AO5),
.O6(CLBLL_L_X4Y101_SLICE_X5Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h157fffff015733ff)
  ) CLBLL_L_X4Y102_SLICE_X4Y102_DLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(CLBLL_L_X4Y102_SLICE_X5Y102_AO6),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(CLBLL_L_X4Y102_SLICE_X4Y102_CO6),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(CLBLL_L_X4Y101_SLICE_X5Y101_DO6),
.O5(CLBLL_L_X4Y102_SLICE_X4Y102_DO5),
.O6(CLBLL_L_X4Y102_SLICE_X4Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb3cb7f074c3480f8)
  ) CLBLL_L_X4Y102_SLICE_X4Y102_CLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(CLBLL_L_X4Y103_SLICE_X5Y103_BO6),
.I3(CLBLM_R_X5Y101_SLICE_X6Y101_AO5),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(CLBLM_R_X3Y102_SLICE_X2Y102_BO6),
.O5(CLBLL_L_X4Y102_SLICE_X4Y102_CO5),
.O6(CLBLL_L_X4Y102_SLICE_X4Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f7f5fff035f137f)
  ) CLBLL_L_X4Y102_SLICE_X4Y102_BLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(CLBLL_L_X4Y103_SLICE_X5Y103_BO6),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(CLBLM_R_X3Y102_SLICE_X2Y102_BO6),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLM_R_X5Y101_SLICE_X6Y101_AO5),
.O5(CLBLL_L_X4Y102_SLICE_X4Y102_BO5),
.O6(CLBLL_L_X4Y102_SLICE_X4Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffff78877887)
  ) CLBLL_L_X4Y102_SLICE_X4Y102_ALUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(RIOB33_X105Y107_IOB_X1Y108_I),
.I2(CLBLL_L_X4Y102_SLICE_X5Y102_AO6),
.I3(CLBLL_L_X4Y101_SLICE_X5Y101_DO6),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y102_SLICE_X4Y102_AO5),
.O6(CLBLL_L_X4Y102_SLICE_X4Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hbc70d61acc000cc0)
  ) CLBLL_L_X4Y102_SLICE_X5Y102_DLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(CLBLM_R_X5Y102_SLICE_X6Y102_CO6),
.I5(RIOB33_X105Y111_IOB_X1Y111_I),
.O5(CLBLL_L_X4Y102_SLICE_X5Y102_DO5),
.O6(CLBLL_L_X4Y102_SLICE_X5Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'he86ac6cc24a60a00)
  ) CLBLL_L_X4Y102_SLICE_X5Y102_CLUT (
.I0(RIOB33_X105Y111_IOB_X1Y111_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(CLBLM_R_X3Y102_SLICE_X3Y102_BO6),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLL_L_X4Y102_SLICE_X5Y102_CO5),
.O6(CLBLL_L_X4Y102_SLICE_X5Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcebb73ff63ff33ff)
  ) CLBLL_L_X4Y102_SLICE_X5Y102_BLUT (
.I0(CLBLM_R_X3Y102_SLICE_X3Y102_BO6),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(RIOB33_X105Y109_IOB_X1Y110_I),
.O5(CLBLL_L_X4Y102_SLICE_X5Y102_BO5),
.O6(CLBLL_L_X4Y102_SLICE_X5Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33c996633cc)
  ) CLBLL_L_X4Y102_SLICE_X5Y102_ALUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(CLBLM_R_X5Y101_SLICE_X6Y101_AO5),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(CLBLL_L_X4Y102_SLICE_X5Y102_BO6),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(RIOB33_X105Y109_IOB_X1Y110_I),
.O5(CLBLL_L_X4Y102_SLICE_X5Y102_AO5),
.O6(CLBLL_L_X4Y102_SLICE_X5Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he619758a4cb3df20)
  ) CLBLL_L_X4Y103_SLICE_X4Y103_DLUT (
.I0(RIOB33_X105Y107_IOB_X1Y108_I),
.I1(CLBLL_L_X4Y101_SLICE_X5Y101_DO6),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(CLBLL_L_X4Y102_SLICE_X4Y102_CO6),
.I4(CLBLL_L_X4Y102_SLICE_X5Y102_AO6),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLL_L_X4Y103_SLICE_X4Y103_DO5),
.O6(CLBLL_L_X4Y103_SLICE_X4Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9fc53f95603ac06a)
  ) CLBLL_L_X4Y103_SLICE_X4Y103_CLUT (
.I0(CLBLL_L_X4Y104_SLICE_X5Y104_AO6),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(CLBLM_R_X5Y104_SLICE_X6Y104_AO5),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(CLBLL_L_X4Y104_SLICE_X5Y104_BO6),
.O5(CLBLL_L_X4Y103_SLICE_X4Y103_CO5),
.O6(CLBLL_L_X4Y103_SLICE_X4Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f66cc9933)
  ) CLBLL_L_X4Y103_SLICE_X4Y103_BLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(CLBLL_L_X4Y102_SLICE_X4Y102_AO5),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(CLBLL_L_X4Y101_SLICE_X5Y101_AO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y103_SLICE_X4Y103_BO5),
.O6(CLBLL_L_X4Y103_SLICE_X4Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff6699aa55)
  ) CLBLL_L_X4Y103_SLICE_X4Y103_ALUT (
.I0(CLBLL_L_X2Y103_SLICE_X1Y103_BO6),
.I1(LIOB33_X0Y113_IOB_X0Y113_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLL_L_X4Y102_SLICE_X4Y102_DO6),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y103_SLICE_X4Y103_AO5),
.O6(CLBLL_L_X4Y103_SLICE_X4Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y103_SLICE_X5Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y103_SLICE_X5Y103_DO5),
.O6(CLBLL_L_X4Y103_SLICE_X5Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f13ff5fdf4c5f00)
  ) CLBLL_L_X4Y103_SLICE_X5Y103_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLL_L_X4Y103_SLICE_X5Y103_AO5),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(CLBLL_L_X4Y104_SLICE_X5Y104_BO6),
.O5(CLBLL_L_X4Y103_SLICE_X5Y103_CO5),
.O6(CLBLL_L_X4Y103_SLICE_X5Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc3333330fff0fff)
  ) CLBLL_L_X4Y103_SLICE_X5Y103_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y102_SLICE_X5Y102_BO6),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y103_SLICE_X5Y103_BO5),
.O6(CLBLL_L_X4Y103_SLICE_X5Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff2baf2baf)
  ) CLBLL_L_X4Y103_SLICE_X5Y103_ALUT (
.I0(CLBLM_R_X5Y104_SLICE_X6Y104_AO5),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(CLBLL_L_X4Y104_SLICE_X5Y104_AO6),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y103_SLICE_X5Y103_AO5),
.O6(CLBLL_L_X4Y103_SLICE_X5Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f7f151f7f7f157f)
  ) CLBLL_L_X4Y104_SLICE_X4Y104_DLUT (
.I0(CLBLL_L_X4Y101_SLICE_X4Y101_BO6),
.I1(LIOB33_X0Y113_IOB_X0Y113_I),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(CLBLL_L_X4Y104_SLICE_X4Y104_AO5),
.I4(CLBLM_R_X5Y105_SLICE_X7Y105_BO5),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLL_L_X4Y104_SLICE_X4Y104_DO5),
.O6(CLBLL_L_X4Y104_SLICE_X4Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9a6a959a6a6a956a)
  ) CLBLL_L_X4Y104_SLICE_X4Y104_CLUT (
.I0(CLBLL_L_X4Y101_SLICE_X4Y101_BO6),
.I1(LIOB33_X0Y113_IOB_X0Y113_I),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(CLBLL_L_X4Y104_SLICE_X4Y104_AO5),
.I4(CLBLM_R_X5Y105_SLICE_X7Y105_BO5),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLL_L_X4Y104_SLICE_X4Y104_CO5),
.O6(CLBLL_L_X4Y104_SLICE_X4Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aaaa5550aaaafff)
  ) CLBLL_L_X4Y104_SLICE_X4Y104_BLUT (
.I0(CLBLL_L_X4Y105_SLICE_X4Y105_CO6),
.I1(1'b1),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(CLBLL_L_X4Y104_SLICE_X4Y104_CO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y104_SLICE_X4Y104_BO5),
.O6(CLBLL_L_X4Y104_SLICE_X4Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a569a5c30fc30f)
  ) CLBLL_L_X4Y104_SLICE_X4Y104_ALUT (
.I0(CLBLM_R_X5Y105_SLICE_X7Y105_BO5),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(CLBLL_L_X4Y101_SLICE_X4Y101_AO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y104_SLICE_X4Y104_AO5),
.O6(CLBLL_L_X4Y104_SLICE_X4Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9f603fc0c53a956a)
  ) CLBLL_L_X4Y104_SLICE_X5Y104_DLUT (
.I0(CLBLL_L_X4Y104_SLICE_X5Y104_AO6),
.I1(LIOB33_X0Y113_IOB_X0Y113_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLL_L_X4Y104_SLICE_X5Y104_CO6),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(CLBLM_R_X5Y104_SLICE_X6Y104_AO5),
.O5(CLBLL_L_X4Y104_SLICE_X5Y104_DO5),
.O6(CLBLL_L_X4Y104_SLICE_X5Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999666996669996)
  ) CLBLL_L_X4Y104_SLICE_X5Y104_CLUT (
.I0(CLBLL_L_X4Y106_SLICE_X5Y106_AO6),
.I1(CLBLM_R_X3Y105_SLICE_X3Y105_CO6),
.I2(CLBLM_R_X5Y103_SLICE_X6Y103_AO5),
.I3(CLBLL_L_X4Y104_SLICE_X5Y104_AO5),
.I4(CLBLM_R_X5Y105_SLICE_X7Y105_CO6),
.I5(CLBLM_R_X5Y102_SLICE_X6Y102_AO6),
.O5(CLBLL_L_X4Y104_SLICE_X5Y104_CO5),
.O6(CLBLL_L_X4Y104_SLICE_X5Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb24d4db2dd22dd22)
  ) CLBLL_L_X4Y104_SLICE_X5Y104_BLUT (
.I0(CLBLM_R_X5Y105_SLICE_X7Y105_CO6),
.I1(CLBLM_R_X5Y103_SLICE_X6Y103_AO5),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(CLBLM_R_X5Y102_SLICE_X6Y102_AO6),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLL_L_X4Y104_SLICE_X5Y104_BO5),
.O6(CLBLL_L_X4Y104_SLICE_X5Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h699969990fff0fff)
  ) CLBLL_L_X4Y104_SLICE_X5Y104_ALUT (
.I0(CLBLM_R_X5Y105_SLICE_X7Y105_CO6),
.I1(CLBLM_R_X5Y103_SLICE_X6Y103_AO5),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y104_SLICE_X5Y104_AO5),
.O6(CLBLL_L_X4Y104_SLICE_X5Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha8feffff0000a8fe)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_DLUT (
.I0(CLBLL_L_X4Y105_SLICE_X4Y105_AO6),
.I1(CLBLL_L_X4Y105_SLICE_X5Y105_CO6),
.I2(CLBLL_L_X4Y107_SLICE_X5Y107_DO6),
.I3(CLBLM_R_X3Y105_SLICE_X3Y105_DO6),
.I4(CLBLL_L_X4Y104_SLICE_X4Y104_BO6),
.I5(CLBLL_L_X4Y105_SLICE_X4Y105_BO6),
.O5(CLBLL_L_X4Y105_SLICE_X4Y105_DO5),
.O6(CLBLL_L_X4Y105_SLICE_X4Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h60f6f6f6a0fafafa)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_CLUT (
.I0(CLBLL_L_X4Y104_SLICE_X4Y104_AO6),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(CLBLL_L_X4Y105_SLICE_X5Y105_BO6),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLL_L_X4Y105_SLICE_X4Y105_CO5),
.O6(CLBLL_L_X4Y105_SLICE_X4Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6cffffff006c6c6c)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(CLBLM_R_X3Y105_SLICE_X3Y105_AO5),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLL_L_X4Y103_SLICE_X5Y103_CO6),
.O5(CLBLL_L_X4Y105_SLICE_X4Y105_BO5),
.O6(CLBLL_L_X4Y105_SLICE_X4Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4dddcfff8eee0ccc)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(CLBLM_R_X5Y103_SLICE_X6Y103_CO6),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(CLBLL_L_X4Y103_SLICE_X4Y103_CO6),
.O5(CLBLL_L_X4Y105_SLICE_X4Y105_AO5),
.O6(CLBLL_L_X4Y105_SLICE_X4Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4bd2b42db42d4bd2)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_DLUT (
.I0(CLBLM_R_X3Y106_SLICE_X3Y106_AO5),
.I1(CLBLM_R_X5Y103_SLICE_X6Y103_DO6),
.I2(CLBLL_L_X4Y104_SLICE_X5Y104_DO6),
.I3(CLBLL_L_X4Y105_SLICE_X5Y105_AO5),
.I4(CLBLL_L_X4Y105_SLICE_X5Y105_AO6),
.I5(CLBLM_R_X5Y103_SLICE_X6Y103_CO6),
.O5(CLBLL_L_X4Y105_SLICE_X5Y105_DO5),
.O6(CLBLL_L_X4Y105_SLICE_X5Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0b02b020b0200b02)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_CLUT (
.I0(CLBLM_R_X3Y106_SLICE_X3Y106_AO5),
.I1(CLBLM_R_X5Y103_SLICE_X6Y103_DO6),
.I2(CLBLL_L_X4Y104_SLICE_X5Y104_DO6),
.I3(CLBLL_L_X4Y105_SLICE_X5Y105_AO5),
.I4(CLBLL_L_X4Y105_SLICE_X5Y105_AO6),
.I5(CLBLM_R_X5Y103_SLICE_X6Y103_CO6),
.O5(CLBLL_L_X4Y105_SLICE_X5Y105_CO5),
.O6(CLBLL_L_X4Y105_SLICE_X5Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1301ff557f37ffff)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_BLUT (
.I0(CLBLM_R_X5Y105_SLICE_X7Y105_CO6),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(CLBLM_R_X5Y103_SLICE_X6Y103_AO5),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(CLBLM_R_X5Y105_SLICE_X7Y105_BO6),
.O5(CLBLL_L_X4Y105_SLICE_X5Y105_BO5),
.O6(CLBLL_L_X4Y105_SLICE_X5Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f0fff0fff)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(1'b1),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y105_SLICE_X5Y105_AO5),
.O6(CLBLL_L_X4Y105_SLICE_X5Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb3fb32b332b32032)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_DLUT (
.I0(CLBLM_R_X5Y103_SLICE_X6Y103_CO6),
.I1(CLBLM_R_X3Y105_SLICE_X3Y105_DO6),
.I2(CLBLL_L_X4Y106_SLICE_X5Y106_DO6),
.I3(CLBLL_L_X4Y104_SLICE_X5Y104_DO6),
.I4(CLBLL_L_X4Y107_SLICE_X4Y107_DO6),
.I5(CLBLL_L_X4Y105_SLICE_X5Y105_AO6),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_DO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c939393936c6c6c)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(CLBLM_R_X5Y103_SLICE_X6Y103_CO6),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLL_L_X4Y103_SLICE_X4Y103_CO6),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_CO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h96969696b24d4db2)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_BLUT (
.I0(CLBLL_L_X4Y107_SLICE_X4Y107_DO6),
.I1(CLBLL_L_X4Y106_SLICE_X4Y106_CO6),
.I2(CLBLL_L_X4Y106_SLICE_X5Y106_DO6),
.I3(CLBLM_R_X3Y105_SLICE_X3Y105_DO6),
.I4(CLBLL_L_X4Y105_SLICE_X4Y105_AO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_BO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h30f3f0ff3cc3f00f)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(CLBLM_R_X5Y106_SLICE_X6Y106_BO6),
.I3(CLBLM_R_X5Y105_SLICE_X6Y105_CO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_AO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h71f3f5ffd4fc50f0)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_DLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(CLBLM_R_X3Y106_SLICE_X3Y106_AO5),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(CLBLM_R_X5Y104_SLICE_X6Y104_BO6),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_DO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887878787787878)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_R_X3Y106_SLICE_X3Y106_AO5),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(CLBLM_R_X5Y104_SLICE_X6Y104_BO6),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_CO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f15ff3fd540ffc0)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(CLBLM_R_X5Y107_SLICE_X6Y107_DO6),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLM_R_X5Y106_SLICE_X6Y106_DO6),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_BO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff0f0fffff)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_AO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000e880fee8fffe)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_DLUT (
.I0(CLBLL_L_X4Y106_SLICE_X5Y106_BO6),
.I1(CLBLL_L_X4Y107_SLICE_X5Y107_AO5),
.I2(CLBLM_R_X5Y107_SLICE_X6Y107_CO6),
.I3(CLBLM_R_X3Y107_SLICE_X3Y107_BO6),
.I4(CLBLM_R_X3Y107_SLICE_X2Y107_AO5),
.I5(CLBLL_L_X4Y106_SLICE_X5Y106_CO6),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_DO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4dcfd4fcd4fcd4fc)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLM_R_X5Y107_SLICE_X6Y107_CO6),
.I2(CLBLM_R_X3Y107_SLICE_X3Y107_DO5),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_CO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a95956a956a956a)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_BLUT (
.I0(CLBLM_R_X5Y107_SLICE_X6Y107_CO6),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(CLBLM_R_X3Y107_SLICE_X3Y107_DO5),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_BO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc639639ca5a55a5a)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_ALUT (
.I0(CLBLL_L_X4Y107_SLICE_X4Y107_BO6),
.I1(CLBLL_L_X4Y107_SLICE_X4Y107_CO6),
.I2(CLBLM_R_X3Y107_SLICE_X3Y107_BO6),
.I3(CLBLL_L_X4Y106_SLICE_X5Y106_CO6),
.I4(CLBLL_L_X4Y106_SLICE_X5Y106_BO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_AO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00dd004d004d0044)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_DLUT (
.I0(CLBLL_L_X4Y106_SLICE_X5Y106_CO6),
.I1(CLBLL_L_X4Y107_SLICE_X4Y107_CO6),
.I2(CLBLL_L_X4Y107_SLICE_X4Y107_BO6),
.I3(CLBLL_L_X4Y105_SLICE_X5Y105_DO6),
.I4(CLBLL_L_X4Y106_SLICE_X5Y106_BO6),
.I5(CLBLM_R_X3Y107_SLICE_X3Y107_BO6),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_DO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1171f3f37177ffff)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(CLBLM_R_X5Y107_SLICE_X7Y107_AO6),
.I2(CLBLL_L_X4Y108_SLICE_X4Y108_DO6),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLM_R_X5Y107_SLICE_X6Y107_AO6),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_CO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c939393936c6c6c)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLM_R_X5Y106_SLICE_X6Y106_DO6),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLM_R_X5Y107_SLICE_X6Y107_DO6),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_BO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffff00ffffff)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(1'b1),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_AO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7080f7f8f7f8f7f8)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_DLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(CLBLM_R_X5Y109_SLICE_X6Y109_DO6),
.I3(CLBLM_R_X7Y108_SLICE_X8Y108_CO6),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_DO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0708080777888877)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_CLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(CLBLM_R_X7Y108_SLICE_X8Y108_CO6),
.I4(CLBLM_R_X5Y109_SLICE_X6Y109_DO6),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_CO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a9696a5a569695a)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_BLUT (
.I0(CLBLM_R_X7Y109_SLICE_X8Y109_CO6),
.I1(CLBLM_R_X5Y109_SLICE_X6Y109_AO6),
.I2(CLBLM_R_X3Y105_SLICE_X3Y105_AO6),
.I3(CLBLM_R_X5Y110_SLICE_X7Y110_BO6),
.I4(CLBLL_L_X4Y108_SLICE_X4Y108_AO6),
.I5(CLBLL_L_X4Y108_SLICE_X4Y108_AO5),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_BO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff77777777)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_ALUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_AO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc66c66cc9933c66c)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_DLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(CLBLM_R_X5Y107_SLICE_X7Y107_CO6),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(CLBLM_R_X5Y107_SLICE_X6Y107_AO6),
.I5(CLBLL_L_X4Y108_SLICE_X4Y108_DO6),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_DO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffb3ff135f20a0)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(CLBLL_L_X4Y108_SLICE_X5Y108_DO6),
.I5(CLBLM_R_X5Y108_SLICE_X6Y108_CO6),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_CO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h87787887e11e1ee1)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_BLUT (
.I0(CLBLM_R_X3Y102_SLICE_X3Y102_AO6),
.I1(CLBLL_L_X4Y109_SLICE_X4Y109_DO6),
.I2(CLBLL_L_X4Y107_SLICE_X5Y107_AO6),
.I3(CLBLM_R_X5Y108_SLICE_X6Y108_CO6),
.I4(CLBLL_L_X4Y108_SLICE_X5Y108_AO6),
.I5(CLBLM_R_X5Y108_SLICE_X6Y108_BO6),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_BO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb78b487477878878)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(CLBLM_R_X5Y107_SLICE_X6Y107_AO6),
.I3(CLBLL_L_X4Y108_SLICE_X4Y108_DO6),
.I4(CLBLM_R_X5Y107_SLICE_X7Y107_AO6),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_AO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f7f05157fff1fff)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_DLUT (
.I0(CLBLL_L_X4Y109_SLICE_X4Y109_AO6),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(CLBLM_R_X3Y110_SLICE_X3Y110_BO6),
.I5(CLBLL_L_X4Y108_SLICE_X4Y108_BO6),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_DO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h956aff00a9560ff0)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(CLBLM_R_X5Y109_SLICE_X6Y109_AO6),
.I3(CLBLM_R_X7Y109_SLICE_X8Y109_CO6),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(CLBLM_R_X5Y110_SLICE_X7Y110_BO6),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_CO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hca6a6f3f359590c0)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_BLUT (
.I0(CLBLM_R_X3Y110_SLICE_X3Y110_BO6),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(CLBLL_L_X4Y109_SLICE_X4Y109_AO6),
.I5(CLBLL_L_X4Y109_SLICE_X4Y109_CO6),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_BO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887877887788778)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_ALUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(CLBLM_R_X7Y109_SLICE_X8Y109_AO6),
.I3(CLBLM_R_X5Y110_SLICE_X7Y110_BO6),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_AO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_DO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_CO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_BO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ca0935f935f6ca0)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_ALUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(LIOB33_X0Y113_IOB_X0Y113_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(CLBLL_L_X4Y109_SLICE_X4Y109_DO6),
.I5(CLBLM_R_X5Y109_SLICE_X6Y109_BO6),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_AO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c39933963c66cc)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(CLBLM_R_X5Y111_SLICE_X7Y111_AO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLL_L_X4Y113_SLICE_X5Y113_BO6),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_DO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb43cd29678f01e5a)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_CLUT (
.I0(CLBLL_L_X4Y111_SLICE_X4Y111_AO6),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(CLBLL_L_X4Y111_SLICE_X5Y111_DO6),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_AO5),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_CO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000064e48808a828)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_BLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(RIOB33_X105Y111_IOB_X1Y112_I),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_BO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3c33333ff03ff33)
  ) CLBLL_L_X4Y111_SLICE_X4Y111_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y110_SLICE_X2Y110_BO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLL_L_X4Y111_SLICE_X4Y111_BO6),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y111_SLICE_X4Y111_AO5),
.O6(CLBLL_L_X4Y111_SLICE_X4Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ef1f50af10ef50a)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_DLUT (
.I0(CLBLM_R_X3Y110_SLICE_X2Y110_BO6),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(CLBLL_L_X4Y111_SLICE_X4Y111_BO6),
.I3(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_DO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaa0a0fafea8a8fe)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_CLUT (
.I0(CLBLL_L_X4Y111_SLICE_X5Y111_AO6),
.I1(CLBLM_R_X3Y111_SLICE_X3Y111_AO6),
.I2(CLBLL_L_X4Y111_SLICE_X4Y111_BO6),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_AO6),
.I4(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I5(CLBLM_R_X3Y110_SLICE_X2Y110_BO6),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_CO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h55aaaa559a65659a)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_BLUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I1(CLBLM_R_X3Y110_SLICE_X2Y110_BO6),
.I2(CLBLM_R_X3Y111_SLICE_X3Y111_AO6),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_AO6),
.I4(CLBLL_L_X4Y111_SLICE_X5Y111_AO6),
.I5(CLBLL_L_X4Y111_SLICE_X4Y111_BO6),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_BO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555ffff5f5f5f5f)
  ) CLBLL_L_X4Y111_SLICE_X5Y111_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(1'b1),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(1'b1),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y111_SLICE_X5Y111_AO5),
.O6(CLBLL_L_X4Y111_SLICE_X5Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a5c30f965a3cf0)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_DLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(CLBLL_L_X4Y111_SLICE_X5Y111_DO6),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLM_R_X3Y111_SLICE_X2Y111_CO6),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_DO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h96f03cf0c30f96f0)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y106_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(CLBLL_L_X4Y112_SLICE_X5Y112_BO6),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_DO6),
.I5(CLBLM_R_X3Y112_SLICE_X2Y112_CO6),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_CO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6696996996996966)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_BLUT (
.I0(CLBLM_R_X3Y111_SLICE_X2Y111_CO6),
.I1(CLBLL_L_X4Y111_SLICE_X5Y111_BO6),
.I2(CLBLM_R_X3Y111_SLICE_X2Y111_DO6),
.I3(CLBLL_L_X2Y111_SLICE_X1Y111_DO6),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_AO6),
.I5(CLBLL_L_X4Y112_SLICE_X4Y112_AO5),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_BO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h777777775f5f5f5f)
  ) CLBLL_L_X4Y112_SLICE_X4Y112_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y112_SLICE_X4Y112_AO5),
.O6(CLBLL_L_X4Y112_SLICE_X4Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hefae8a088a08efae)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_DLUT (
.I0(CLBLL_L_X4Y112_SLICE_X5Y112_AO6),
.I1(CLBLM_R_X3Y113_SLICE_X2Y113_BO6),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_DO6),
.I3(CLBLM_R_X3Y112_SLICE_X2Y112_CO6),
.I4(CLBLL_L_X4Y112_SLICE_X5Y112_BO6),
.I5(CLBLM_R_X5Y112_SLICE_X6Y112_AO6),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_DO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7d14f550ff3cfff0)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(CLBLL_L_X4Y111_SLICE_X5Y111_DO6),
.I3(CLBLM_R_X3Y111_SLICE_X2Y111_CO6),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_CO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6966969999696696)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_BLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_AO6),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_BO6),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_AO6),
.I3(CLBLL_L_X4Y111_SLICE_X5Y111_BO6),
.I4(CLBLL_L_X4Y111_SLICE_X5Y111_CO6),
.I5(CLBLM_R_X3Y111_SLICE_X2Y111_CO6),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_BO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff00ffffff)
  ) CLBLL_L_X4Y112_SLICE_X5Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y112_SLICE_X5Y112_AO5),
.O6(CLBLL_L_X4Y112_SLICE_X5Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_DO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_CO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fbfff3f152a3f00)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(CLBLL_L_X4Y111_SLICE_X4Y111_CO6),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(CLBLM_R_X3Y112_SLICE_X2Y112_CO6),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_BO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb78b778748748878)
  ) CLBLL_L_X4Y113_SLICE_X4Y113_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(CLBLL_L_X4Y113_SLICE_X5Y113_AO6),
.I3(CLBLL_L_X4Y113_SLICE_X4Y113_BO6),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(CLBLM_R_X5Y112_SLICE_X6Y112_CO6),
.O5(CLBLL_L_X4Y113_SLICE_X4Y113_AO5),
.O6(CLBLL_L_X4Y113_SLICE_X4Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_DO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_CO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4d8ecf0cddeeffcc)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(CLBLL_L_X4Y112_SLICE_X5Y112_DO6),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(CLBLM_R_X5Y112_SLICE_X6Y112_CO6),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_BO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887878787787878)
  ) CLBLL_L_X4Y113_SLICE_X5Y113_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(CLBLM_R_X5Y112_SLICE_X7Y112_AO6),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLL_L_X4Y112_SLICE_X5Y112_CO6),
.O5(CLBLL_L_X4Y113_SLICE_X5Y113_AO5),
.O6(CLBLL_L_X4Y113_SLICE_X5Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y101_SLICE_X10Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y101_SLICE_X10Y101_DO5),
.O6(CLBLM_L_X8Y101_SLICE_X10Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y101_SLICE_X10Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y101_SLICE_X10Y101_CO5),
.O6(CLBLM_L_X8Y101_SLICE_X10Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y101_SLICE_X10Y101_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y101_SLICE_X10Y101_BO5),
.O6(CLBLM_L_X8Y101_SLICE_X10Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h57157f1f5f17ff3f)
  ) CLBLM_L_X8Y101_SLICE_X10Y101_ALUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(CLBLM_L_X8Y103_SLICE_X10Y103_BO6),
.I2(CLBLM_R_X7Y101_SLICE_X9Y101_BO6),
.I3(CLBLM_L_X10Y101_SLICE_X12Y101_BO6),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_L_X8Y101_SLICE_X10Y101_AO5),
.O6(CLBLM_L_X8Y101_SLICE_X10Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y101_SLICE_X11Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y101_SLICE_X11Y101_DO5),
.O6(CLBLM_L_X8Y101_SLICE_X11Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y101_SLICE_X11Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y101_SLICE_X11Y101_CO5),
.O6(CLBLM_L_X8Y101_SLICE_X11Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y101_SLICE_X11Y101_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y101_SLICE_X11Y101_BO5),
.O6(CLBLM_L_X8Y101_SLICE_X11Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y101_SLICE_X11Y101_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y101_SLICE_X11Y101_AO5),
.O6(CLBLM_L_X8Y101_SLICE_X11Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha96965a56a66a6aa)
  ) CLBLM_L_X8Y102_SLICE_X10Y102_DLUT (
.I0(CLBLM_R_X7Y102_SLICE_X9Y102_CO6),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(CLBLM_L_X10Y101_SLICE_X12Y101_BO6),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(CLBLM_L_X8Y103_SLICE_X10Y103_BO6),
.O5(CLBLM_L_X8Y102_SLICE_X10Y102_DO5),
.O6(CLBLM_L_X8Y102_SLICE_X10Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf80bbbb82dd7777)
  ) CLBLM_L_X8Y102_SLICE_X10Y102_CLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(RIOB33_X105Y109_IOB_X1Y109_I),
.O5(CLBLM_L_X8Y102_SLICE_X10Y102_CO5),
.O6(CLBLM_L_X8Y102_SLICE_X10Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9699aa556696aaaa)
  ) CLBLM_L_X8Y102_SLICE_X10Y102_BLUT (
.I0(CLBLM_L_X8Y102_SLICE_X10Y102_DO6),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y101_SLICE_X12Y101_CO6),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLM_L_X8Y102_SLICE_X10Y102_AO5),
.O5(CLBLM_L_X8Y102_SLICE_X10Y102_BO5),
.O6(CLBLM_L_X8Y102_SLICE_X10Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777777778877887)
  ) CLBLM_L_X8Y102_SLICE_X10Y102_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(CLBLM_L_X10Y101_SLICE_X12Y101_BO6),
.I3(CLBLM_L_X8Y103_SLICE_X10Y103_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y102_SLICE_X10Y102_AO5),
.O6(CLBLM_L_X8Y102_SLICE_X10Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f3f3f3f3f)
  ) CLBLM_L_X8Y102_SLICE_X11Y102_DLUT (
.I0(1'b1),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y102_SLICE_X11Y102_DO5),
.O6(CLBLM_L_X8Y102_SLICE_X11Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h666699c6cccc336c)
  ) CLBLM_L_X8Y102_SLICE_X11Y102_CLUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(CLBLM_L_X8Y102_SLICE_X10Y102_CO6),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(CLBLM_L_X10Y101_SLICE_X13Y101_AO6),
.I4(CLBLM_R_X7Y101_SLICE_X9Y101_CO6),
.I5(RIOB33_X105Y109_IOB_X1Y109_I),
.O5(CLBLM_L_X8Y102_SLICE_X11Y102_CO5),
.O6(CLBLM_L_X8Y102_SLICE_X11Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h59a69a65a659659a)
  ) CLBLM_L_X8Y102_SLICE_X11Y102_BLUT (
.I0(CLBLM_L_X8Y102_SLICE_X11Y102_DO6),
.I1(CLBLM_L_X8Y103_SLICE_X10Y103_BO6),
.I2(CLBLM_L_X8Y102_SLICE_X10Y102_AO6),
.I3(CLBLM_R_X7Y102_SLICE_X9Y102_CO6),
.I4(CLBLM_L_X10Y101_SLICE_X12Y101_BO6),
.I5(CLBLM_L_X10Y102_SLICE_X13Y102_AO5),
.O5(CLBLM_L_X8Y102_SLICE_X11Y102_BO5),
.O6(CLBLM_L_X8Y102_SLICE_X11Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hababbbbbc3c33333)
  ) CLBLM_L_X8Y102_SLICE_X11Y102_ALUT (
.I0(CLBLM_R_X7Y101_SLICE_X9Y101_CO6),
.I1(CLBLM_L_X10Y101_SLICE_X13Y101_AO6),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(1'b1),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y102_SLICE_X11Y102_AO5),
.O6(CLBLM_L_X8Y102_SLICE_X11Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0d4f0ddf4dffddff)
  ) CLBLM_L_X8Y103_SLICE_X10Y103_DLUT (
.I0(CLBLM_R_X7Y107_SLICE_X9Y107_BO6),
.I1(CLBLM_L_X8Y102_SLICE_X11Y102_AO6),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(CLBLM_L_X8Y103_SLICE_X10Y103_CO6),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_L_X8Y103_SLICE_X10Y103_DO5),
.O6(CLBLM_L_X8Y103_SLICE_X10Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ef1f30cf10ef30c)
  ) CLBLM_L_X8Y103_SLICE_X10Y103_CLUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(CLBLM_L_X8Y102_SLICE_X10Y102_CO6),
.I2(CLBLM_L_X8Y104_SLICE_X10Y104_DO6),
.I3(CLBLM_L_X8Y104_SLICE_X10Y104_CO6),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_L_X8Y103_SLICE_X10Y103_CO5),
.O6(CLBLM_L_X8Y103_SLICE_X10Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd57fad072a8052f8)
  ) CLBLM_L_X8Y103_SLICE_X10Y103_BLUT (
.I0(RIOB33_X105Y107_IOB_X1Y108_I),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_BO6),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLM_L_X8Y102_SLICE_X11Y102_AO6),
.I5(CLBLM_L_X8Y103_SLICE_X10Y103_CO6),
.O5(CLBLM_L_X8Y103_SLICE_X10Y103_BO5),
.O6(CLBLM_L_X8Y103_SLICE_X10Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a00ff6aff6aff6a)
  ) CLBLM_L_X8Y103_SLICE_X10Y103_ALUT (
.I0(CLBLM_L_X8Y102_SLICE_X10Y102_DO6),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(CLBLM_L_X10Y102_SLICE_X12Y102_CO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_L_X8Y103_SLICE_X10Y103_AO5),
.O6(CLBLM_L_X8Y103_SLICE_X10Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y103_SLICE_X11Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y103_SLICE_X11Y103_DO5),
.O6(CLBLM_L_X8Y103_SLICE_X11Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y103_SLICE_X11Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y103_SLICE_X11Y103_CO5),
.O6(CLBLM_L_X8Y103_SLICE_X11Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y103_SLICE_X11Y103_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y103_SLICE_X11Y103_BO5),
.O6(CLBLM_L_X8Y103_SLICE_X11Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y103_SLICE_X11Y103_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y103_SLICE_X11Y103_AO5),
.O6(CLBLM_L_X8Y103_SLICE_X11Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c5373730453737)
  ) CLBLM_L_X8Y104_SLICE_X10Y104_DLUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_L_X8Y104_SLICE_X10Y104_DO5),
.O6(CLBLM_L_X8Y104_SLICE_X10Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hea4466cc2688aa00)
  ) CLBLM_L_X8Y104_SLICE_X10Y104_CLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(LIOB33_X0Y101_IOB_X0Y101_I),
.O5(CLBLM_L_X8Y104_SLICE_X10Y104_CO5),
.O6(CLBLM_L_X8Y104_SLICE_X10Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb8787b7747878488)
  ) CLBLM_L_X8Y104_SLICE_X10Y104_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(CLBLM_L_X10Y104_SLICE_X12Y104_AO6),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(CLBLM_L_X10Y104_SLICE_X12Y104_CO6),
.I5(CLBLM_L_X10Y104_SLICE_X12Y104_BO6),
.O5(CLBLM_L_X8Y104_SLICE_X10Y104_BO5),
.O6(CLBLM_L_X8Y104_SLICE_X10Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0bbbbbafbfffff)
  ) CLBLM_L_X8Y104_SLICE_X10Y104_ALUT (
.I0(CLBLM_L_X8Y104_SLICE_X10Y104_DO6),
.I1(CLBLM_L_X8Y102_SLICE_X10Y102_CO6),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(CLBLM_L_X8Y104_SLICE_X10Y104_CO6),
.O5(CLBLM_L_X8Y104_SLICE_X10Y104_AO5),
.O6(CLBLM_L_X8Y104_SLICE_X10Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y104_SLICE_X11Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y104_SLICE_X11Y104_DO5),
.O6(CLBLM_L_X8Y104_SLICE_X11Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y104_SLICE_X11Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y104_SLICE_X11Y104_CO5),
.O6(CLBLM_L_X8Y104_SLICE_X11Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3963c993366cc)
  ) CLBLM_L_X8Y104_SLICE_X11Y104_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(CLBLM_L_X10Y103_SLICE_X12Y103_BO6),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(CLBLM_L_X10Y104_SLICE_X12Y104_AO6),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_L_X8Y104_SLICE_X11Y104_BO5),
.O6(CLBLM_L_X8Y104_SLICE_X11Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6f06cf0cff66ffcc)
  ) CLBLM_L_X8Y104_SLICE_X11Y104_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(CLBLM_L_X10Y103_SLICE_X12Y103_BO6),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLM_L_X10Y104_SLICE_X12Y104_AO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_L_X8Y104_SLICE_X11Y104_AO5),
.O6(CLBLM_L_X8Y104_SLICE_X11Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7ddd1444ffff3ccc)
  ) CLBLM_L_X8Y105_SLICE_X10Y105_DLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(CLBLM_L_X10Y105_SLICE_X13Y105_DO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(CLBLM_L_X10Y106_SLICE_X13Y106_CO6),
.I5(RIOB33_X105Y101_IOB_X1Y102_I),
.O5(CLBLM_L_X8Y105_SLICE_X10Y105_DO5),
.O6(CLBLM_L_X8Y105_SLICE_X10Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69999666c3333ccc)
  ) CLBLM_L_X8Y105_SLICE_X10Y105_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(CLBLM_L_X10Y105_SLICE_X13Y105_DO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(CLBLM_L_X10Y106_SLICE_X13Y106_CO6),
.I5(RIOB33_X105Y101_IOB_X1Y102_I),
.O5(CLBLM_L_X8Y105_SLICE_X10Y105_CO5),
.O6(CLBLM_L_X8Y105_SLICE_X10Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb4d22dd24bd2d2d2)
  ) CLBLM_L_X8Y105_SLICE_X10Y105_BLUT (
.I0(CLBLM_L_X10Y105_SLICE_X12Y105_DO6),
.I1(CLBLM_L_X10Y106_SLICE_X13Y106_CO6),
.I2(CLBLM_L_X10Y104_SLICE_X12Y104_DO6),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_L_X8Y105_SLICE_X10Y105_BO5),
.O6(CLBLM_L_X8Y105_SLICE_X10Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff33ff33ff)
  ) CLBLM_L_X8Y105_SLICE_X10Y105_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(1'b1),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y105_SLICE_X10Y105_AO5),
.O6(CLBLM_L_X8Y105_SLICE_X10Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y105_SLICE_X11Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y105_SLICE_X11Y105_DO5),
.O6(CLBLM_L_X8Y105_SLICE_X11Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y105_SLICE_X11Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y105_SLICE_X11Y105_CO5),
.O6(CLBLM_L_X8Y105_SLICE_X11Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y105_SLICE_X11Y105_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y105_SLICE_X11Y105_BO5),
.O6(CLBLM_L_X8Y105_SLICE_X11Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y105_SLICE_X11Y105_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y105_SLICE_X11Y105_AO5),
.O6(CLBLM_L_X8Y105_SLICE_X11Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdf7c431dc734010)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_DLUT (
.I0(CLBLM_L_X10Y105_SLICE_X12Y105_DO6),
.I1(CLBLM_L_X8Y105_SLICE_X10Y105_AO5),
.I2(CLBLM_L_X10Y106_SLICE_X13Y106_CO6),
.I3(CLBLM_L_X10Y104_SLICE_X12Y104_DO6),
.I4(CLBLM_L_X8Y107_SLICE_X10Y107_AO5),
.I5(CLBLM_R_X7Y106_SLICE_X9Y106_AO6),
.O5(CLBLM_L_X8Y106_SLICE_X10Y106_DO5),
.O6(CLBLM_L_X8Y106_SLICE_X10Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9cc639c663c6c6c6)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_CLUT (
.I0(CLBLM_L_X8Y106_SLICE_X11Y106_BO6),
.I1(CLBLM_L_X8Y106_SLICE_X11Y106_CO6),
.I2(CLBLM_L_X8Y107_SLICE_X10Y107_BO6),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_L_X8Y106_SLICE_X10Y106_CO5),
.O6(CLBLM_L_X8Y106_SLICE_X10Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fb31320ffff5fa0)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_L_X10Y106_SLICE_X13Y106_DO6),
.I4(CLBLM_L_X10Y107_SLICE_X12Y107_DO6),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_L_X8Y106_SLICE_X10Y106_BO5),
.O6(CLBLM_L_X8Y106_SLICE_X10Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a55a69965aa596)
  ) CLBLM_L_X8Y106_SLICE_X10Y106_ALUT (
.I0(CLBLM_L_X8Y107_SLICE_X10Y107_AO5),
.I1(CLBLM_L_X10Y106_SLICE_X13Y106_CO6),
.I2(CLBLM_L_X8Y105_SLICE_X10Y105_AO5),
.I3(CLBLM_R_X7Y106_SLICE_X9Y106_AO6),
.I4(CLBLM_L_X10Y105_SLICE_X12Y105_DO6),
.I5(CLBLM_L_X10Y104_SLICE_X12Y104_DO6),
.O5(CLBLM_L_X8Y106_SLICE_X10Y106_AO5),
.O6(CLBLM_L_X8Y106_SLICE_X10Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hefae8a08df5d4504)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_DLUT (
.I0(CLBLM_L_X10Y105_SLICE_X12Y105_CO6),
.I1(CLBLM_L_X10Y107_SLICE_X12Y107_DO6),
.I2(CLBLM_L_X10Y106_SLICE_X13Y106_BO6),
.I3(CLBLM_L_X8Y107_SLICE_X11Y107_AO5),
.I4(CLBLM_R_X7Y104_SLICE_X8Y104_BO6),
.I5(CLBLM_R_X7Y106_SLICE_X9Y106_AO6),
.O5(CLBLM_L_X8Y106_SLICE_X11Y106_DO5),
.O6(CLBLM_L_X8Y106_SLICE_X11Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h965aa596aaaa55aa)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_CLUT (
.I0(CLBLM_L_X10Y105_SLICE_X12Y105_CO6),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(CLBLM_L_X10Y106_SLICE_X13Y106_BO6),
.I4(CLBLM_L_X10Y107_SLICE_X12Y107_DO6),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLM_L_X8Y106_SLICE_X11Y106_CO5),
.O6(CLBLM_L_X8Y106_SLICE_X11Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999c33396663ccc)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLM_L_X10Y107_SLICE_X12Y107_DO6),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(CLBLM_L_X10Y106_SLICE_X13Y106_DO6),
.O5(CLBLM_L_X8Y106_SLICE_X11Y106_BO5),
.O6(CLBLM_L_X8Y106_SLICE_X11Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h788787781ee1e11e)
  ) CLBLM_L_X8Y106_SLICE_X11Y106_ALUT (
.I0(CLBLM_L_X10Y107_SLICE_X12Y107_DO6),
.I1(CLBLM_L_X8Y107_SLICE_X11Y107_AO5),
.I2(CLBLM_R_X7Y104_SLICE_X8Y104_BO6),
.I3(CLBLM_R_X7Y106_SLICE_X9Y106_AO6),
.I4(CLBLM_L_X10Y105_SLICE_X12Y105_CO6),
.I5(CLBLM_L_X10Y106_SLICE_X13Y106_BO6),
.O5(CLBLM_L_X8Y106_SLICE_X11Y106_AO5),
.O6(CLBLM_L_X8Y106_SLICE_X11Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h965aaaaaa59655aa)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_DLUT (
.I0(CLBLM_L_X8Y106_SLICE_X11Y106_AO6),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(CLBLM_L_X8Y106_SLICE_X11Y106_BO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_L_X8Y107_SLICE_X10Y107_BO6),
.O5(CLBLM_L_X8Y107_SLICE_X10Y107_DO5),
.O6(CLBLM_L_X8Y107_SLICE_X10Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h175fffff051755ff)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_CLUT (
.I0(CLBLM_L_X8Y106_SLICE_X11Y106_AO6),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(CLBLM_L_X8Y106_SLICE_X11Y106_BO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_L_X8Y107_SLICE_X10Y107_BO6),
.O5(CLBLM_L_X8Y107_SLICE_X10Y107_CO5),
.O6(CLBLM_L_X8Y107_SLICE_X10Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7bfff3ff125a30f0)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(CLBLM_R_X11Y107_SLICE_X14Y107_BO6),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(CLBLM_L_X10Y108_SLICE_X12Y108_AO6),
.O5(CLBLM_L_X8Y107_SLICE_X10Y107_BO5),
.O6(CLBLM_L_X8Y107_SLICE_X10Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff0f0fffff)
  ) CLBLM_L_X8Y107_SLICE_X10Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y107_SLICE_X10Y107_AO5),
.O6(CLBLM_L_X8Y107_SLICE_X10Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h78871ee18778e11e)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_DLUT (
.I0(CLBLM_L_X8Y107_SLICE_X11Y107_AO6),
.I1(CLBLM_L_X10Y108_SLICE_X12Y108_AO6),
.I2(CLBLM_L_X10Y107_SLICE_X12Y107_DO6),
.I3(CLBLM_L_X8Y107_SLICE_X11Y107_AO5),
.I4(CLBLM_L_X10Y107_SLICE_X12Y107_CO6),
.I5(CLBLM_L_X10Y106_SLICE_X13Y106_BO6),
.O5(CLBLM_L_X8Y107_SLICE_X11Y107_DO5),
.O6(CLBLM_L_X8Y107_SLICE_X11Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hebff82c3c3eb0082)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_CLUT (
.I0(CLBLM_L_X8Y107_SLICE_X11Y107_AO6),
.I1(CLBLM_L_X10Y107_SLICE_X12Y107_BO6),
.I2(CLBLM_L_X8Y107_SLICE_X11Y107_AO5),
.I3(CLBLM_L_X10Y107_SLICE_X12Y107_CO6),
.I4(CLBLM_L_X8Y107_SLICE_X10Y107_AO6),
.I5(CLBLM_L_X10Y108_SLICE_X12Y108_AO6),
.O5(CLBLM_L_X8Y107_SLICE_X11Y107_CO5),
.O6(CLBLM_L_X8Y107_SLICE_X11Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c9696c3c369693c)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_BLUT (
.I0(CLBLM_L_X10Y107_SLICE_X12Y107_CO6),
.I1(CLBLM_L_X10Y107_SLICE_X12Y107_BO6),
.I2(CLBLM_L_X8Y107_SLICE_X10Y107_AO6),
.I3(CLBLM_L_X10Y108_SLICE_X12Y108_AO6),
.I4(CLBLM_L_X8Y107_SLICE_X11Y107_AO6),
.I5(CLBLM_L_X8Y107_SLICE_X11Y107_AO5),
.O5(CLBLM_L_X8Y107_SLICE_X11Y107_BO5),
.O6(CLBLM_L_X8Y107_SLICE_X11Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff00ffffff)
  ) CLBLM_L_X8Y107_SLICE_X11Y107_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(1'b1),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y107_SLICE_X11Y107_AO5),
.O6(CLBLM_L_X8Y107_SLICE_X11Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h956aa956ff0033cc)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_DLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_L_X10Y108_SLICE_X12Y108_CO6),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(CLBLM_L_X10Y108_SLICE_X12Y108_BO6),
.I4(CLBLM_L_X8Y109_SLICE_X10Y109_DO6),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_DO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hefdfae5d8a450804)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_CLUT (
.I0(CLBLM_L_X8Y107_SLICE_X11Y107_AO6),
.I1(CLBLM_R_X7Y109_SLICE_X9Y109_AO5),
.I2(CLBLM_L_X10Y108_SLICE_X12Y108_CO6),
.I3(CLBLM_L_X10Y108_SLICE_X12Y108_BO6),
.I4(CLBLM_L_X8Y109_SLICE_X10Y109_DO6),
.I5(CLBLM_R_X7Y108_SLICE_X9Y108_AO6),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_CO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7b12ff5abb22ffaa)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_BLUT (
.I0(CLBLM_L_X10Y108_SLICE_X12Y108_DO6),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_L_X8Y109_SLICE_X10Y109_DO6),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_BO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4bb4b44bd22d2dd2)
  ) CLBLM_L_X8Y108_SLICE_X10Y108_ALUT (
.I0(CLBLM_L_X8Y109_SLICE_X10Y109_DO6),
.I1(CLBLM_L_X10Y108_SLICE_X12Y108_CO6),
.I2(CLBLM_L_X8Y107_SLICE_X11Y107_AO6),
.I3(CLBLM_R_X7Y108_SLICE_X9Y108_AO6),
.I4(CLBLM_L_X10Y108_SLICE_X12Y108_BO6),
.I5(CLBLM_R_X7Y109_SLICE_X9Y109_AO5),
.O5(CLBLM_L_X8Y108_SLICE_X10Y108_AO5),
.O6(CLBLM_L_X8Y108_SLICE_X10Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_DO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_CO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_BO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y108_SLICE_X11Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y108_SLICE_X11Y108_AO5),
.O6(CLBLM_L_X8Y108_SLICE_X11Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4dcfddff8e0ceecc)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_DLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLM_L_X10Y110_SLICE_X12Y110_CO6),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_DO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a5965a995566aa)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_CLUT (
.I0(CLBLM_L_X10Y108_SLICE_X12Y108_DO6),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(CLBLM_L_X8Y109_SLICE_X10Y109_DO6),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_CO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h15403fc04015c03f)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_L_X10Y110_SLICE_X12Y110_CO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_BO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a95c03f956a3fc0)
  ) CLBLM_L_X8Y109_SLICE_X10Y109_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_L_X10Y110_SLICE_X12Y110_CO6),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.O5(CLBLM_L_X8Y109_SLICE_X10Y109_AO5),
.O6(CLBLM_L_X8Y109_SLICE_X10Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_DO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_CO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69963cc3c33c6996)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_BLUT (
.I0(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I1(CLBLM_L_X10Y110_SLICE_X12Y110_BO6),
.I2(CLBLM_L_X10Y108_SLICE_X13Y108_AO6),
.I3(CLBLM_L_X10Y107_SLICE_X12Y107_AO6),
.I4(CLBLM_L_X10Y110_SLICE_X12Y110_AO6),
.I5(CLBLM_R_X7Y110_SLICE_X9Y110_AO5),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_BO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff77777777)
  ) CLBLM_L_X8Y109_SLICE_X11Y109_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(1'b1),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y109_SLICE_X11Y109_AO5),
.O6(CLBLM_L_X8Y109_SLICE_X11Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_DO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_CO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_BO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y110_SLICE_X10Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y110_SLICE_X10Y110_AO5),
.O6(CLBLM_L_X8Y110_SLICE_X10Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ac0953f953f6ac0)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_DLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLM_L_X10Y110_SLICE_X13Y110_CO6),
.I5(CLBLM_L_X8Y111_SLICE_X11Y111_BO6),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_DO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hebc3ffeb8200c382)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_CLUT (
.I0(CLBLM_L_X8Y109_SLICE_X11Y109_AO5),
.I1(CLBLM_L_X10Y110_SLICE_X12Y110_DO6),
.I2(CLBLM_L_X10Y111_SLICE_X12Y111_AO5),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_BO6),
.I4(CLBLM_L_X8Y110_SLICE_X11Y110_DO6),
.I5(CLBLM_R_X7Y110_SLICE_X8Y110_AO5),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_CO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h93cc6cccc9663666)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_BLUT (
.I0(CLBLM_L_X8Y110_SLICE_X11Y110_DO6),
.I1(CLBLM_L_X10Y110_SLICE_X12Y110_DO6),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_L_X8Y112_SLICE_X10Y112_BO6),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_BO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h39c6c6399c63639c)
  ) CLBLM_L_X8Y110_SLICE_X11Y110_ALUT (
.I0(CLBLM_L_X8Y110_SLICE_X11Y110_DO6),
.I1(CLBLM_L_X10Y110_SLICE_X12Y110_DO6),
.I2(CLBLM_L_X8Y109_SLICE_X11Y109_AO5),
.I3(CLBLM_R_X7Y110_SLICE_X8Y110_AO5),
.I4(CLBLM_L_X10Y111_SLICE_X12Y111_AO5),
.I5(CLBLM_L_X8Y112_SLICE_X10Y112_BO6),
.O5(CLBLM_L_X8Y110_SLICE_X11Y110_AO5),
.O6(CLBLM_L_X8Y110_SLICE_X11Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h69969966c33c33cc)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_DLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_L_X8Y112_SLICE_X10Y112_BO6),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(CLBLM_L_X10Y111_SLICE_X12Y111_BO6),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_DO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffccff33ce083b02)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_CLUT (
.I0(CLBLM_L_X8Y111_SLICE_X10Y111_AO6),
.I1(CLBLM_L_X8Y112_SLICE_X11Y112_AO5),
.I2(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I3(CLBLM_L_X8Y111_SLICE_X10Y111_AO5),
.I4(CLBLM_R_X7Y112_SLICE_X9Y112_BO6),
.I5(CLBLM_R_X7Y111_SLICE_X9Y111_AO6),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_CO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a965aa5a569a55a)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_BLUT (
.I0(CLBLM_L_X8Y112_SLICE_X11Y112_AO5),
.I1(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_BO6),
.I3(CLBLM_R_X7Y111_SLICE_X9Y111_AO6),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_AO6),
.I5(CLBLM_L_X8Y111_SLICE_X10Y111_AO5),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_BO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555ffff5f5f5f5f)
  ) CLBLM_L_X8Y111_SLICE_X10Y111_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(1'b1),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(1'b1),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLM_L_X8Y111_SLICE_X10Y111_AO5),
.O6(CLBLM_L_X8Y111_SLICE_X10Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6f06ff66cf0cffcc)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_DLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_L_X10Y111_SLICE_X12Y111_BO6),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_BO6),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_DO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h96cc993366cc96cc)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_L_X10Y110_SLICE_X12Y110_CO6),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(CLBLM_L_X8Y111_SLICE_X11Y111_DO6),
.I5(CLBLM_L_X10Y111_SLICE_X12Y111_CO6),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_CO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hef8a8aefee8888ee)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_BLUT (
.I0(CLBLL_L_X4Y111_SLICE_X5Y111_AO5),
.I1(CLBLM_L_X8Y112_SLICE_X11Y112_CO6),
.I2(CLBLM_R_X7Y112_SLICE_X9Y112_BO6),
.I3(CLBLM_L_X10Y109_SLICE_X12Y109_BO6),
.I4(CLBLM_R_X11Y110_SLICE_X14Y110_AO5),
.I5(CLBLM_L_X8Y112_SLICE_X11Y112_AO5),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_BO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h39c6c6399c63639c)
  ) CLBLM_L_X8Y111_SLICE_X11Y111_ALUT (
.I0(CLBLM_L_X8Y112_SLICE_X11Y112_DO6),
.I1(CLBLM_L_X10Y110_SLICE_X13Y110_BO6),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_CO6),
.I3(CLBLM_L_X8Y111_SLICE_X11Y111_BO6),
.I4(CLBLM_L_X10Y111_SLICE_X12Y111_AO6),
.I5(CLBLM_R_X7Y112_SLICE_X9Y112_AO5),
.O5(CLBLM_L_X8Y111_SLICE_X11Y111_AO5),
.O6(CLBLM_L_X8Y111_SLICE_X11Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_DO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_CO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h71f3d4fcd4fcd4fc)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLM_L_X8Y112_SLICE_X11Y112_BO6),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_CO6),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_BO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3963c963c963c)
  ) CLBLM_L_X8Y112_SLICE_X10Y112_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLM_L_X8Y112_SLICE_X11Y112_BO6),
.I2(CLBLM_L_X8Y111_SLICE_X10Y111_CO6),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_L_X8Y112_SLICE_X10Y112_AO5),
.O6(CLBLM_L_X8Y112_SLICE_X10Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4b5ab4a5b4a54b5a)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_DLUT (
.I0(CLBLM_L_X8Y112_SLICE_X11Y112_CO6),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_BO6),
.I2(CLBLM_R_X11Y110_SLICE_X14Y110_AO5),
.I3(CLBLM_L_X8Y112_SLICE_X11Y112_AO5),
.I4(CLBLL_L_X4Y111_SLICE_X5Y111_AO5),
.I5(CLBLM_L_X10Y109_SLICE_X12Y109_BO6),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_DO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h080c783c0000cc00)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_CLUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_CO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ccccccc9663666)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_BLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_BO6),
.I1(CLBLM_L_X10Y109_SLICE_X12Y109_BO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(CLBLM_L_X8Y112_SLICE_X11Y112_CO6),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_BO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff05550fff0fff)
  ) CLBLM_L_X8Y112_SLICE_X11Y112_ALUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_BO6),
.I1(1'b1),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(CLBLM_L_X8Y112_SLICE_X11Y112_CO6),
.I5(1'b1),
.O5(CLBLM_L_X8Y112_SLICE_X11Y112_AO5),
.O6(CLBLM_L_X8Y112_SLICE_X11Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he14b78d269c35af0)
  ) CLBLM_L_X10Y101_SLICE_X12Y101_DLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(CLBLM_L_X10Y103_SLICE_X13Y103_AO5),
.I2(CLBLM_L_X8Y102_SLICE_X11Y102_CO6),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(CLBLM_L_X8Y102_SLICE_X11Y102_AO5),
.I5(RIOB33_X105Y107_IOB_X1Y107_I),
.O5(CLBLM_L_X10Y101_SLICE_X12Y101_DO5),
.O6(CLBLM_L_X10Y101_SLICE_X12Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f07f770ff777700)
  ) CLBLM_L_X10Y101_SLICE_X12Y101_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLM_R_X11Y103_SLICE_X14Y103_AO6),
.I4(CLBLM_L_X10Y101_SLICE_X12Y101_DO6),
.I5(RIOB33_X105Y107_IOB_X1Y107_I),
.O5(CLBLM_L_X10Y101_SLICE_X12Y101_CO5),
.O6(CLBLM_L_X10Y101_SLICE_X12Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f15bf2abf2abf2a)
  ) CLBLM_L_X10Y101_SLICE_X12Y101_BLUT (
.I0(CLBLM_L_X8Y102_SLICE_X11Y102_CO6),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLM_L_X10Y103_SLICE_X13Y103_BO6),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(RIOB33_X105Y107_IOB_X1Y108_I),
.O5(CLBLM_L_X10Y101_SLICE_X12Y101_BO5),
.O6(CLBLM_L_X10Y101_SLICE_X12Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a95956a956a956a)
  ) CLBLM_L_X10Y101_SLICE_X12Y101_ALUT (
.I0(CLBLM_L_X8Y102_SLICE_X11Y102_CO6),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLM_L_X10Y103_SLICE_X13Y103_BO6),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(RIOB33_X105Y107_IOB_X1Y108_I),
.O5(CLBLM_L_X10Y101_SLICE_X12Y101_AO5),
.O6(CLBLM_L_X10Y101_SLICE_X12Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y101_SLICE_X13Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y101_SLICE_X13Y101_DO5),
.O6(CLBLM_L_X10Y101_SLICE_X13Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y101_SLICE_X13Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y101_SLICE_X13Y101_CO5),
.O6(CLBLM_L_X10Y101_SLICE_X13Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h226602c600a000a0)
  ) CLBLM_L_X10Y101_SLICE_X13Y101_BLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(RIOB33_X105Y107_IOB_X1Y108_I),
.O5(CLBLM_L_X10Y101_SLICE_X13Y101_BO5),
.O6(CLBLM_L_X10Y101_SLICE_X13Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h242e04ae6a60ca60)
  ) CLBLM_L_X10Y101_SLICE_X13Y101_ALUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(RIOB33_X105Y107_IOB_X1Y108_I),
.O5(CLBLM_L_X10Y101_SLICE_X13Y101_AO5),
.O6(CLBLM_L_X10Y101_SLICE_X13Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8e71f3f3718e0c0c)
  ) CLBLM_L_X10Y102_SLICE_X12Y102_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y101_SLICE_X12Y101_AO6),
.I2(CLBLM_R_X11Y103_SLICE_X14Y103_AO6),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(CLBLM_L_X10Y102_SLICE_X12Y102_BO6),
.O5(CLBLM_L_X10Y102_SLICE_X12Y102_DO5),
.O6(CLBLM_L_X10Y102_SLICE_X12Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfab2b2a0f5717150)
  ) CLBLM_L_X10Y102_SLICE_X12Y102_CLUT (
.I0(CLBLM_L_X8Y102_SLICE_X10Y102_AO6),
.I1(CLBLM_L_X10Y101_SLICE_X12Y101_AO6),
.I2(CLBLM_L_X10Y102_SLICE_X13Y102_AO6),
.I3(CLBLM_L_X10Y102_SLICE_X13Y102_BO6),
.I4(CLBLM_R_X11Y103_SLICE_X14Y103_AO6),
.I5(CLBLM_L_X10Y102_SLICE_X12Y102_BO6),
.O5(CLBLM_L_X10Y102_SLICE_X12Y102_CO5),
.O6(CLBLM_L_X10Y102_SLICE_X12Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a9556a9956aa956)
  ) CLBLM_L_X10Y102_SLICE_X12Y102_BLUT (
.I0(CLBLM_L_X8Y103_SLICE_X10Y103_CO6),
.I1(CLBLM_L_X10Y103_SLICE_X13Y103_BO6),
.I2(CLBLM_L_X10Y102_SLICE_X13Y102_CO6),
.I3(CLBLM_R_X7Y102_SLICE_X9Y102_AO6),
.I4(CLBLM_R_X7Y102_SLICE_X9Y102_BO6),
.I5(CLBLL_L_X4Y103_SLICE_X4Y103_AO6),
.O5(CLBLM_L_X10Y102_SLICE_X12Y102_BO5),
.O6(CLBLM_L_X10Y102_SLICE_X12Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h788787781ee1e11e)
  ) CLBLM_L_X10Y102_SLICE_X12Y102_ALUT (
.I0(CLBLM_R_X11Y103_SLICE_X14Y103_AO6),
.I1(CLBLM_L_X10Y102_SLICE_X13Y102_BO6),
.I2(CLBLM_L_X10Y102_SLICE_X13Y102_AO6),
.I3(CLBLM_L_X10Y102_SLICE_X12Y102_BO6),
.I4(CLBLM_L_X8Y102_SLICE_X10Y102_AO6),
.I5(CLBLM_L_X10Y101_SLICE_X12Y101_AO6),
.O5(CLBLM_L_X10Y102_SLICE_X12Y102_AO5),
.O6(CLBLM_L_X10Y102_SLICE_X12Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6966996996996696)
  ) CLBLM_L_X10Y102_SLICE_X13Y102_DLUT (
.I0(CLBLM_L_X10Y102_SLICE_X13Y102_CO6),
.I1(CLBLM_R_X7Y102_SLICE_X9Y102_BO6),
.I2(CLBLM_R_X11Y104_SLICE_X14Y104_DO6),
.I3(CLBLM_L_X10Y103_SLICE_X13Y103_DO6),
.I4(CLBLM_L_X10Y102_SLICE_X13Y102_BO5),
.I5(CLBLM_L_X10Y103_SLICE_X13Y103_BO6),
.O5(CLBLM_L_X10Y102_SLICE_X13Y102_DO5),
.O6(CLBLM_L_X10Y102_SLICE_X13Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff77777777)
  ) CLBLM_L_X10Y102_SLICE_X13Y102_CLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(1'b1),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y102_SLICE_X13Y102_CO5),
.O6(CLBLM_L_X10Y102_SLICE_X13Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff5f5f5f5f)
  ) CLBLM_L_X10Y102_SLICE_X13Y102_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(1'b1),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y102_SLICE_X13Y102_BO5),
.O6(CLBLM_L_X10Y102_SLICE_X13Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f77777777)
  ) CLBLM_L_X10Y102_SLICE_X13Y102_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y102_SLICE_X13Y102_AO5),
.O6(CLBLM_L_X10Y102_SLICE_X13Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y103_SLICE_X12Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y103_SLICE_X12Y103_DO5),
.O6(CLBLM_L_X10Y103_SLICE_X12Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69969696c33c3c3c)
  ) CLBLM_L_X10Y103_SLICE_X12Y103_CLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(CLBLM_L_X10Y101_SLICE_X12Y101_DO6),
.I2(CLBLM_R_X11Y103_SLICE_X14Y103_AO6),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_L_X10Y103_SLICE_X12Y103_CO5),
.O6(CLBLM_L_X10Y103_SLICE_X12Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha6956a956aa66a6a)
  ) CLBLM_L_X10Y103_SLICE_X12Y103_BLUT (
.I0(CLBLM_L_X10Y102_SLICE_X12Y102_DO6),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X11Y103_SLICE_X14Y103_BO6),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(CLBLM_L_X10Y103_SLICE_X12Y103_CO6),
.O5(CLBLM_L_X10Y103_SLICE_X12Y103_BO5),
.O6(CLBLM_L_X10Y103_SLICE_X12Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a00ff6aff6aff6a)
  ) CLBLM_L_X10Y103_SLICE_X12Y103_ALUT (
.I0(CLBLM_L_X10Y102_SLICE_X12Y102_DO6),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y104_SLICE_X13Y104_AO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_L_X10Y103_SLICE_X12Y103_AO5),
.O6(CLBLM_L_X10Y103_SLICE_X12Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699996636c9c936)
  ) CLBLM_L_X10Y103_SLICE_X13Y103_DLUT (
.I0(CLBLM_L_X10Y101_SLICE_X13Y101_BO6),
.I1(CLBLM_R_X5Y101_SLICE_X7Y101_AO6),
.I2(CLBLL_L_X4Y103_SLICE_X4Y103_BO6),
.I3(CLBLM_L_X10Y102_SLICE_X13Y102_CO5),
.I4(CLBLM_L_X10Y101_SLICE_X13Y101_AO6),
.I5(CLBLM_L_X12Y104_SLICE_X16Y104_BO6),
.O5(CLBLM_L_X10Y103_SLICE_X13Y103_DO5),
.O6(CLBLM_L_X10Y103_SLICE_X13Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ffff000e3131cec)
  ) CLBLM_L_X10Y103_SLICE_X13Y103_CLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(CLBLM_L_X12Y104_SLICE_X16Y104_BO6),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(CLBLM_L_X10Y101_SLICE_X13Y101_AO6),
.I5(CLBLM_L_X10Y101_SLICE_X13Y101_BO6),
.O5(CLBLM_L_X10Y103_SLICE_X13Y103_CO5),
.O6(CLBLM_L_X10Y103_SLICE_X13Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaf5b271faf5a050)
  ) CLBLM_L_X10Y103_SLICE_X13Y103_BLUT (
.I0(CLBLM_L_X10Y101_SLICE_X13Y101_AO6),
.I1(CLBLM_L_X12Y104_SLICE_X16Y104_BO6),
.I2(CLBLM_L_X10Y102_SLICE_X13Y102_CO5),
.I3(CLBLM_R_X5Y101_SLICE_X7Y101_AO6),
.I4(CLBLM_L_X10Y101_SLICE_X13Y101_BO6),
.I5(CLBLL_L_X4Y103_SLICE_X4Y103_BO6),
.O5(CLBLM_L_X10Y103_SLICE_X13Y103_BO5),
.O6(CLBLM_L_X10Y103_SLICE_X13Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3c33333ff03ff33)
  ) CLBLM_L_X10Y103_SLICE_X13Y103_ALUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y104_SLICE_X16Y104_BO6),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(CLBLM_L_X10Y101_SLICE_X13Y101_BO6),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y103_SLICE_X13Y103_AO5),
.O6(CLBLM_L_X10Y103_SLICE_X13Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6696969999696966)
  ) CLBLM_L_X10Y104_SLICE_X12Y104_DLUT (
.I0(CLBLM_L_X10Y102_SLICE_X12Y102_AO6),
.I1(CLBLM_L_X10Y104_SLICE_X13Y104_AO6),
.I2(CLBLM_L_X10Y104_SLICE_X13Y104_BO6),
.I3(CLBLM_R_X11Y105_SLICE_X14Y105_BO6),
.I4(CLBLM_L_X8Y105_SLICE_X10Y105_AO6),
.I5(CLBLM_L_X10Y105_SLICE_X12Y105_BO6),
.O5(CLBLM_L_X10Y104_SLICE_X12Y104_DO5),
.O6(CLBLM_L_X10Y104_SLICE_X12Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3963c993366cc)
  ) CLBLM_L_X10Y104_SLICE_X12Y104_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_L_X10Y104_SLICE_X13Y104_AO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X10Y102_SLICE_X12Y102_DO6),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_L_X10Y104_SLICE_X12Y104_CO5),
.O6(CLBLM_L_X10Y104_SLICE_X12Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999666996669996)
  ) CLBLM_L_X10Y104_SLICE_X12Y104_BLUT (
.I0(CLBLM_L_X10Y105_SLICE_X12Y105_AO5),
.I1(CLBLM_L_X8Y102_SLICE_X11Y102_BO6),
.I2(CLBLM_L_X10Y104_SLICE_X13Y104_AO6),
.I3(CLBLM_L_X10Y105_SLICE_X12Y105_BO6),
.I4(CLBLM_L_X10Y102_SLICE_X12Y102_AO6),
.I5(CLBLM_L_X10Y102_SLICE_X12Y102_CO6),
.O5(CLBLM_L_X10Y104_SLICE_X12Y104_BO5),
.O6(CLBLM_L_X10Y104_SLICE_X12Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6affffff006a6a6a)
  ) CLBLM_L_X10Y104_SLICE_X12Y104_ALUT (
.I0(CLBLM_L_X10Y104_SLICE_X13Y104_CO6),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_R_X11Y105_SLICE_X14Y105_BO6),
.O5(CLBLM_L_X10Y104_SLICE_X12Y104_AO5),
.O6(CLBLM_L_X10Y104_SLICE_X12Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3963c3c69c396)
  ) CLBLM_L_X10Y104_SLICE_X13Y104_DLUT (
.I0(CLBLM_L_X10Y106_SLICE_X12Y106_CO6),
.I1(CLBLM_R_X11Y104_SLICE_X14Y104_DO6),
.I2(CLBLM_L_X10Y103_SLICE_X13Y103_DO6),
.I3(CLBLM_L_X10Y105_SLICE_X13Y105_AO5),
.I4(CLBLM_L_X10Y102_SLICE_X13Y102_BO5),
.I5(CLBLM_R_X11Y104_SLICE_X14Y104_CO6),
.O5(CLBLM_L_X10Y104_SLICE_X13Y104_DO5),
.O6(CLBLM_L_X10Y104_SLICE_X13Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h93ffc9556c0036aa)
  ) CLBLM_L_X10Y104_SLICE_X13Y104_CLUT (
.I0(CLBLM_R_X11Y104_SLICE_X14Y104_BO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(CLBLM_R_X11Y104_SLICE_X15Y104_CO6),
.I5(CLBLM_L_X10Y102_SLICE_X13Y102_DO6),
.O5(CLBLM_L_X10Y104_SLICE_X13Y104_CO5),
.O6(CLBLM_L_X10Y104_SLICE_X13Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996669999666996)
  ) CLBLM_L_X10Y104_SLICE_X13Y104_BLUT (
.I0(CLBLM_L_X10Y105_SLICE_X12Y105_BO5),
.I1(CLBLM_L_X10Y102_SLICE_X13Y102_BO6),
.I2(CLBLM_L_X10Y105_SLICE_X13Y105_AO6),
.I3(CLBLM_L_X10Y102_SLICE_X13Y102_DO6),
.I4(CLBLM_R_X11Y104_SLICE_X14Y104_BO6),
.I5(CLBLM_R_X11Y104_SLICE_X15Y104_CO6),
.O5(CLBLM_L_X10Y104_SLICE_X13Y104_BO5),
.O6(CLBLM_L_X10Y104_SLICE_X13Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he88efaafa00ae88e)
  ) CLBLM_L_X10Y104_SLICE_X13Y104_ALUT (
.I0(CLBLM_L_X10Y105_SLICE_X12Y105_BO5),
.I1(CLBLM_L_X10Y105_SLICE_X13Y105_AO6),
.I2(CLBLM_L_X10Y102_SLICE_X13Y102_DO6),
.I3(CLBLM_L_X10Y102_SLICE_X13Y102_BO6),
.I4(CLBLM_R_X11Y104_SLICE_X14Y104_BO6),
.I5(CLBLM_R_X11Y104_SLICE_X15Y104_CO6),
.O5(CLBLM_L_X10Y104_SLICE_X13Y104_AO5),
.O6(CLBLM_L_X10Y104_SLICE_X13Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93936c936c936c)
  ) CLBLM_L_X10Y105_SLICE_X12Y105_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_L_X10Y104_SLICE_X13Y104_CO6),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(CLBLM_R_X11Y105_SLICE_X14Y105_BO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_L_X10Y105_SLICE_X12Y105_DO5),
.O6(CLBLM_L_X10Y105_SLICE_X12Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h639cc6399c6339c6)
  ) CLBLM_L_X10Y105_SLICE_X12Y105_CLUT (
.I0(CLBLM_L_X10Y105_SLICE_X12Y105_AO6),
.I1(CLBLM_L_X8Y105_SLICE_X10Y105_AO6),
.I2(CLBLM_R_X11Y105_SLICE_X14Y105_CO6),
.I3(CLBLM_L_X10Y104_SLICE_X13Y104_BO6),
.I4(CLBLM_R_X11Y107_SLICE_X15Y107_BO6),
.I5(CLBLM_R_X11Y105_SLICE_X14Y105_BO6),
.O5(CLBLM_L_X10Y105_SLICE_X12Y105_CO5),
.O6(CLBLM_L_X10Y105_SLICE_X12Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffff0f0fffff)
  ) CLBLM_L_X10Y105_SLICE_X12Y105_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(1'b1),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y105_SLICE_X12Y105_BO5),
.O6(CLBLM_L_X10Y105_SLICE_X12Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f33ff33ff)
  ) CLBLM_L_X10Y105_SLICE_X12Y105_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y105_SLICE_X12Y105_AO5),
.O6(CLBLM_L_X10Y105_SLICE_X12Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc69c6c366696cc3c)
  ) CLBLM_L_X10Y105_SLICE_X13Y105_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_L_X10Y104_SLICE_X13Y104_CO6),
.I2(CLBLM_R_X11Y104_SLICE_X14Y104_AO6),
.I3(CLBLM_L_X10Y105_SLICE_X13Y105_CO6),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_L_X10Y105_SLICE_X13Y105_DO5),
.O6(CLBLM_L_X10Y105_SLICE_X13Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h71d4f550f3fcfff0)
  ) CLBLM_L_X10Y105_SLICE_X13Y105_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(CLBLM_R_X11Y106_SLICE_X15Y106_DO6),
.I3(CLBLM_R_X11Y105_SLICE_X15Y105_DO6),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_L_X10Y105_SLICE_X13Y105_CO5),
.O6(CLBLM_L_X10Y105_SLICE_X13Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6ca0935f935f6ca0)
  ) CLBLM_L_X10Y105_SLICE_X13Y105_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(CLBLM_R_X11Y106_SLICE_X15Y106_DO6),
.I5(CLBLM_R_X11Y105_SLICE_X15Y105_DO6),
.O5(CLBLM_L_X10Y105_SLICE_X13Y105_BO5),
.O6(CLBLM_L_X10Y105_SLICE_X13Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff0f0fffff)
  ) CLBLM_L_X10Y105_SLICE_X13Y105_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y105_SLICE_X13Y105_AO5),
.O6(CLBLM_L_X10Y105_SLICE_X13Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5aa5a596a5695a)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_DLUT (
.I0(CLBLM_L_X10Y106_SLICE_X12Y106_AO6),
.I1(CLBLM_R_X11Y106_SLICE_X15Y106_BO6),
.I2(CLBLM_R_X11Y105_SLICE_X15Y105_AO6),
.I3(CLBLM_L_X10Y106_SLICE_X12Y106_AO5),
.I4(CLBLM_R_X11Y104_SLICE_X15Y104_AO6),
.I5(CLBLM_R_X11Y105_SLICE_X15Y105_BO6),
.O5(CLBLM_L_X10Y106_SLICE_X12Y106_DO5),
.O6(CLBLM_L_X10Y106_SLICE_X12Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafaafafb2a02b0a)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_CLUT (
.I0(CLBLM_L_X10Y106_SLICE_X12Y106_AO6),
.I1(CLBLM_R_X11Y106_SLICE_X15Y106_BO6),
.I2(CLBLM_R_X11Y105_SLICE_X15Y105_AO6),
.I3(CLBLM_L_X10Y106_SLICE_X12Y106_AO5),
.I4(CLBLM_R_X11Y104_SLICE_X15Y104_AO6),
.I5(CLBLM_R_X11Y105_SLICE_X15Y105_BO6),
.O5(CLBLM_L_X10Y106_SLICE_X12Y106_CO5),
.O6(CLBLM_L_X10Y106_SLICE_X12Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h155a25aac050f0a0)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O5(CLBLM_L_X10Y106_SLICE_X12Y106_BO5),
.O6(CLBLM_L_X10Y106_SLICE_X12Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff5f5f5f5f)
  ) CLBLM_L_X10Y106_SLICE_X12Y106_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(1'b1),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(1'b1),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y106_SLICE_X12Y106_AO5),
.O6(CLBLM_L_X10Y106_SLICE_X12Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc6aa395563ff9c00)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_DLUT (
.I0(CLBLM_R_X11Y106_SLICE_X14Y106_BO6),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(CLBLM_R_X11Y105_SLICE_X14Y105_DO6),
.I5(CLBLM_L_X10Y105_SLICE_X13Y105_BO6),
.O5(CLBLM_L_X10Y106_SLICE_X13Y106_DO5),
.O6(CLBLM_L_X10Y106_SLICE_X13Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h032bbbbb2b3fffff)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_CLUT (
.I0(CLBLM_R_X11Y106_SLICE_X14Y106_BO6),
.I1(CLBLM_R_X11Y105_SLICE_X14Y105_CO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(CLBLM_L_X10Y105_SLICE_X13Y105_BO6),
.O5(CLBLM_L_X10Y106_SLICE_X13Y106_CO5),
.O6(CLBLM_L_X10Y106_SLICE_X13Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h96cc993366cc96cc)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLM_R_X11Y105_SLICE_X14Y105_CO6),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(CLBLM_R_X11Y106_SLICE_X14Y106_BO6),
.I5(CLBLM_L_X10Y105_SLICE_X13Y105_BO6),
.O5(CLBLM_L_X10Y106_SLICE_X13Y106_BO5),
.O6(CLBLM_L_X10Y106_SLICE_X13Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4bd2b42db42d4bd2)
  ) CLBLM_L_X10Y106_SLICE_X13Y106_ALUT (
.I0(CLBLM_L_X10Y107_SLICE_X13Y107_AO5),
.I1(CLBLM_L_X10Y106_SLICE_X12Y106_DO6),
.I2(CLBLM_L_X10Y106_SLICE_X12Y106_CO6),
.I3(CLBLM_L_X10Y107_SLICE_X13Y107_CO6),
.I4(CLBLM_L_X10Y105_SLICE_X13Y105_AO5),
.I5(CLBLM_R_X11Y104_SLICE_X14Y104_CO6),
.O5(CLBLM_L_X10Y106_SLICE_X13Y106_AO5),
.O6(CLBLM_L_X10Y106_SLICE_X13Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2b8e8e8ebbeeeeee)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_DLUT (
.I0(CLBLM_L_X10Y108_SLICE_X13Y108_DO6),
.I1(CLBLM_R_X11Y107_SLICE_X15Y107_CO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_L_X10Y107_SLICE_X12Y107_DO5),
.O6(CLBLM_L_X10Y107_SLICE_X12Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996969699666666)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_CLUT (
.I0(CLBLM_L_X10Y108_SLICE_X13Y108_DO6),
.I1(CLBLM_R_X11Y107_SLICE_X15Y107_CO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_L_X10Y107_SLICE_X12Y107_CO5),
.O6(CLBLM_L_X10Y107_SLICE_X12Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa596699669a55a)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_BLUT (
.I0(CLBLM_R_X11Y105_SLICE_X14Y105_CO6),
.I1(CLBLM_R_X11Y107_SLICE_X15Y107_DO6),
.I2(CLBLM_L_X10Y105_SLICE_X12Y105_AO6),
.I3(CLBLM_R_X11Y107_SLICE_X15Y107_BO6),
.I4(CLBLM_L_X10Y108_SLICE_X13Y108_DO6),
.I5(CLBLM_L_X10Y107_SLICE_X12Y107_AO5),
.O5(CLBLM_L_X10Y107_SLICE_X12Y107_BO5),
.O6(CLBLM_L_X10Y107_SLICE_X12Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff5f5f5f5f)
  ) CLBLM_L_X10Y107_SLICE_X12Y107_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(1'b1),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y107_SLICE_X12Y107_AO5),
.O6(CLBLM_L_X10Y107_SLICE_X12Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6699669999669669)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_DLUT (
.I0(CLBLM_L_X10Y107_SLICE_X13Y107_AO6),
.I1(CLBLM_L_X10Y106_SLICE_X12Y106_AO5),
.I2(CLBLM_R_X11Y106_SLICE_X14Y106_AO6),
.I3(CLBLM_R_X11Y106_SLICE_X15Y106_BO6),
.I4(CLBLM_R_X5Y109_SLICE_X7Y109_AO5),
.I5(CLBLM_L_X10Y107_SLICE_X13Y107_BO6),
.O5(CLBLM_L_X10Y107_SLICE_X13Y107_DO5),
.O6(CLBLM_L_X10Y107_SLICE_X13Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'heebbeebb88228e2b)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_CLUT (
.I0(CLBLM_L_X10Y107_SLICE_X13Y107_AO6),
.I1(CLBLM_L_X10Y106_SLICE_X12Y106_AO5),
.I2(CLBLM_R_X11Y106_SLICE_X14Y106_AO6),
.I3(CLBLM_R_X11Y106_SLICE_X15Y106_BO6),
.I4(CLBLM_R_X5Y109_SLICE_X7Y109_AO5),
.I5(CLBLM_L_X10Y107_SLICE_X13Y107_BO6),
.O5(CLBLM_L_X10Y107_SLICE_X13Y107_CO5),
.O6(CLBLM_L_X10Y107_SLICE_X13Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h406a505a00f00000)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_BLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_L_X10Y107_SLICE_X13Y107_BO5),
.O6(CLBLM_L_X10Y107_SLICE_X13Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff00ffffff)
  ) CLBLM_L_X10Y107_SLICE_X13Y107_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(1'b1),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y107_SLICE_X13Y107_AO5),
.O6(CLBLM_L_X10Y107_SLICE_X13Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd52a7f80ad5207f8)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_R_X11Y108_SLICE_X14Y108_CO6),
.I3(CLBLM_R_X11Y108_SLICE_X14Y108_BO6),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(CLBLM_L_X10Y111_SLICE_X13Y111_AO6),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_DO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93a05f936c5fa0)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLM_R_X11Y108_SLICE_X14Y108_BO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_L_X10Y110_SLICE_X12Y110_BO6),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_CO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6696969999696966)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_BLUT (
.I0(CLBLM_R_X11Y107_SLICE_X15Y107_DO6),
.I1(CLBLM_L_X10Y108_SLICE_X13Y108_DO6),
.I2(CLBLM_L_X10Y108_SLICE_X13Y108_AO6),
.I3(CLBLM_L_X10Y110_SLICE_X12Y110_BO6),
.I4(CLBLM_L_X10Y107_SLICE_X12Y107_AO6),
.I5(CLBLM_L_X10Y107_SLICE_X12Y107_AO5),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_BO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f13ff5fb320ffa0)
  ) CLBLM_L_X10Y108_SLICE_X12Y108_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_L_X10Y110_SLICE_X12Y110_BO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_R_X11Y108_SLICE_X14Y108_BO6),
.O5(CLBLM_L_X10Y108_SLICE_X12Y108_AO5),
.O6(CLBLM_L_X10Y108_SLICE_X12Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hef8c8cefce0808ce)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_DLUT (
.I0(CLBLM_L_X8Y109_SLICE_X11Y109_AO6),
.I1(CLBLM_L_X10Y109_SLICE_X12Y109_AO5),
.I2(CLBLM_R_X11Y108_SLICE_X15Y108_CO6),
.I3(CLBLM_L_X10Y108_SLICE_X13Y108_CO6),
.I4(CLBLM_R_X11Y107_SLICE_X15Y107_AO6),
.I5(CLBLM_R_X11Y109_SLICE_X14Y109_BO6),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_DO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h65a69a599a5965a6)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_CLUT (
.I0(CLBLM_L_X10Y107_SLICE_X13Y107_AO5),
.I1(CLBLM_R_X11Y107_SLICE_X15Y107_AO5),
.I2(CLBLM_L_X10Y107_SLICE_X13Y107_DO6),
.I3(CLBLM_L_X10Y109_SLICE_X13Y109_DO6),
.I4(CLBLM_L_X10Y106_SLICE_X12Y106_DO6),
.I5(CLBLM_L_X10Y107_SLICE_X13Y107_CO6),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_CO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h280aa02882a00a82)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_BLUT (
.I0(CLBLM_L_X10Y109_SLICE_X12Y109_AO5),
.I1(CLBLM_R_X11Y109_SLICE_X14Y109_BO6),
.I2(CLBLM_R_X11Y107_SLICE_X15Y107_AO6),
.I3(CLBLM_R_X11Y108_SLICE_X15Y108_CO6),
.I4(CLBLM_L_X8Y109_SLICE_X11Y109_AO6),
.I5(CLBLM_L_X10Y108_SLICE_X13Y108_CO6),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_BO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h695aa56996a55a96)
  ) CLBLM_L_X10Y108_SLICE_X13Y108_ALUT (
.I0(CLBLM_L_X10Y109_SLICE_X12Y109_AO5),
.I1(CLBLM_R_X11Y109_SLICE_X14Y109_BO6),
.I2(CLBLM_R_X11Y107_SLICE_X15Y107_AO6),
.I3(CLBLM_R_X11Y108_SLICE_X15Y108_CO6),
.I4(CLBLM_L_X8Y109_SLICE_X11Y109_AO6),
.I5(CLBLM_L_X10Y108_SLICE_X13Y108_CO6),
.O5(CLBLM_L_X10Y108_SLICE_X13Y108_AO5),
.O6(CLBLM_L_X10Y108_SLICE_X13Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887878787787878)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_DLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(CLBLM_L_X10Y110_SLICE_X13Y110_DO6),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(CLBLM_R_X11Y109_SLICE_X14Y109_CO6),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_DO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4bb4d22db44b2dd2)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_CLUT (
.I0(CLBLM_L_X10Y109_SLICE_X12Y109_AO6),
.I1(CLBLM_L_X10Y109_SLICE_X13Y109_CO6),
.I2(CLBLM_L_X10Y109_SLICE_X13Y109_DO6),
.I3(CLBLM_R_X11Y107_SLICE_X15Y107_AO5),
.I4(CLBLM_L_X10Y110_SLICE_X13Y110_DO6),
.I5(CLBLM_L_X10Y107_SLICE_X13Y107_DO6),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_CO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h12665a66de001e00)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_BO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h777777775f5f5f5f)
  ) CLBLM_L_X10Y109_SLICE_X12Y109_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y109_SLICE_X12Y109_AO5),
.O6(CLBLM_L_X10Y109_SLICE_X12Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfef458addee4488)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_DLUT (
.I0(CLBLM_R_X11Y106_SLICE_X14Y106_AO6),
.I1(CLBLM_R_X11Y108_SLICE_X15Y108_AO6),
.I2(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I3(CLBLM_R_X5Y109_SLICE_X7Y109_AO5),
.I4(CLBLM_L_X10Y109_SLICE_X13Y109_BO5),
.I5(CLBLM_L_X10Y109_SLICE_X13Y109_BO6),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_DO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9a65659a99666699)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_CLUT (
.I0(CLBLM_R_X11Y106_SLICE_X14Y106_AO6),
.I1(CLBLM_R_X11Y108_SLICE_X15Y108_AO6),
.I2(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I3(CLBLM_R_X5Y109_SLICE_X7Y109_AO5),
.I4(CLBLM_L_X10Y109_SLICE_X13Y109_BO5),
.I5(CLBLM_L_X10Y109_SLICE_X13Y109_BO6),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_CO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff00ffffff)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(1'b1),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_BO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff0fff0fff)
  ) CLBLM_L_X10Y109_SLICE_X13Y109_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y109_SLICE_X13Y109_AO5),
.O6(CLBLM_L_X10Y109_SLICE_X13Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h639c9c63c63939c6)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_DLUT (
.I0(CLBLM_L_X8Y111_SLICE_X11Y111_BO6),
.I1(CLBLM_L_X10Y109_SLICE_X13Y109_CO6),
.I2(CLBLM_L_X10Y110_SLICE_X13Y110_BO6),
.I3(CLBLM_L_X10Y110_SLICE_X13Y110_DO6),
.I4(CLBLM_L_X10Y109_SLICE_X12Y109_AO6),
.I5(CLBLM_L_X10Y111_SLICE_X12Y111_AO6),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_DO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h96ccc3333ccc96cc)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_L_X10Y109_SLICE_X12Y109_CO6),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(CLBLM_L_X10Y111_SLICE_X12Y111_DO6),
.I5(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_CO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hebc38200ffebc382)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_BLUT (
.I0(CLBLM_L_X10Y111_SLICE_X12Y111_AO5),
.I1(CLBLM_L_X8Y109_SLICE_X11Y109_AO6),
.I2(CLBLM_L_X10Y109_SLICE_X12Y109_CO6),
.I3(CLBLM_L_X10Y111_SLICE_X12Y111_DO6),
.I4(CLBLM_L_X10Y109_SLICE_X13Y109_AO6),
.I5(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_BO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3963c3c69c396)
  ) CLBLM_L_X10Y110_SLICE_X12Y110_ALUT (
.I0(CLBLM_L_X10Y111_SLICE_X12Y111_AO5),
.I1(CLBLM_L_X8Y109_SLICE_X11Y109_AO6),
.I2(CLBLM_L_X10Y109_SLICE_X12Y109_CO6),
.I3(CLBLM_L_X10Y111_SLICE_X12Y111_DO6),
.I4(CLBLM_L_X10Y109_SLICE_X13Y109_AO6),
.I5(CLBLM_L_X10Y109_SLICE_X12Y109_DO6),
.O5(CLBLM_L_X10Y110_SLICE_X12Y110_AO5),
.O6(CLBLM_L_X10Y110_SLICE_X12Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee88e8bbbb22b2)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_DLUT (
.I0(CLBLM_R_X11Y110_SLICE_X14Y110_AO6),
.I1(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I2(CLBLM_R_X11Y110_SLICE_X14Y110_AO5),
.I3(CLBLM_L_X10Y109_SLICE_X12Y109_BO6),
.I4(CLBLM_R_X11Y109_SLICE_X15Y109_AO6),
.I5(CLBLM_L_X10Y109_SLICE_X13Y109_BO6),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_DO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h66cc9c3666cc963c)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_CLUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I2(CLBLM_L_X10Y109_SLICE_X12Y109_BO6),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(CLBLM_R_X11Y109_SLICE_X15Y109_AO6),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_CO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ff0f00fb44b4bb4)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_BLUT (
.I0(CLBLM_L_X10Y109_SLICE_X12Y109_BO6),
.I1(CLBLM_R_X11Y110_SLICE_X14Y110_AO5),
.I2(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I3(CLBLM_L_X10Y109_SLICE_X13Y109_BO6),
.I4(CLBLM_R_X11Y110_SLICE_X14Y110_AO6),
.I5(CLBLM_R_X11Y109_SLICE_X15Y109_AO6),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_BO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0055fff0f0f5ff)
  ) CLBLM_L_X10Y110_SLICE_X13Y110_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(1'b1),
.I2(CLBLM_R_X11Y109_SLICE_X15Y109_AO6),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(CLBLM_L_X10Y109_SLICE_X12Y109_BO6),
.I5(1'b1),
.O5(CLBLM_L_X10Y110_SLICE_X13Y110_AO5),
.O6(CLBLM_L_X10Y110_SLICE_X13Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fdfdfdf134c4c4c)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_DLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_L_X10Y110_SLICE_X13Y110_CO6),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLM_L_X8Y111_SLICE_X11Y111_BO6),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_DO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93936c93936c6c)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_R_X11Y110_SLICE_X14Y110_BO6),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLM_L_X10Y111_SLICE_X12Y111_DO6),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_CO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he64c75df19b38a20)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_BLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(CLBLM_L_X8Y112_SLICE_X11Y112_AO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLM_L_X10Y110_SLICE_X13Y110_AO6),
.I5(CLBLM_L_X10Y110_SLICE_X13Y110_CO6),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_BO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffff0f0fffff)
  ) CLBLM_L_X10Y111_SLICE_X12Y111_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(1'b1),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLM_L_X10Y111_SLICE_X12Y111_AO5),
.O6(CLBLM_L_X10Y111_SLICE_X12Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_DO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_CO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_BO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fdf134cff5f5f00)
  ) CLBLM_L_X10Y111_SLICE_X13Y111_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_R_X11Y110_SLICE_X14Y110_BO6),
.I4(CLBLM_L_X10Y111_SLICE_X12Y111_DO6),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_L_X10Y111_SLICE_X13Y111_AO5),
.O6(CLBLM_L_X10Y111_SLICE_X13Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y104_SLICE_X16Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y104_SLICE_X16Y104_DO5),
.O6(CLBLM_L_X12Y104_SLICE_X16Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0b4b00f000cc0000)
  ) CLBLM_L_X12Y104_SLICE_X16Y104_CLUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(RIOB33_X105Y107_IOB_X1Y108_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(RIOB33_X105Y107_IOB_X1Y107_I),
.O5(CLBLM_L_X12Y104_SLICE_X16Y104_CO5),
.O6(CLBLM_L_X12Y104_SLICE_X16Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h407b7f4422882288)
  ) CLBLM_L_X12Y104_SLICE_X16Y104_BLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y107_IOB_X1Y108_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(RIOB33_X105Y113_IOB_X1Y113_I),
.O5(CLBLM_L_X12Y104_SLICE_X16Y104_BO5),
.O6(CLBLM_L_X12Y104_SLICE_X16Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h778877888d728778)
  ) CLBLM_L_X12Y104_SLICE_X16Y104_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(CLBLM_R_X11Y105_SLICE_X15Y105_AO6),
.I3(CLBLM_L_X12Y104_SLICE_X16Y104_BO6),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X12Y104_SLICE_X16Y104_CO6),
.O5(CLBLM_L_X12Y104_SLICE_X16Y104_AO5),
.O6(CLBLM_L_X12Y104_SLICE_X16Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y104_SLICE_X17Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y104_SLICE_X17Y104_DO5),
.O6(CLBLM_L_X12Y104_SLICE_X17Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y104_SLICE_X17Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y104_SLICE_X17Y104_CO5),
.O6(CLBLM_L_X12Y104_SLICE_X17Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y104_SLICE_X17Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y104_SLICE_X17Y104_BO5),
.O6(CLBLM_L_X12Y104_SLICE_X17Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_L_X12Y104_SLICE_X17Y104_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_L_X12Y104_SLICE_X17Y104_AO5),
.O6(CLBLM_L_X12Y104_SLICE_X17Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y102_SLICE_X2Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y102_SLICE_X2Y102_DO5),
.O6(CLBLM_R_X3Y102_SLICE_X2Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y102_SLICE_X2Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y102_SLICE_X2Y102_CO5),
.O6(CLBLM_R_X3Y102_SLICE_X2Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he2c06ac09548e248)
  ) CLBLM_R_X3Y102_SLICE_X2Y102_BLUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(CLBLM_R_X3Y102_SLICE_X2Y102_AO6),
.O5(CLBLM_R_X3Y102_SLICE_X2Y102_BO5),
.O6(CLBLM_R_X3Y102_SLICE_X2Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4d5f5ddfdfdfffff)
  ) CLBLM_R_X3Y102_SLICE_X2Y102_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLM_R_X3Y102_SLICE_X3Y102_BO6),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(RIOB33_X105Y111_IOB_X1Y111_I),
.O5(CLBLM_R_X3Y102_SLICE_X2Y102_AO5),
.O6(CLBLM_R_X3Y102_SLICE_X2Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y102_SLICE_X3Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y102_SLICE_X3Y102_DO5),
.O6(CLBLM_R_X3Y102_SLICE_X3Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y102_SLICE_X3Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y102_SLICE_X3Y102_CO5),
.O6(CLBLM_R_X3Y102_SLICE_X3Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f7fffff171f3fff)
  ) CLBLM_R_X3Y102_SLICE_X3Y102_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(RIOB33_X105Y111_IOB_X1Y111_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(CLBLM_R_X5Y102_SLICE_X6Y102_CO6),
.O5(CLBLM_R_X3Y102_SLICE_X3Y102_BO5),
.O6(CLBLM_R_X3Y102_SLICE_X3Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffffff71f571f5)
  ) CLBLM_R_X3Y102_SLICE_X3Y102_ALUT (
.I0(CLBLL_L_X4Y103_SLICE_X4Y103_AO5),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(CLBLM_R_X3Y103_SLICE_X3Y103_CO6),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y102_SLICE_X3Y102_AO5),
.O6(CLBLM_R_X3Y102_SLICE_X3Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc33cf00fc33cf00f)
  ) CLBLM_R_X3Y103_SLICE_X2Y103_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y103_SLICE_X3Y103_AO5),
.I2(CLBLM_R_X3Y103_SLICE_X3Y103_DO6),
.I3(CLBLM_R_X3Y102_SLICE_X3Y102_AO5),
.I4(CLBLM_R_X3Y104_SLICE_X2Y104_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y103_SLICE_X2Y103_DO5),
.O6(CLBLM_R_X3Y103_SLICE_X2Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf5dff5f45045505)
  ) CLBLM_R_X3Y103_SLICE_X2Y103_CLUT (
.I0(CLBLL_L_X2Y103_SLICE_X0Y103_CO6),
.I1(CLBLM_R_X3Y103_SLICE_X3Y103_AO5),
.I2(CLBLM_R_X3Y103_SLICE_X3Y103_DO6),
.I3(CLBLM_R_X3Y102_SLICE_X3Y102_AO5),
.I4(CLBLM_R_X3Y104_SLICE_X2Y104_CO6),
.I5(CLBLM_R_X3Y103_SLICE_X2Y103_BO6),
.O5(CLBLM_R_X3Y103_SLICE_X2Y103_CO5),
.O6(CLBLM_R_X3Y103_SLICE_X2Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h557f7fff055707ff)
  ) CLBLM_R_X3Y103_SLICE_X2Y103_BLUT (
.I0(RIOB33_X105Y107_IOB_X1Y108_I),
.I1(LIOB33_X0Y113_IOB_X0Y113_I),
.I2(CLBLL_L_X2Y103_SLICE_X1Y103_BO6),
.I3(CLBLL_L_X2Y103_SLICE_X0Y103_AO6),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLL_L_X4Y102_SLICE_X4Y102_DO6),
.O5(CLBLM_R_X3Y103_SLICE_X2Y103_BO5),
.O6(CLBLM_R_X3Y103_SLICE_X2Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf70808f731cece31)
  ) CLBLM_R_X3Y103_SLICE_X2Y103_ALUT (
.I0(CLBLM_R_X3Y104_SLICE_X2Y104_CO6),
.I1(CLBLM_R_X3Y103_SLICE_X3Y103_DO6),
.I2(CLBLM_R_X3Y103_SLICE_X3Y103_AO5),
.I3(CLBLM_R_X3Y103_SLICE_X2Y103_BO6),
.I4(CLBLL_L_X2Y103_SLICE_X0Y103_CO6),
.I5(CLBLM_R_X3Y102_SLICE_X3Y102_AO5),
.O5(CLBLM_R_X3Y103_SLICE_X2Y103_AO5),
.O6(CLBLM_R_X3Y103_SLICE_X2Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9f5fa39360a05c6c)
  ) CLBLM_R_X3Y103_SLICE_X3Y103_DLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLL_L_X2Y103_SLICE_X1Y103_BO6),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(CLBLL_L_X4Y102_SLICE_X4Y102_DO6),
.I5(CLBLL_L_X2Y103_SLICE_X0Y103_AO6),
.O5(CLBLM_R_X3Y103_SLICE_X3Y103_DO5),
.O6(CLBLM_R_X3Y103_SLICE_X3Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f7f7fff031f13ff)
  ) CLBLM_R_X3Y103_SLICE_X3Y103_CLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(CLBLL_L_X4Y102_SLICE_X4Y102_AO5),
.I2(RIOB33_X105Y107_IOB_X1Y107_I),
.I3(CLBLL_L_X4Y103_SLICE_X4Y103_DO6),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(CLBLL_L_X4Y101_SLICE_X5Y101_AO6),
.O5(CLBLM_R_X3Y103_SLICE_X3Y103_CO5),
.O6(CLBLM_R_X3Y103_SLICE_X3Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha599699969aa5aaa)
  ) CLBLM_R_X3Y103_SLICE_X3Y103_BLUT (
.I0(CLBLL_L_X4Y103_SLICE_X4Y103_DO6),
.I1(CLBLL_L_X4Y101_SLICE_X5Y101_AO6),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(CLBLL_L_X4Y102_SLICE_X4Y102_AO5),
.O5(CLBLM_R_X3Y103_SLICE_X3Y103_BO5),
.O6(CLBLM_R_X3Y103_SLICE_X3Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h9666699982222888)
  ) CLBLM_R_X3Y103_SLICE_X3Y103_ALUT (
.I0(CLBLM_R_X3Y104_SLICE_X3Y104_DO6),
.I1(CLBLL_L_X4Y103_SLICE_X4Y103_AO5),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(CLBLM_R_X3Y103_SLICE_X3Y103_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y103_SLICE_X3Y103_AO5),
.O6(CLBLM_R_X3Y103_SLICE_X3Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc33cc33cc33cc33c)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y104_SLICE_X3Y104_CO6),
.I2(CLBLM_R_X3Y104_SLICE_X3Y104_BO6),
.I3(CLBLM_R_X3Y104_SLICE_X2Y104_AO5),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y104_SLICE_X2Y104_DO5),
.O6(CLBLM_R_X3Y104_SLICE_X2Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haafaeafeeafefaff)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_CLUT (
.I0(CLBLM_R_X3Y103_SLICE_X3Y103_AO6),
.I1(CLBLM_R_X3Y104_SLICE_X2Y104_AO6),
.I2(CLBLM_R_X3Y104_SLICE_X3Y104_BO6),
.I3(CLBLM_R_X3Y104_SLICE_X2Y104_AO5),
.I4(CLBLL_L_X4Y105_SLICE_X4Y105_DO6),
.I5(CLBLL_L_X4Y104_SLICE_X4Y104_BO5),
.O5(CLBLM_R_X3Y104_SLICE_X2Y104_CO5),
.O6(CLBLM_R_X3Y104_SLICE_X2Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbf3b3b233b232302)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_BLUT (
.I0(CLBLL_L_X4Y105_SLICE_X4Y105_DO6),
.I1(CLBLM_R_X3Y104_SLICE_X3Y104_BO6),
.I2(CLBLM_R_X3Y105_SLICE_X3Y105_BO5),
.I3(CLBLL_L_X4Y104_SLICE_X4Y104_BO5),
.I4(CLBLL_L_X4Y104_SLICE_X4Y104_DO6),
.I5(CLBLM_R_X3Y105_SLICE_X3Y105_CO5),
.O5(CLBLM_R_X3Y104_SLICE_X2Y104_BO5),
.O6(CLBLM_R_X3Y104_SLICE_X2Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6969c3c34d4dcfcf)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_ALUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLL_L_X4Y104_SLICE_X4Y104_DO6),
.I2(CLBLM_R_X3Y105_SLICE_X3Y105_BO5),
.I3(1'b1),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y104_SLICE_X2Y104_AO5),
.O6(CLBLM_R_X3Y104_SLICE_X2Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0f4cdf4fdfffff)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_DLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(CLBLL_L_X4Y101_SLICE_X4Y101_CO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLL_L_X4Y103_SLICE_X4Y103_BO5),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLM_R_X3Y103_SLICE_X3Y103_BO6),
.O5(CLBLM_R_X3Y104_SLICE_X3Y104_DO5),
.O6(CLBLM_R_X3Y104_SLICE_X3Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd440fffd4000fdd4)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_CLUT (
.I0(CLBLL_L_X4Y104_SLICE_X4Y104_CO6),
.I1(CLBLL_L_X4Y105_SLICE_X4Y105_BO6),
.I2(CLBLL_L_X4Y106_SLICE_X4Y106_DO6),
.I3(CLBLL_L_X4Y105_SLICE_X4Y105_CO6),
.I4(CLBLM_R_X3Y104_SLICE_X2Y104_AO6),
.I5(CLBLL_L_X4Y106_SLICE_X5Y106_AO5),
.O5(CLBLM_R_X3Y104_SLICE_X3Y104_CO5),
.O6(CLBLM_R_X3Y104_SLICE_X3Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha699599965aa9aaa)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_BLUT (
.I0(CLBLM_R_X3Y103_SLICE_X3Y103_BO6),
.I1(CLBLL_L_X4Y101_SLICE_X4Y101_CO6),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLL_L_X4Y103_SLICE_X4Y103_BO5),
.O5(CLBLM_R_X3Y104_SLICE_X3Y104_BO5),
.O6(CLBLM_R_X3Y104_SLICE_X3Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h9966996687e1781e)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_ALUT (
.I0(CLBLL_L_X4Y106_SLICE_X4Y106_DO6),
.I1(CLBLL_L_X4Y105_SLICE_X4Y105_BO6),
.I2(CLBLM_R_X3Y104_SLICE_X2Y104_AO6),
.I3(CLBLL_L_X4Y104_SLICE_X4Y104_BO6),
.I4(CLBLL_L_X4Y104_SLICE_X4Y104_BO5),
.I5(1'b1),
.O5(CLBLM_R_X3Y104_SLICE_X3Y104_AO5),
.O6(CLBLM_R_X3Y104_SLICE_X3Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y105_SLICE_X2Y105_DO5),
.O6(CLBLM_R_X3Y105_SLICE_X2Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y105_SLICE_X2Y105_CO5),
.O6(CLBLM_R_X3Y105_SLICE_X2Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y105_SLICE_X2Y105_BO5),
.O6(CLBLM_R_X3Y105_SLICE_X2Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0f00f0ff0f0)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X3Y103_SLICE_X3Y103_AO6),
.I3(1'b1),
.I4(CLBLM_R_X3Y104_SLICE_X2Y104_BO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y105_SLICE_X2Y105_AO5),
.O6(CLBLM_R_X3Y105_SLICE_X2Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93936ca05f5fa0)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_DLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(CLBLM_R_X3Y105_SLICE_X3Y105_AO5),
.I4(CLBLL_L_X4Y103_SLICE_X5Y103_CO6),
.I5(LIOB33_X0Y113_IOB_X0Y113_I),
.O5(CLBLM_R_X3Y105_SLICE_X3Y105_DO5),
.O6(CLBLM_R_X3Y105_SLICE_X3Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff5f5f5f5f)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_CLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(1'b1),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(LIOB33_X0Y111_IOB_X0Y111_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y105_SLICE_X3Y105_CO5),
.O6(CLBLM_R_X3Y105_SLICE_X3Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff66cc9933)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLL_L_X4Y103_SLICE_X4Y103_BO5),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(CLBLL_L_X4Y101_SLICE_X4Y101_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y105_SLICE_X3Y105_BO5),
.O6(CLBLM_R_X3Y105_SLICE_X3Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff69699999)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_ALUT (
.I0(CLBLL_L_X4Y105_SLICE_X5Y105_BO6),
.I1(CLBLL_L_X4Y104_SLICE_X4Y104_AO6),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y105_SLICE_X3Y105_AO5),
.O6(CLBLM_R_X3Y105_SLICE_X3Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_DO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_CO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_BO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_AO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_DO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_CO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_BO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0ccc03330ccccfff)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y106_SLICE_X4Y106_AO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(CLBLM_R_X5Y105_SLICE_X6Y105_BO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_AO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555aaaaaaaa)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_DLUT (
.I0(CLBLL_L_X4Y107_SLICE_X5Y107_BO6),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLM_R_X3Y107_SLICE_X2Y107_BO6),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_DO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999a55596665aaa)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_CLUT (
.I0(CLBLM_R_X5Y106_SLICE_X7Y106_DO6),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLL_L_X4Y107_SLICE_X5Y107_CO6),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_CO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f13df4cff5f5f00)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(LIOB33_X0Y113_IOB_X0Y113_I),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(CLBLL_L_X4Y107_SLICE_X5Y107_CO6),
.I4(CLBLM_R_X5Y106_SLICE_X7Y106_DO6),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_BO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa5500ff93939393)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(CLBLM_R_X3Y107_SLICE_X3Y107_DO5),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLL_L_X4Y109_SLICE_X4Y109_BO6),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_AO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33cc33cc5555aaaa)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_DLUT (
.I0(CLBLM_R_X5Y105_SLICE_X6Y105_BO6),
.I1(CLBLM_R_X3Y107_SLICE_X2Y107_CO6),
.I2(1'b1),
.I3(CLBLL_L_X4Y108_SLICE_X5Y108_CO6),
.I4(CLBLL_L_X4Y106_SLICE_X4Y106_AO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_DO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h8000000000008000)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_CLUT (
.I0(CLBLM_R_X3Y105_SLICE_X3Y105_BO6),
.I1(CLBLL_L_X4Y108_SLICE_X4Y108_CO6),
.I2(CLBLM_R_X5Y105_SLICE_X6Y105_AO6),
.I3(CLBLM_R_X5Y108_SLICE_X7Y108_BO6),
.I4(CLBLL_L_X4Y106_SLICE_X4Y106_AO6),
.I5(CLBLM_R_X5Y105_SLICE_X6Y105_BO6),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_CO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc48ffde088cceef)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_BLUT (
.I0(CLBLL_L_X4Y108_SLICE_X5Y108_CO6),
.I1(CLBLM_R_X3Y107_SLICE_X2Y107_BO6),
.I2(CLBLM_R_X3Y107_SLICE_X2Y107_CO6),
.I3(CLBLL_L_X4Y108_SLICE_X5Y108_BO6),
.I4(CLBLL_L_X4Y107_SLICE_X5Y107_BO6),
.I5(CLBLM_R_X3Y107_SLICE_X3Y107_CO6),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_BO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'he999999999999999)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_ALUT (
.I0(CLBLM_R_X3Y107_SLICE_X3Y107_DO6),
.I1(CLBLL_L_X4Y108_SLICE_X5Y108_BO6),
.I2(CLBLM_R_X3Y106_SLICE_X3Y106_AO6),
.I3(CLBLM_R_X5Y105_SLICE_X6Y105_AO6),
.I4(CLBLL_L_X4Y108_SLICE_X4Y108_CO6),
.I5(CLBLM_R_X5Y108_SLICE_X7Y108_BO6),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_AO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_DO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_CO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_BO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_AO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_DO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_CO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_BO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aaa566696666555)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_ALUT (
.I0(CLBLM_R_X3Y107_SLICE_X2Y107_DO6),
.I1(CLBLL_L_X4Y108_SLICE_X5Y108_CO6),
.I2(CLBLM_R_X3Y106_SLICE_X3Y106_AO6),
.I3(CLBLM_R_X5Y108_SLICE_X6Y108_DO6),
.I4(CLBLM_R_X3Y107_SLICE_X2Y107_CO6),
.I5(CLBLL_L_X4Y108_SLICE_X5Y108_BO6),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_AO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_DO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_CO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2a200a20959f359f)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_BLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_BO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a555550f0fffff)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_ALUT (
.I0(CLBLL_L_X2Y111_SLICE_X0Y111_DO6),
.I1(1'b1),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(1'b1),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_AO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_DO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_CO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_BO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aa5aa553f3f3f3f)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_ALUT (
.I0(CLBLM_R_X3Y110_SLICE_X3Y110_BO6),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(CLBLL_L_X4Y109_SLICE_X4Y109_AO6),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_AO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3963ca50f5af0)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_DLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I2(CLBLM_R_X3Y111_SLICE_X3Y111_DO6),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(CLBLM_R_X5Y110_SLICE_X6Y110_DO6),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_DO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0b4b00f000cc0000)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_CLUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_CO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h138a1b0a64a8e428)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_BLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_BO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h02a25da277228888)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_ALUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_AO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_DO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_CO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2bb2bb22affaffaa)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_BLUT (
.I0(CLBLM_R_X3Y111_SLICE_X3Y111_DO6),
.I1(LIOB33_X0Y111_IOB_X0Y111_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(CLBLM_R_X5Y110_SLICE_X6Y110_DO6),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_BO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h999933330f0fffff)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_ALUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(CLBLM_R_X3Y111_SLICE_X3Y111_CO6),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(1'b1),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_AO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a56a5a9a5a95a56)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_DLUT (
.I0(CLBLM_R_X3Y110_SLICE_X2Y110_BO6),
.I1(CLBLM_R_X3Y111_SLICE_X3Y111_AO5),
.I2(CLBLM_R_X3Y110_SLICE_X2Y110_CO6),
.I3(CLBLM_R_X3Y110_SLICE_X2Y110_AO6),
.I4(CLBLM_R_X3Y111_SLICE_X3Y111_AO6),
.I5(CLBLL_L_X2Y111_SLICE_X1Y111_AO6),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_DO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfafef5fda0a85054)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_CLUT (
.I0(CLBLM_R_X3Y110_SLICE_X2Y110_BO6),
.I1(CLBLM_R_X3Y111_SLICE_X3Y111_AO5),
.I2(CLBLM_R_X3Y110_SLICE_X2Y110_CO6),
.I3(CLBLM_R_X3Y110_SLICE_X2Y110_AO6),
.I4(CLBLM_R_X3Y111_SLICE_X3Y111_AO6),
.I5(CLBLL_L_X2Y111_SLICE_X1Y111_AO6),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_CO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cf0c30f3bf7c408)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(CLBLM_R_X3Y110_SLICE_X2Y110_CO6),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(CLBLM_R_X3Y110_SLICE_X2Y110_BO6),
.I5(CLBLM_R_X3Y110_SLICE_X2Y110_AO6),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_BO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha50fa50fcdcfcdcf)
  ) CLBLM_R_X3Y111_SLICE_X2Y111_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(CLBLM_R_X3Y110_SLICE_X2Y110_CO6),
.I2(CLBLM_R_X3Y110_SLICE_X2Y110_AO6),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y111_SLICE_X2Y111_AO5),
.O6(CLBLM_R_X3Y111_SLICE_X2Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h57155f177f1fff3f)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_DLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(CLBLL_L_X4Y111_SLICE_X4Y111_DO6),
.I2(CLBLM_R_X5Y111_SLICE_X6Y111_DO6),
.I3(CLBLM_R_X3Y113_SLICE_X3Y113_CO6),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_DO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h93c9cc3c6c36cc3c)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_CLUT (
.I0(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I1(CLBLM_R_X5Y111_SLICE_X6Y111_BO6),
.I2(CLBLL_L_X4Y111_SLICE_X4Y111_DO6),
.I3(CLBLM_R_X3Y113_SLICE_X3Y113_CO6),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_CO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff69699999)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_BLUT (
.I0(CLBLM_R_X3Y113_SLICE_X3Y113_CO6),
.I1(CLBLL_L_X4Y111_SLICE_X4Y111_DO6),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_BO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff3333ffff)
  ) CLBLM_R_X3Y111_SLICE_X3Y111_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(1'b1),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y111_SLICE_X3Y111_AO5),
.O6(CLBLM_R_X3Y111_SLICE_X3Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_DO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4d8e8e8eddeeeeee)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_CLUT (
.I0(CLBLM_R_X3Y111_SLICE_X2Y111_BO6),
.I1(CLBLL_L_X2Y111_SLICE_X1Y111_DO6),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_CO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2bafbbff8e0aeeaa)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_BLUT (
.I0(CLBLL_L_X2Y112_SLICE_X1Y112_CO6),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I5(CLBLL_L_X2Y111_SLICE_X1Y111_CO6),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_BO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3963ca50f5af0)
  ) CLBLM_R_X3Y112_SLICE_X2Y112_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(CLBLL_L_X2Y111_SLICE_X1Y111_DO6),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(CLBLM_R_X3Y111_SLICE_X2Y111_BO6),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_R_X3Y112_SLICE_X2Y112_AO5),
.O6(CLBLM_R_X3Y112_SLICE_X2Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_DO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3963c993366cc)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(CLBLL_L_X4Y111_SLICE_X4Y111_CO6),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLM_R_X3Y112_SLICE_X2Y112_CO6),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_CO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he6194cb3758adf20)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X3Y112_SLICE_X2Y112_BO6),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(CLBLL_L_X4Y112_SLICE_X4Y112_CO6),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(CLBLM_R_X3Y112_SLICE_X3Y112_CO6),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_BO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf00f00ff5555ffff)
  ) CLBLM_R_X3Y112_SLICE_X3Y112_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(1'b1),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_BO6),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y112_SLICE_X3Y112_AO5),
.O6(CLBLM_R_X3Y112_SLICE_X3Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdc4dc40f7317310)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_DLUT (
.I0(CLBLM_R_X3Y112_SLICE_X2Y112_AO6),
.I1(CLBLL_L_X4Y112_SLICE_X4Y112_BO6),
.I2(CLBLL_L_X2Y112_SLICE_X1Y112_CO6),
.I3(CLBLM_R_X3Y113_SLICE_X2Y113_AO5),
.I4(CLBLM_R_X3Y113_SLICE_X2Y113_BO5),
.I5(CLBLM_R_X3Y113_SLICE_X2Y113_BO6),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_DO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb43cd29678f01e5a)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_CLUT (
.I0(CLBLM_R_X3Y112_SLICE_X2Y112_AO6),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(CLBLL_L_X4Y112_SLICE_X4Y112_BO6),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(CLBLL_L_X2Y112_SLICE_X1Y112_CO6),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_CO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffff00ffffff)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_BLUT (
.I0(1'b1),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(1'b1),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_BO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0000fff0fff0fff)
  ) CLBLM_R_X3Y113_SLICE_X2Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(CLBLM_R_X3Y113_SLICE_X2Y113_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y113_SLICE_X2Y113_AO5),
.O6(CLBLM_R_X3Y113_SLICE_X2Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_DO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6affffff006a6a6a)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_CLUT (
.I0(CLBLL_L_X4Y113_SLICE_X4Y113_AO6),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(CLBLM_R_X3Y113_SLICE_X3Y113_BO6),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_CO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffbf3f153f2a00)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(CLBLL_L_X4Y112_SLICE_X4Y112_CO6),
.I5(CLBLM_R_X3Y113_SLICE_X2Y113_DO6),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_BO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a95956a956a956a)
  ) CLBLM_R_X3Y113_SLICE_X3Y113_ALUT (
.I0(CLBLM_R_X3Y113_SLICE_X3Y113_BO6),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(CLBLL_L_X4Y113_SLICE_X4Y113_AO6),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.O5(CLBLM_R_X3Y113_SLICE_X3Y113_AO5),
.O6(CLBLM_R_X3Y113_SLICE_X3Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y100_SLICE_X6Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y100_SLICE_X6Y100_DO5),
.O6(CLBLM_R_X5Y100_SLICE_X6Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y100_SLICE_X6Y100_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y100_SLICE_X6Y100_CO5),
.O6(CLBLM_R_X5Y100_SLICE_X6Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h87f078f0e13c1e3c)
  ) CLBLM_R_X5Y100_SLICE_X6Y100_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(CLBLM_R_X7Y100_SLICE_X8Y100_AO6),
.I2(CLBLM_R_X5Y100_SLICE_X7Y100_AO6),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(CLBLM_R_X7Y100_SLICE_X8Y100_BO6),
.O5(CLBLM_R_X5Y100_SLICE_X6Y100_BO5),
.O6(CLBLM_R_X5Y100_SLICE_X6Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h07017f1fff3fff3f)
  ) CLBLM_R_X5Y100_SLICE_X6Y100_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(CLBLM_R_X7Y100_SLICE_X8Y100_AO6),
.I2(CLBLM_R_X5Y100_SLICE_X7Y100_AO6),
.I3(CLBLM_R_X7Y100_SLICE_X8Y100_BO6),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(RIOB33_X105Y107_IOB_X1Y107_I),
.O5(CLBLM_R_X5Y100_SLICE_X6Y100_AO5),
.O6(CLBLM_R_X5Y100_SLICE_X6Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y100_SLICE_X7Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y100_SLICE_X7Y100_DO5),
.O6(CLBLM_R_X5Y100_SLICE_X7Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y100_SLICE_X7Y100_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y100_SLICE_X7Y100_CO5),
.O6(CLBLM_R_X5Y100_SLICE_X7Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y100_SLICE_X7Y100_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y100_SLICE_X7Y100_BO5),
.O6(CLBLM_R_X5Y100_SLICE_X7Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h9a6a6a6a95959a6a)
  ) CLBLM_R_X5Y100_SLICE_X7Y100_ALUT (
.I0(CLBLM_R_X5Y102_SLICE_X7Y102_CO6),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(RIOB33_X105Y107_IOB_X1Y108_I),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(CLBLM_R_X7Y102_SLICE_X9Y102_DO6),
.I5(CLBLM_R_X7Y101_SLICE_X8Y101_AO5),
.O5(CLBLM_R_X5Y100_SLICE_X7Y100_AO5),
.O6(CLBLM_R_X5Y100_SLICE_X7Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7df51450ffff3cf0)
  ) CLBLM_R_X5Y101_SLICE_X6Y101_DLUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(CLBLM_R_X5Y102_SLICE_X6Y102_BO6),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(CLBLM_R_X5Y102_SLICE_X7Y102_AO5),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLM_R_X5Y101_SLICE_X6Y101_DO5),
.O6(CLBLM_R_X5Y101_SLICE_X6Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc66c93936c6cc66c)
  ) CLBLM_R_X5Y101_SLICE_X6Y101_CLUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(CLBLL_L_X4Y102_SLICE_X5Y102_CO6),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(CLBLM_R_X5Y102_SLICE_X7Y102_AO5),
.I5(CLBLM_R_X5Y102_SLICE_X7Y102_BO6),
.O5(CLBLM_R_X5Y101_SLICE_X6Y101_CO5),
.O6(CLBLM_R_X5Y101_SLICE_X6Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a959595956a6a6a)
  ) CLBLM_R_X5Y101_SLICE_X6Y101_BLUT (
.I0(CLBLM_R_X5Y102_SLICE_X7Y102_AO5),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(CLBLM_R_X5Y102_SLICE_X6Y102_BO6),
.O5(CLBLM_R_X5Y101_SLICE_X6Y101_BO5),
.O6(CLBLM_R_X5Y101_SLICE_X6Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff2b2bbbbb)
  ) CLBLM_R_X5Y101_SLICE_X6Y101_ALUT (
.I0(CLBLM_R_X5Y101_SLICE_X6Y101_DO6),
.I1(CLBLL_L_X4Y102_SLICE_X5Y102_CO6),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y101_SLICE_X6Y101_AO5),
.O6(CLBLM_R_X5Y101_SLICE_X6Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h571177577f33ff7f)
  ) CLBLM_R_X5Y101_SLICE_X7Y101_DLUT (
.I0(RIOB33_X105Y107_IOB_X1Y108_I),
.I1(CLBLM_R_X5Y102_SLICE_X7Y102_CO6),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(CLBLM_R_X7Y101_SLICE_X8Y101_AO5),
.I4(CLBLM_R_X7Y102_SLICE_X9Y102_DO6),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLM_R_X5Y101_SLICE_X7Y101_DO5),
.O6(CLBLM_R_X5Y101_SLICE_X7Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h04df0ddf4fdfdfdf)
  ) CLBLM_R_X5Y101_SLICE_X7Y101_CLUT (
.I0(CLBLM_R_X7Y101_SLICE_X8Y101_CO5),
.I1(CLBLM_R_X7Y102_SLICE_X8Y102_AO5),
.I2(CLBLM_R_X5Y100_SLICE_X6Y100_BO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X5Y101_SLICE_X7Y101_CO5),
.O6(CLBLM_R_X5Y101_SLICE_X7Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he64c75df19b38a20)
  ) CLBLM_R_X5Y101_SLICE_X7Y101_BLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_R_X7Y102_SLICE_X8Y102_AO5),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(CLBLM_R_X7Y101_SLICE_X8Y101_CO5),
.I5(CLBLM_R_X5Y100_SLICE_X6Y100_BO6),
.O5(CLBLM_R_X5Y101_SLICE_X7Y101_BO5),
.O6(CLBLM_R_X5Y101_SLICE_X7Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffffff69996999)
  ) CLBLM_R_X5Y101_SLICE_X7Y101_ALUT (
.I0(CLBLM_R_X5Y101_SLICE_X7Y101_DO6),
.I1(CLBLM_R_X5Y101_SLICE_X6Y101_BO6),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y101_SLICE_X7Y101_AO5),
.O6(CLBLM_R_X5Y101_SLICE_X7Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff00ffffffffff)
  ) CLBLM_R_X5Y102_SLICE_X6Y102_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(1'b1),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X5Y102_SLICE_X6Y102_DO5),
.O6(CLBLM_R_X5Y102_SLICE_X6Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h44dfdfff5ddfffff)
  ) CLBLM_R_X5Y102_SLICE_X6Y102_CLUT (
.I0(RIOB33_X105Y109_IOB_X1Y110_I),
.I1(CLBLM_R_X7Y105_SLICE_X8Y105_AO6),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(LIOB33_X0Y101_IOB_X0Y101_I),
.O5(CLBLM_R_X5Y102_SLICE_X6Y102_CO5),
.O6(CLBLM_R_X5Y102_SLICE_X6Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd333cb93ffff3fff)
  ) CLBLM_R_X5Y102_SLICE_X6Y102_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(CLBLM_R_X5Y102_SLICE_X6Y102_CO6),
.I5(RIOB33_X105Y111_IOB_X1Y111_I),
.O5(CLBLM_R_X5Y102_SLICE_X6Y102_BO5),
.O6(CLBLM_R_X5Y102_SLICE_X6Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999966666699996)
  ) CLBLM_R_X5Y102_SLICE_X6Y102_ALUT (
.I0(CLBLM_R_X5Y102_SLICE_X6Y102_DO6),
.I1(CLBLM_R_X7Y102_SLICE_X8Y102_CO6),
.I2(CLBLM_R_X7Y104_SLICE_X8Y104_AO5),
.I3(CLBLM_R_X7Y103_SLICE_X8Y103_DO6),
.I4(CLBLM_R_X5Y100_SLICE_X6Y100_BO6),
.I5(CLBLM_R_X7Y102_SLICE_X8Y102_BO6),
.O5(CLBLM_R_X5Y102_SLICE_X6Y102_AO5),
.O6(CLBLM_R_X5Y102_SLICE_X6Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h60a0f6faf6faf6fa)
  ) CLBLM_R_X5Y102_SLICE_X7Y102_DLUT (
.I0(CLBLM_R_X5Y103_SLICE_X7Y103_AO6),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(CLBLM_R_X7Y103_SLICE_X8Y103_AO5),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_R_X5Y102_SLICE_X7Y102_DO5),
.O6(CLBLM_R_X5Y102_SLICE_X7Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9c6339c6c3c3cccc)
  ) CLBLM_R_X5Y102_SLICE_X7Y102_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLL_L_X4Y102_SLICE_X5Y102_DO6),
.I2(CLBLM_R_X7Y103_SLICE_X8Y103_AO5),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(CLBLM_R_X5Y102_SLICE_X7Y102_BO5),
.I5(RIOB33_X105Y109_IOB_X1Y109_I),
.O5(CLBLM_R_X5Y102_SLICE_X7Y102_CO5),
.O6(CLBLM_R_X5Y102_SLICE_X7Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h99339933f00f0f0f)
  ) CLBLM_R_X5Y102_SLICE_X7Y102_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLM_R_X5Y102_SLICE_X6Y102_BO6),
.I2(CLBLM_R_X5Y103_SLICE_X7Y103_AO6),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y102_SLICE_X7Y102_BO5),
.O6(CLBLM_R_X5Y102_SLICE_X7Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffffff2b2bafaf)
  ) CLBLM_R_X5Y102_SLICE_X7Y102_ALUT (
.I0(CLBLM_R_X5Y102_SLICE_X7Y102_DO6),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(CLBLL_L_X4Y102_SLICE_X5Y102_DO6),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(RIOB33_X105Y109_IOB_X1Y109_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y102_SLICE_X7Y102_AO5),
.O6(CLBLM_R_X5Y102_SLICE_X7Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb4d23c96781ef05a)
  ) CLBLM_R_X5Y103_SLICE_X6Y103_DLUT (
.I0(CLBLM_R_X5Y104_SLICE_X6Y104_AO6),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(CLBLM_R_X5Y104_SLICE_X6Y104_DO6),
.I3(CLBLM_R_X5Y105_SLICE_X6Y105_DO6),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(LIOB33_X0Y113_IOB_X0Y113_I),
.O5(CLBLM_R_X5Y103_SLICE_X6Y103_DO5),
.O6(CLBLM_R_X5Y103_SLICE_X6Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h37133f177f1fff5f)
  ) CLBLM_R_X5Y103_SLICE_X6Y103_CLUT (
.I0(CLBLM_R_X5Y104_SLICE_X6Y104_AO6),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(CLBLM_R_X5Y104_SLICE_X6Y104_DO6),
.I3(CLBLM_R_X5Y105_SLICE_X6Y105_DO6),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(LIOB33_X0Y113_IOB_X0Y113_I),
.O5(CLBLM_R_X5Y103_SLICE_X6Y103_CO5),
.O6(CLBLM_R_X5Y103_SLICE_X6Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h639cc6399c6339c6)
  ) CLBLM_R_X5Y103_SLICE_X6Y103_BLUT (
.I0(CLBLM_R_X7Y104_SLICE_X9Y104_AO5),
.I1(CLBLM_R_X7Y103_SLICE_X8Y103_DO6),
.I2(CLBLM_R_X7Y103_SLICE_X8Y103_CO6),
.I3(CLBLM_R_X7Y102_SLICE_X8Y102_BO6),
.I4(CLBLM_R_X5Y103_SLICE_X6Y103_AO6),
.I5(CLBLM_R_X7Y104_SLICE_X8Y104_AO5),
.O5(CLBLM_R_X5Y103_SLICE_X6Y103_BO5),
.O6(CLBLM_R_X5Y103_SLICE_X6Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff2baf2baf)
  ) CLBLM_R_X5Y103_SLICE_X6Y103_ALUT (
.I0(CLBLM_R_X7Y104_SLICE_X9Y104_AO5),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(CLBLM_R_X7Y103_SLICE_X8Y103_CO6),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y103_SLICE_X6Y103_AO5),
.O6(CLBLM_R_X5Y103_SLICE_X6Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y103_SLICE_X7Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y103_SLICE_X7Y103_DO5),
.O6(CLBLM_R_X5Y103_SLICE_X7Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y103_SLICE_X7Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y103_SLICE_X7Y103_CO5),
.O6(CLBLM_R_X5Y103_SLICE_X7Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y103_SLICE_X7Y103_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y103_SLICE_X7Y103_BO5),
.O6(CLBLM_R_X5Y103_SLICE_X7Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb79b77f7f7977777)
  ) CLBLM_R_X5Y103_SLICE_X7Y103_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(RIOB33_X105Y111_IOB_X1Y111_I),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(CLBLM_R_X7Y105_SLICE_X8Y105_AO6),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(LIOB33_X0Y101_IOB_X0Y101_I),
.O5(CLBLM_R_X5Y103_SLICE_X7Y103_AO5),
.O6(CLBLM_R_X5Y103_SLICE_X7Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a9696a5a569695a)
  ) CLBLM_R_X5Y104_SLICE_X6Y104_DLUT (
.I0(CLBLL_L_X4Y103_SLICE_X5Y103_AO6),
.I1(CLBLM_R_X5Y104_SLICE_X7Y104_AO6),
.I2(CLBLL_L_X4Y104_SLICE_X5Y104_AO5),
.I3(CLBLM_R_X7Y104_SLICE_X9Y104_BO6),
.I4(CLBLM_R_X5Y105_SLICE_X6Y105_AO5),
.I5(CLBLM_R_X5Y103_SLICE_X6Y103_BO6),
.O5(CLBLM_R_X5Y104_SLICE_X6Y104_DO5),
.O6(CLBLM_R_X5Y104_SLICE_X6Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h87e1ff33781e00cc)
  ) CLBLM_R_X5Y104_SLICE_X6Y104_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(CLBLM_R_X5Y104_SLICE_X7Y104_AO6),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(CLBLM_R_X7Y104_SLICE_X9Y104_BO6),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(CLBLM_R_X5Y103_SLICE_X6Y103_BO6),
.O5(CLBLM_R_X5Y104_SLICE_X6Y104_CO5),
.O6(CLBLM_R_X5Y104_SLICE_X6Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9af059ff650fa600)
  ) CLBLM_R_X5Y104_SLICE_X6Y104_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(CLBLM_R_X5Y105_SLICE_X6Y105_DO6),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(CLBLM_R_X5Y104_SLICE_X6Y104_AO6),
.I5(CLBLM_R_X5Y104_SLICE_X6Y104_CO6),
.O5(CLBLM_R_X5Y104_SLICE_X6Y104_BO5),
.O6(CLBLM_R_X5Y104_SLICE_X6Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h999955553f03ff0f)
  ) CLBLM_R_X5Y104_SLICE_X6Y104_ALUT (
.I0(CLBLM_R_X5Y104_SLICE_X7Y104_AO5),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(CLBLM_R_X5Y104_SLICE_X7Y104_AO6),
.I3(CLBLM_R_X7Y104_SLICE_X9Y104_BO6),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y104_SLICE_X6Y104_AO5),
.O6(CLBLM_R_X5Y104_SLICE_X6Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y104_SLICE_X7Y104_DO5),
.O6(CLBLM_R_X5Y104_SLICE_X7Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y104_SLICE_X7Y104_CO5),
.O6(CLBLM_R_X5Y104_SLICE_X7Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y104_SLICE_X7Y104_BO5),
.O6(CLBLM_R_X5Y104_SLICE_X7Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5af0a50f963c69c3)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_ALUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(CLBLM_R_X7Y104_SLICE_X9Y104_BO6),
.I2(CLBLM_R_X7Y104_SLICE_X9Y104_AO5),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(CLBLM_R_X7Y103_SLICE_X8Y103_CO6),
.I5(1'b1),
.O5(CLBLM_R_X5Y104_SLICE_X7Y104_AO5),
.O6(CLBLM_R_X5Y104_SLICE_X7Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h48dedede88eeeeee)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_DLUT (
.I0(CLBLM_R_X7Y104_SLICE_X9Y104_DO6),
.I1(CLBLM_R_X7Y106_SLICE_X9Y106_CO6),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_DO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999966696669666)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_CLUT (
.I0(CLBLM_R_X7Y104_SLICE_X9Y104_DO6),
.I1(CLBLM_R_X7Y106_SLICE_X9Y106_CO6),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_CO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3963c963c963c)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_BLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(CLBLM_R_X5Y105_SLICE_X6Y105_DO6),
.I2(CLBLM_R_X5Y104_SLICE_X7Y104_AO5),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(LIOB33_X0Y111_IOB_X0Y112_I),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_BO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5050f0f05555ffff)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(1'b1),
.I2(CLBLM_R_X5Y104_SLICE_X7Y104_AO5),
.I3(1'b1),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_AO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7df51450ffff3cf0)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_DLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(LIOB33_X0Y109_IOB_X0Y109_I),
.I2(CLBLM_R_X7Y102_SLICE_X8Y102_DO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X7Y103_SLICE_X8Y103_DO6),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_DO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3963ca50f5af0)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(CLBLM_R_X7Y102_SLICE_X8Y102_DO6),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(CLBLM_R_X7Y103_SLICE_X8Y103_DO6),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_CO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h696999992b2bbbbb)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_BLUT (
.I0(CLBLM_R_X5Y105_SLICE_X7Y105_DO6),
.I1(CLBLM_R_X5Y101_SLICE_X7Y101_BO6),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(1'b1),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_BO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff5f5f5f5f)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_ALUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(1'b1),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_AO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdb24718e59a6f30c)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_DLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(CLBLM_R_X5Y107_SLICE_X6Y107_BO6),
.I2(CLBLM_R_X5Y106_SLICE_X7Y106_BO6),
.I3(CLBLM_R_X5Y106_SLICE_X6Y106_CO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_DO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'ha956956a956aa956)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_CLUT (
.I0(CLBLM_R_X7Y106_SLICE_X9Y106_DO6),
.I1(CLBLM_R_X5Y105_SLICE_X7Y105_AO5),
.I2(CLBLM_L_X8Y107_SLICE_X10Y107_CO6),
.I3(CLBLM_R_X5Y106_SLICE_X6Y106_AO5),
.I4(CLBLM_R_X7Y107_SLICE_X9Y107_AO5),
.I5(CLBLM_R_X7Y106_SLICE_X9Y106_BO6),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_CO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f15ff3fd540ffc0)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_BLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(CLBLM_L_X8Y107_SLICE_X10Y107_CO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_R_X7Y106_SLICE_X9Y106_BO6),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_BO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h55ff55ff5f5f5f5f)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_ALUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(1'b1),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_AO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6966969999696696)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_DLUT (
.I0(CLBLM_R_X5Y106_SLICE_X7Y106_AO6),
.I1(CLBLM_R_X5Y106_SLICE_X7Y106_BO6),
.I2(CLBLM_R_X5Y106_SLICE_X7Y106_AO5),
.I3(CLBLM_R_X5Y106_SLICE_X7Y106_CO6),
.I4(CLBLM_R_X5Y107_SLICE_X6Y107_BO6),
.I5(CLBLM_R_X5Y107_SLICE_X7Y107_BO6),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_DO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887877887788778)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_CLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_R_X7Y107_SLICE_X8Y107_CO6),
.I3(CLBLM_L_X8Y106_SLICE_X10Y106_CO6),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_CO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f07ff77f7707700)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_BLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_R_X7Y107_SLICE_X8Y107_CO6),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLM_L_X8Y106_SLICE_X10Y106_CO6),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_BO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff3f3f3f3f)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_AO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h71d4f3fcd471fcf3)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_DLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(CLBLM_R_X5Y106_SLICE_X7Y106_BO6),
.I2(CLBLM_R_X5Y107_SLICE_X7Y107_DO6),
.I3(CLBLM_R_X5Y106_SLICE_X7Y106_AO6),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(CLBLM_R_X5Y107_SLICE_X6Y107_BO6),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_DO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h507570ff55f7f7ff)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(CLBLM_R_X5Y106_SLICE_X7Y106_BO6),
.I3(CLBLL_L_X4Y106_SLICE_X4Y106_AO5),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(CLBLM_R_X5Y107_SLICE_X6Y107_BO6),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_CO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c939393936c6c6c)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_BLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(CLBLM_R_X7Y106_SLICE_X9Y106_BO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(CLBLM_L_X8Y107_SLICE_X10Y107_CO6),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_BO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887878787787878)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_ALUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(CLBLM_R_X7Y107_SLICE_X8Y107_BO6),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLM_R_X7Y108_SLICE_X8Y108_AO6),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_AO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8808f08fee0ef0e)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_DLUT (
.I0(CLBLM_R_X5Y106_SLICE_X6Y106_AO6),
.I1(CLBLM_R_X7Y108_SLICE_X8Y108_AO6),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_DO6),
.I3(CLBLM_R_X5Y106_SLICE_X7Y106_AO5),
.I4(CLBLM_R_X5Y105_SLICE_X7Y105_AO6),
.I5(CLBLM_R_X7Y107_SLICE_X8Y107_AO6),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_DO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h788787781ee1e11e)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_CLUT (
.I0(CLBLM_R_X5Y106_SLICE_X6Y106_AO6),
.I1(CLBLM_R_X7Y108_SLICE_X8Y108_AO6),
.I2(CLBLM_L_X8Y107_SLICE_X10Y107_DO6),
.I3(CLBLM_R_X7Y107_SLICE_X8Y107_CO6),
.I4(CLBLM_R_X5Y105_SLICE_X7Y105_AO6),
.I5(CLBLM_R_X7Y107_SLICE_X8Y107_AO6),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_CO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4cdf80ecdfdfecec)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLM_R_X7Y108_SLICE_X8Y108_AO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(CLBLM_R_X7Y107_SLICE_X8Y107_BO6),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_BO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a9556a9956aa956)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_ALUT (
.I0(CLBLM_R_X5Y105_SLICE_X7Y105_AO6),
.I1(CLBLM_R_X7Y108_SLICE_X8Y108_AO6),
.I2(CLBLM_R_X5Y106_SLICE_X6Y106_AO6),
.I3(CLBLM_R_X7Y107_SLICE_X9Y107_DO6),
.I4(CLBLM_R_X7Y107_SLICE_X8Y107_AO6),
.I5(CLBLM_R_X5Y106_SLICE_X7Y106_AO5),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_AO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0080000000000000)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_DLUT (
.I0(CLBLM_R_X5Y105_SLICE_X6Y105_AO6),
.I1(CLBLL_L_X4Y108_SLICE_X4Y108_CO6),
.I2(CLBLM_R_X5Y108_SLICE_X7Y108_DO6),
.I3(CLBLM_R_X7Y106_SLICE_X9Y106_BO6),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_DO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f7f07373fff1777)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_CLUT (
.I0(CLBLM_R_X5Y108_SLICE_X6Y108_AO6),
.I1(CLBLM_R_X5Y108_SLICE_X7Y108_CO6),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(LIOB33_X0Y113_IOB_X0Y113_I),
.I4(CLBLM_R_X5Y109_SLICE_X6Y109_CO6),
.I5(LIOB33_X0Y111_IOB_X0Y112_I),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_CO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he169783c2da5b4f0)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_BLUT (
.I0(CLBLM_R_X5Y109_SLICE_X6Y109_CO6),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(CLBLM_R_X5Y108_SLICE_X7Y108_CO6),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(CLBLM_R_X5Y108_SLICE_X6Y108_AO6),
.I5(LIOB33_X0Y113_IOB_X0Y113_I),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_BO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a5965a965a965a)
  ) CLBLM_R_X5Y108_SLICE_X6Y108_ALUT (
.I0(CLBLM_R_X5Y109_SLICE_X6Y109_DO6),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(CLBLM_R_X7Y108_SLICE_X8Y108_CO6),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLM_R_X5Y108_SLICE_X6Y108_AO5),
.O6(CLBLM_R_X5Y108_SLICE_X6Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0400040000000000)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_DLUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_AO6),
.I1(CLBLM_L_X10Y108_SLICE_X13Y108_BO6),
.I2(CLBLM_R_X7Y112_SLICE_X8Y112_AO6),
.I3(CLBLM_R_X5Y109_SLICE_X7Y109_DO6),
.I4(1'b1),
.I5(CLBLM_L_X8Y109_SLICE_X10Y109_BO6),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_DO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h599aa665a665599a)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_CLUT (
.I0(CLBLM_R_X5Y106_SLICE_X6Y106_AO6),
.I1(CLBLM_R_X7Y108_SLICE_X8Y108_BO6),
.I2(CLBLM_R_X5Y109_SLICE_X6Y109_DO6),
.I3(CLBLL_L_X4Y108_SLICE_X4Y108_AO5),
.I4(CLBLM_R_X7Y108_SLICE_X9Y108_CO6),
.I5(CLBLM_R_X3Y109_SLICE_X3Y109_AO5),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_CO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000080000000)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_BLUT (
.I0(CLBLM_R_X5Y109_SLICE_X7Y109_BO6),
.I1(CLBLM_L_X8Y109_SLICE_X10Y109_BO6),
.I2(CLBLM_L_X10Y108_SLICE_X13Y108_BO6),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(CLBLM_R_X7Y106_SLICE_X9Y106_BO6),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_BO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h4bb4b44bd22d2dd2)
  ) CLBLM_R_X5Y108_SLICE_X7Y108_ALUT (
.I0(CLBLM_R_X5Y109_SLICE_X6Y109_DO6),
.I1(CLBLM_R_X7Y108_SLICE_X8Y108_BO6),
.I2(CLBLM_R_X5Y106_SLICE_X6Y106_AO6),
.I3(CLBLM_R_X7Y108_SLICE_X8Y108_AO6),
.I4(CLBLM_R_X7Y107_SLICE_X8Y107_AO6),
.I5(CLBLL_L_X4Y108_SLICE_X4Y108_AO5),
.O5(CLBLM_R_X5Y108_SLICE_X7Y108_AO5),
.O6(CLBLM_R_X5Y108_SLICE_X7Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0f4fdf4cdfffff)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_DLUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_DO6),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(CLBLM_R_X7Y109_SLICE_X8Y109_BO6),
.I4(CLBLM_R_X7Y109_SLICE_X9Y109_DO6),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_DO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h70f7f770f770f770)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_CLUT (
.I0(LIOB33_X0Y111_IOB_X0Y111_I),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(CLBLM_R_X5Y110_SLICE_X7Y110_BO6),
.I3(CLBLM_R_X7Y109_SLICE_X8Y109_AO6),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_CO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha66a66aa9a56965a)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_BLUT (
.I0(CLBLM_R_X5Y108_SLICE_X7Y108_AO6),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(CLBLM_R_X5Y108_SLICE_X6Y108_AO6),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(RIOB33_X105Y105_IOB_X1Y106_I),
.I5(CLBLM_R_X5Y109_SLICE_X6Y109_CO6),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_BO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha66599aa599a99aa)
  ) CLBLM_R_X5Y109_SLICE_X6Y109_ALUT (
.I0(CLBLM_R_X7Y109_SLICE_X9Y109_DO6),
.I1(CLBLM_R_X7Y110_SLICE_X8Y110_DO6),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(CLBLM_R_X7Y109_SLICE_X8Y109_BO6),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(LIOB33_X0Y109_IOB_X0Y110_I),
.O5(CLBLM_R_X5Y109_SLICE_X6Y109_AO5),
.O6(CLBLM_R_X5Y109_SLICE_X6Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000020000000000)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_DLUT (
.I0(CLBLM_R_X5Y109_SLICE_X7Y109_AO6),
.I1(CLBLM_R_X7Y103_SLICE_X9Y103_AO5),
.I2(CLBLL_L_X2Y111_SLICE_X0Y111_DO6),
.I3(RIOB33_SING_X105Y100_IOB_X1Y100_I),
.I4(CLBLM_R_X11Y106_SLICE_X15Y106_DO6),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_DO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0013005f00000000)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_CLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(RIOB33_X105Y103_IOB_X1Y103_I),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(CLBLM_R_X7Y103_SLICE_X9Y103_AO5),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(CLBLM_R_X3Y109_SLICE_X2Y109_BO6),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_CO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000100000000)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_BLUT (
.I0(CLBLL_L_X2Y111_SLICE_X0Y111_DO6),
.I1(CLBLM_R_X3Y109_SLICE_X2Y109_AO5),
.I2(CLBLM_R_X11Y106_SLICE_X15Y106_DO6),
.I3(CLBLM_R_X7Y112_SLICE_X8Y112_AO6),
.I4(CLBLM_L_X8Y112_SLICE_X10Y112_AO6),
.I5(CLBLM_R_X5Y109_SLICE_X7Y109_CO6),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_BO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h07007700f0f00000)
  ) CLBLM_R_X5Y109_SLICE_X7Y109_ALUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(CLBLM_R_X3Y109_SLICE_X2Y109_BO6),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y109_SLICE_X7Y109_AO5),
.O6(CLBLM_R_X5Y109_SLICE_X7Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc66699c66ccc336c)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_DLUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(CLBLM_R_X5Y110_SLICE_X7Y110_AO6),
.I2(RIOB33_X105Y105_IOB_X1Y106_I),
.I3(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_CO6),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_DO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdc4dc40f7317310)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_CLUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_AO6),
.I1(CLBLM_L_X8Y109_SLICE_X11Y109_AO5),
.I2(CLBLM_R_X5Y112_SLICE_X6Y112_AO5),
.I3(CLBLM_R_X7Y110_SLICE_X8Y110_AO6),
.I4(CLBLM_R_X7Y112_SLICE_X8Y112_AO6),
.I5(CLBLM_L_X8Y111_SLICE_X11Y111_AO6),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_CO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c33c69963cc396)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_BLUT (
.I0(CLBLM_R_X5Y112_SLICE_X6Y112_DO6),
.I1(CLBLM_L_X8Y110_SLICE_X11Y110_AO6),
.I2(CLBLM_R_X7Y110_SLICE_X9Y110_AO6),
.I3(CLBLM_R_X3Y112_SLICE_X3Y112_AO5),
.I4(CLBLM_R_X5Y110_SLICE_X6Y110_AO6),
.I5(CLBLM_R_X5Y110_SLICE_X6Y110_CO6),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_BO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h78871ee18778e11e)
  ) CLBLM_R_X5Y110_SLICE_X6Y110_ALUT (
.I0(CLBLM_R_X7Y112_SLICE_X8Y112_AO6),
.I1(CLBLM_R_X5Y112_SLICE_X6Y112_AO5),
.I2(CLBLM_R_X7Y110_SLICE_X8Y110_AO6),
.I3(CLBLM_L_X8Y109_SLICE_X11Y109_AO5),
.I4(CLBLM_L_X8Y112_SLICE_X10Y112_AO6),
.I5(CLBLM_L_X8Y111_SLICE_X11Y111_AO6),
.O5(CLBLM_R_X5Y110_SLICE_X6Y110_AO5),
.O6(CLBLM_R_X5Y110_SLICE_X6Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdc4dc40f7317310)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_DLUT (
.I0(CLBLM_R_X7Y110_SLICE_X8Y110_BO6),
.I1(CLBLM_R_X7Y110_SLICE_X9Y110_BO6),
.I2(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I3(CLBLL_L_X4Y103_SLICE_X5Y103_BO5),
.I4(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.I5(CLBLM_R_X7Y109_SLICE_X9Y109_AO6),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_DO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2bd4d42bd42b2bd4)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_CLUT (
.I0(CLBLM_R_X7Y110_SLICE_X8Y110_BO6),
.I1(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.I2(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I3(CLBLM_R_X7Y110_SLICE_X9Y110_BO6),
.I4(CLBLL_L_X4Y103_SLICE_X5Y103_BO5),
.I5(CLBLM_R_X7Y109_SLICE_X9Y109_AO6),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_CO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h33117f157f37ffff)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_BLUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_DO6),
.I1(RIOB33_X105Y105_IOB_X1Y106_I),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(CLBLM_R_X5Y111_SLICE_X6Y111_CO6),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLM_R_X5Y110_SLICE_X7Y110_CO6),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_BO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc639639c9999cccc)
  ) CLBLM_R_X5Y110_SLICE_X7Y110_ALUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I1(CLBLM_R_X7Y110_SLICE_X9Y110_BO6),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(CLBLM_R_X7Y110_SLICE_X8Y110_BO6),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLM_R_X5Y110_SLICE_X7Y110_AO5),
.O6(CLBLM_R_X5Y110_SLICE_X7Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a55a69965aa596)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_DLUT (
.I0(CLBLM_R_X5Y111_SLICE_X6Y111_AO6),
.I1(CLBLL_L_X4Y113_SLICE_X5Y113_BO6),
.I2(CLBLM_R_X5Y110_SLICE_X6Y110_BO6),
.I3(CLBLM_R_X5Y111_SLICE_X6Y111_AO5),
.I4(CLBLM_R_X5Y111_SLICE_X7Y111_CO6),
.I5(CLBLM_R_X3Y111_SLICE_X3Y111_BO6),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_DO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h60f6c0fcf6f6fcfc)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(CLBLM_R_X5Y111_SLICE_X7Y111_AO6),
.I2(CLBLL_L_X4Y113_SLICE_X5Y113_BO6),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_CO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hbd424db22dd2dd22)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_BLUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_CO6),
.I1(CLBLL_L_X4Y113_SLICE_X5Y113_BO6),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(CLBLM_R_X5Y110_SLICE_X6Y110_BO6),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(RIOB33_X105Y105_IOB_X1Y106_I),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_BO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff0fff0fff)
  ) CLBLM_R_X5Y111_SLICE_X6Y111_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(RIOB33_X105Y105_IOB_X1Y106_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y111_SLICE_X6Y111_AO5),
.O6(CLBLM_R_X5Y111_SLICE_X6Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1777ffff111755ff)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_DLUT (
.I0(CLBLM_R_X5Y110_SLICE_X6Y110_AO6),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_R_X7Y111_SLICE_X8Y111_AO5),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLM_R_X5Y112_SLICE_X7Y112_BO6),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_DO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9666aaaa999655aa)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_CLUT (
.I0(CLBLM_R_X5Y110_SLICE_X6Y110_AO6),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_R_X7Y111_SLICE_X8Y111_AO5),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(CLBLM_R_X5Y112_SLICE_X7Y112_BO6),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_CO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb73fc0b748c03f48)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_BLUT (
.I0(LIOB33_X0Y113_IOB_X0Y114_I),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(CLBLM_L_X8Y112_SLICE_X10Y112_AO6),
.I4(CLBLM_R_X7Y112_SLICE_X8Y112_AO6),
.I5(CLBLM_L_X8Y111_SLICE_X11Y111_AO6),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_BO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h9699aa556696aaaa)
  ) CLBLM_R_X5Y111_SLICE_X7Y111_ALUT (
.I0(CLBLM_R_X5Y111_SLICE_X7Y111_BO6),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(CLBLM_R_X5Y112_SLICE_X7Y112_BO6),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLM_R_X7Y111_SLICE_X8Y111_AO5),
.O5(CLBLM_R_X5Y111_SLICE_X7Y111_AO5),
.O6(CLBLM_R_X5Y111_SLICE_X7Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hecb38020fefbc832)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_DLUT (
.I0(CLBLM_R_X5Y112_SLICE_X6Y112_AO6),
.I1(CLBLM_R_X7Y112_SLICE_X9Y112_CO6),
.I2(CLBLL_L_X4Y112_SLICE_X5Y112_CO6),
.I3(CLBLM_R_X5Y112_SLICE_X6Y112_AO5),
.I4(CLBLL_L_X4Y112_SLICE_X5Y112_AO5),
.I5(CLBLM_R_X5Y112_SLICE_X6Y112_BO6),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_DO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93936c36c9c936)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_CLUT (
.I0(CLBLM_R_X5Y112_SLICE_X6Y112_AO6),
.I1(CLBLM_R_X7Y112_SLICE_X8Y112_AO6),
.I2(CLBLL_L_X4Y112_SLICE_X5Y112_CO6),
.I3(CLBLM_R_X5Y112_SLICE_X6Y112_AO5),
.I4(CLBLM_L_X8Y112_SLICE_X10Y112_AO6),
.I5(CLBLM_R_X5Y112_SLICE_X6Y112_BO6),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_CO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6a95956a95956a6a)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_BLUT (
.I0(CLBLM_R_X7Y111_SLICE_X9Y111_BO6),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(CLBLL_L_X4Y111_SLICE_X5Y111_CO6),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_BO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f5f5f5f0fff0fff)
  ) CLBLM_R_X5Y112_SLICE_X6Y112_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(1'b1),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X6Y112_AO5),
.O6(CLBLM_R_X5Y112_SLICE_X6Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_DO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_CO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h4cdfdf4cdfdf4c4c)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(CLBLL_L_X4Y112_SLICE_X5Y112_CO6),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(CLBLM_R_X5Y112_SLICE_X7Y112_AO6),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_BO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h965aaaaaa5966666)
  ) CLBLM_R_X5Y112_SLICE_X7Y112_ALUT (
.I0(CLBLM_R_X7Y111_SLICE_X9Y111_BO6),
.I1(CLBLM_R_X7Y107_SLICE_X9Y107_BO5),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLL_L_X4Y111_SLICE_X4Y111_AO5),
.O5(CLBLM_R_X5Y112_SLICE_X7Y112_AO5),
.O6(CLBLM_R_X5Y112_SLICE_X7Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y100_SLICE_X8Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y100_SLICE_X8Y100_DO5),
.O6(CLBLM_R_X7Y100_SLICE_X8Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc396699669c33c)
  ) CLBLM_R_X7Y100_SLICE_X8Y100_CLUT (
.I0(CLBLM_R_X7Y101_SLICE_X8Y101_AO6),
.I1(CLBLM_R_X7Y101_SLICE_X8Y101_AO5),
.I2(CLBLM_R_X7Y102_SLICE_X9Y102_DO6),
.I3(CLBLM_R_X7Y100_SLICE_X8Y100_AO5),
.I4(CLBLM_R_X7Y100_SLICE_X8Y100_BO5),
.I5(CLBLM_L_X8Y101_SLICE_X10Y101_AO6),
.O5(CLBLM_R_X7Y100_SLICE_X8Y100_CO5),
.O6(CLBLM_R_X7Y100_SLICE_X8Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f077f0777777777)
  ) CLBLM_R_X7Y100_SLICE_X8Y100_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(CLBLM_R_X7Y101_SLICE_X8Y101_AO6),
.I3(CLBLM_L_X8Y101_SLICE_X10Y101_AO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y100_SLICE_X8Y100_BO5),
.O6(CLBLM_R_X7Y100_SLICE_X8Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h699969990fff0fff)
  ) CLBLM_R_X7Y100_SLICE_X8Y100_ALUT (
.I0(CLBLM_R_X7Y102_SLICE_X9Y102_DO6),
.I1(CLBLM_R_X7Y101_SLICE_X8Y101_AO5),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y100_SLICE_X8Y100_AO5),
.O6(CLBLM_R_X7Y100_SLICE_X8Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y100_SLICE_X9Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y100_SLICE_X9Y100_DO5),
.O6(CLBLM_R_X7Y100_SLICE_X9Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y100_SLICE_X9Y100_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y100_SLICE_X9Y100_CO5),
.O6(CLBLM_R_X7Y100_SLICE_X9Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y100_SLICE_X9Y100_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y100_SLICE_X9Y100_BO5),
.O6(CLBLM_R_X7Y100_SLICE_X9Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y100_SLICE_X9Y100_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y100_SLICE_X9Y100_AO5),
.O6(CLBLM_R_X7Y100_SLICE_X9Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y101_SLICE_X8Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y101_SLICE_X8Y101_DO5),
.O6(CLBLM_R_X7Y101_SLICE_X8Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffffffcc333333)
  ) CLBLM_R_X7Y101_SLICE_X8Y101_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y100_SLICE_X8Y100_CO6),
.I2(1'b1),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y101_SLICE_X8Y101_CO5),
.O6(CLBLM_R_X7Y101_SLICE_X8Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h963c69c366cc9933)
  ) CLBLM_R_X7Y101_SLICE_X8Y101_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLM_L_X8Y101_SLICE_X10Y101_AO6),
.I2(CLBLM_L_X8Y103_SLICE_X10Y103_AO6),
.I3(RIOB33_X105Y107_IOB_X1Y107_I),
.I4(CLBLM_R_X7Y101_SLICE_X8Y101_AO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y101_SLICE_X8Y101_BO5),
.O6(CLBLM_R_X7Y101_SLICE_X8Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c369c371f371f3)
  ) CLBLM_R_X7Y101_SLICE_X8Y101_ALUT (
.I0(RIOB33_X105Y107_IOB_X1Y108_I),
.I1(CLBLM_R_X7Y103_SLICE_X8Y103_AO6),
.I2(CLBLM_R_X7Y101_SLICE_X9Y101_AO6),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y101_SLICE_X8Y101_AO5),
.O6(CLBLM_R_X7Y101_SLICE_X8Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y101_SLICE_X9Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y101_SLICE_X9Y101_DO5),
.O6(CLBLM_R_X7Y101_SLICE_X9Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00a25da200008888)
  ) CLBLM_R_X7Y101_SLICE_X9Y101_CLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(RIOB33_X105Y109_IOB_X1Y110_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(RIOB33_X105Y109_IOB_X1Y109_I),
.O5(CLBLM_R_X7Y101_SLICE_X9Y101_CO5),
.O6(CLBLM_R_X7Y101_SLICE_X9Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69a59955965a66aa)
  ) CLBLM_R_X7Y101_SLICE_X9Y101_BLUT (
.I0(CLBLM_L_X8Y103_SLICE_X10Y103_DO6),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(CLBLM_R_X7Y103_SLICE_X9Y103_AO5),
.O5(CLBLM_R_X7Y101_SLICE_X9Y101_BO5),
.O6(CLBLM_R_X7Y101_SLICE_X9Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2bafbbff8e0aeeaa)
  ) CLBLM_R_X7Y101_SLICE_X9Y101_ALUT (
.I0(CLBLM_L_X8Y103_SLICE_X10Y103_DO6),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(RIOB33_X105Y107_IOB_X1Y108_I),
.I5(CLBLM_R_X7Y103_SLICE_X9Y103_AO5),
.O5(CLBLM_R_X7Y101_SLICE_X9Y101_AO5),
.O6(CLBLM_R_X7Y101_SLICE_X9Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9c6c93936c6c9c6c)
  ) CLBLM_R_X7Y102_SLICE_X8Y102_DLUT (
.I0(RIOB33_X105Y107_IOB_X1Y107_I),
.I1(CLBLM_R_X7Y100_SLICE_X8Y100_CO6),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_L_X8Y103_SLICE_X10Y103_AO6),
.I5(CLBLM_R_X7Y101_SLICE_X8Y101_BO5),
.O5(CLBLM_R_X7Y102_SLICE_X8Y102_DO5),
.O6(CLBLM_R_X7Y102_SLICE_X8Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf88f8008feefe00e)
  ) CLBLM_R_X7Y102_SLICE_X8Y102_CLUT (
.I0(CLBLM_R_X7Y102_SLICE_X8Y102_AO6),
.I1(CLBLM_L_X8Y103_SLICE_X10Y103_AO6),
.I2(CLBLM_R_X7Y101_SLICE_X8Y101_CO6),
.I3(CLBLM_R_X7Y100_SLICE_X8Y100_CO6),
.I4(CLBLM_R_X7Y104_SLICE_X8Y104_BO5),
.I5(CLBLM_R_X7Y101_SLICE_X8Y101_BO5),
.O5(CLBLM_R_X7Y102_SLICE_X8Y102_CO5),
.O6(CLBLM_R_X7Y102_SLICE_X8Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h695aa56996a55a96)
  ) CLBLM_R_X7Y102_SLICE_X8Y102_BLUT (
.I0(CLBLM_R_X7Y104_SLICE_X8Y104_BO5),
.I1(CLBLM_L_X8Y103_SLICE_X10Y103_AO6),
.I2(CLBLM_R_X7Y101_SLICE_X8Y101_CO6),
.I3(CLBLM_R_X7Y101_SLICE_X8Y101_BO5),
.I4(CLBLM_R_X7Y102_SLICE_X8Y102_AO6),
.I5(CLBLM_R_X7Y100_SLICE_X8Y100_CO6),
.O5(CLBLM_R_X7Y102_SLICE_X8Y102_BO5),
.O6(CLBLM_R_X7Y102_SLICE_X8Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333ffff22bbaaff)
  ) CLBLM_R_X7Y102_SLICE_X8Y102_ALUT (
.I0(CLBLM_L_X8Y103_SLICE_X10Y103_AO6),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(1'b1),
.I3(CLBLM_R_X7Y101_SLICE_X8Y101_BO5),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y102_SLICE_X8Y102_AO5),
.O6(CLBLM_R_X7Y102_SLICE_X8Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h69969966c33c33cc)
  ) CLBLM_R_X7Y102_SLICE_X9Y102_DLUT (
.I0(RIOB33_X105Y109_IOB_X1Y109_I),
.I1(CLBLM_R_X5Y103_SLICE_X7Y103_AO6),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(CLBLM_R_X7Y103_SLICE_X8Y103_AO5),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_R_X7Y102_SLICE_X9Y102_DO5),
.O6(CLBLM_R_X7Y102_SLICE_X9Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6966996996996696)
  ) CLBLM_R_X7Y102_SLICE_X9Y102_CLUT (
.I0(CLBLM_R_X7Y103_SLICE_X9Y103_AO6),
.I1(CLBLM_L_X8Y104_SLICE_X10Y104_AO6),
.I2(CLBLL_L_X4Y103_SLICE_X4Y103_AO6),
.I3(CLBLM_L_X8Y103_SLICE_X10Y103_CO6),
.I4(CLBLM_R_X7Y102_SLICE_X9Y102_AO6),
.I5(CLBLM_R_X5Y102_SLICE_X7Y102_AO6),
.O5(CLBLM_R_X7Y102_SLICE_X9Y102_CO5),
.O6(CLBLM_R_X7Y102_SLICE_X9Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996699669696996)
  ) CLBLM_R_X7Y102_SLICE_X9Y102_BLUT (
.I0(CLBLM_L_X8Y102_SLICE_X10Y102_CO6),
.I1(CLBLL_L_X4Y102_SLICE_X4Y102_AO6),
.I2(CLBLM_R_X5Y101_SLICE_X6Y101_AO6),
.I3(CLBLM_R_X7Y101_SLICE_X9Y101_CO6),
.I4(CLBLM_R_X5Y101_SLICE_X7Y101_AO6),
.I5(CLBLM_L_X10Y101_SLICE_X13Y101_AO6),
.O5(CLBLM_R_X7Y102_SLICE_X9Y102_BO5),
.O6(CLBLM_R_X7Y102_SLICE_X9Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa5a500ffeda584)
  ) CLBLM_R_X7Y102_SLICE_X9Y102_ALUT (
.I0(CLBLM_L_X8Y102_SLICE_X10Y102_CO6),
.I1(CLBLM_R_X5Y101_SLICE_X7Y101_AO6),
.I2(CLBLM_R_X5Y101_SLICE_X6Y101_AO6),
.I3(CLBLM_R_X7Y101_SLICE_X9Y101_CO6),
.I4(CLBLL_L_X4Y102_SLICE_X4Y102_AO6),
.I5(CLBLM_L_X10Y101_SLICE_X13Y101_AO6),
.O5(CLBLM_R_X7Y102_SLICE_X9Y102_AO5),
.O6(CLBLM_R_X7Y102_SLICE_X9Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h48de88eededeeeee)
  ) CLBLM_R_X7Y103_SLICE_X8Y103_DLUT (
.I0(CLBLM_R_X7Y101_SLICE_X8Y101_BO6),
.I1(CLBLM_R_X7Y104_SLICE_X8Y104_CO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_R_X7Y103_SLICE_X8Y103_DO5),
.O6(CLBLM_R_X7Y103_SLICE_X8Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996996696966666)
  ) CLBLM_R_X7Y103_SLICE_X8Y103_CLUT (
.I0(CLBLM_R_X7Y101_SLICE_X8Y101_BO6),
.I1(CLBLM_R_X7Y104_SLICE_X8Y104_CO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_R_X7Y103_SLICE_X8Y103_CO5),
.O6(CLBLM_R_X7Y103_SLICE_X8Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h9aa6f30ca5aa0000)
  ) CLBLM_R_X7Y103_SLICE_X8Y103_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(CLBLM_R_X7Y105_SLICE_X8Y105_AO6),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(RIOB33_X105Y111_IOB_X1Y111_I),
.O5(CLBLM_R_X7Y103_SLICE_X8Y103_BO5),
.O6(CLBLM_R_X7Y103_SLICE_X8Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc3f00f30f3f0ff)
  ) CLBLM_R_X7Y103_SLICE_X8Y103_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(CLBLM_R_X7Y103_SLICE_X9Y103_CO6),
.I3(CLBLM_R_X7Y103_SLICE_X8Y103_BO6),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y103_SLICE_X8Y103_AO5),
.O6(CLBLM_R_X7Y103_SLICE_X8Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y103_SLICE_X9Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y103_SLICE_X9Y103_DO5),
.O6(CLBLM_R_X7Y103_SLICE_X9Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2abfbfbfbf2a2a2a)
  ) CLBLM_R_X7Y103_SLICE_X9Y103_CLUT (
.I0(CLBLM_L_X8Y104_SLICE_X10Y104_AO6),
.I1(RIOB33_X105Y109_IOB_X1Y109_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(RIOB33_X105Y109_IOB_X1Y110_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLM_R_X7Y103_SLICE_X9Y103_BO6),
.O5(CLBLM_R_X7Y103_SLICE_X9Y103_CO5),
.O6(CLBLM_R_X7Y103_SLICE_X9Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc73ff3ff33ff33ff)
  ) CLBLM_R_X7Y103_SLICE_X9Y103_BLUT (
.I0(RIOB33_X105Y111_IOB_X1Y112_I),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(RIOB33_X105Y111_IOB_X1Y111_I),
.I4(RIOB33_X105Y113_IOB_X1Y113_I),
.I5(RIOB33_X105Y109_IOB_X1Y110_I),
.O5(CLBLM_R_X7Y103_SLICE_X9Y103_BO5),
.O6(CLBLM_R_X7Y103_SLICE_X9Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc03fc03f3fc0c03f)
  ) CLBLM_R_X7Y103_SLICE_X9Y103_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(RIOB33_X105Y109_IOB_X1Y110_I),
.I3(CLBLM_R_X7Y103_SLICE_X9Y103_BO6),
.I4(CLBLM_L_X8Y104_SLICE_X10Y104_AO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y103_SLICE_X9Y103_AO5),
.O6(CLBLM_R_X7Y103_SLICE_X9Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h69969696a55a5a5a)
  ) CLBLM_R_X7Y104_SLICE_X8Y104_DLUT (
.I0(CLBLM_L_X8Y102_SLICE_X10Y102_BO6),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(CLBLM_L_X10Y103_SLICE_X12Y103_AO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_R_X7Y104_SLICE_X8Y104_DO5),
.O6(CLBLM_R_X7Y104_SLICE_X8Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h71b2b2b2f5fafafa)
  ) CLBLM_R_X7Y104_SLICE_X8Y104_CLUT (
.I0(CLBLM_L_X8Y102_SLICE_X10Y102_BO6),
.I1(LIOB33_X0Y107_IOB_X0Y108_I),
.I2(CLBLM_L_X10Y103_SLICE_X12Y103_AO6),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(RIOB33_X105Y103_IOB_X1Y104_I),
.O5(CLBLM_R_X7Y104_SLICE_X8Y104_CO5),
.O6(CLBLM_R_X7Y104_SLICE_X8Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff00ffffff)
  ) CLBLM_R_X7Y104_SLICE_X8Y104_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y104_SLICE_X8Y104_BO5),
.O6(CLBLM_R_X7Y104_SLICE_X8Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff55ff55ff)
  ) CLBLM_R_X7Y104_SLICE_X8Y104_ALUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(1'b1),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(RIOB33_X105Y103_IOB_X1Y104_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y104_SLICE_X8Y104_AO5),
.O6(CLBLM_R_X7Y104_SLICE_X8Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8778e11eff0033cc)
  ) CLBLM_R_X7Y104_SLICE_X9Y104_DLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(CLBLM_L_X8Y104_SLICE_X11Y104_BO6),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(CLBLM_L_X8Y104_SLICE_X10Y104_BO6),
.I4(CLBLM_L_X8Y105_SLICE_X10Y105_DO6),
.I5(LIOB33_X0Y109_IOB_X0Y109_I),
.O5(CLBLM_R_X7Y104_SLICE_X9Y104_DO5),
.O6(CLBLM_R_X7Y104_SLICE_X9Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a96a56996a5695a)
  ) CLBLM_R_X7Y104_SLICE_X9Y104_CLUT (
.I0(CLBLM_R_X7Y104_SLICE_X9Y104_AO6),
.I1(CLBLM_L_X10Y104_SLICE_X12Y104_CO6),
.I2(CLBLM_L_X10Y104_SLICE_X12Y104_BO6),
.I3(CLBLM_L_X8Y105_SLICE_X10Y105_AO5),
.I4(CLBLM_R_X7Y104_SLICE_X8Y104_AO6),
.I5(CLBLM_L_X10Y104_SLICE_X12Y104_AO6),
.O5(CLBLM_R_X7Y104_SLICE_X9Y104_CO5),
.O6(CLBLM_R_X7Y104_SLICE_X9Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f5f03137fff5f7f)
  ) CLBLM_R_X7Y104_SLICE_X9Y104_BLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(CLBLM_L_X8Y104_SLICE_X11Y104_BO6),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(CLBLM_L_X8Y105_SLICE_X10Y105_DO6),
.I5(CLBLM_R_X7Y104_SLICE_X9Y104_CO6),
.O5(CLBLM_R_X7Y104_SLICE_X9Y104_BO5),
.O6(CLBLM_R_X7Y104_SLICE_X9Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff3f03ff33)
  ) CLBLM_R_X7Y104_SLICE_X9Y104_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X7Y104_SLICE_X8Y104_DO6),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(CLBLM_L_X8Y104_SLICE_X11Y104_AO6),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y104_SLICE_X9Y104_AO5),
.O6(CLBLM_R_X7Y104_SLICE_X9Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y105_SLICE_X8Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y105_SLICE_X8Y105_DO5),
.O6(CLBLM_R_X7Y105_SLICE_X8Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y105_SLICE_X8Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y105_SLICE_X8Y105_CO5),
.O6(CLBLM_R_X7Y105_SLICE_X8Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y105_SLICE_X8Y105_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y105_SLICE_X8Y105_BO5),
.O6(CLBLM_R_X7Y105_SLICE_X8Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0d5fffff5fffffff)
  ) CLBLM_R_X7Y105_SLICE_X8Y105_ALUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(RIOB33_X105Y109_IOB_X1Y110_I),
.I5(RIOB33_X105Y111_IOB_X1Y111_I),
.O5(CLBLM_R_X7Y105_SLICE_X8Y105_AO5),
.O6(CLBLM_R_X7Y105_SLICE_X8Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y105_SLICE_X9Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y105_SLICE_X9Y105_DO5),
.O6(CLBLM_R_X7Y105_SLICE_X9Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y105_SLICE_X9Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y105_SLICE_X9Y105_CO5),
.O6(CLBLM_R_X7Y105_SLICE_X9Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y105_SLICE_X9Y105_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y105_SLICE_X9Y105_BO5),
.O6(CLBLM_R_X7Y105_SLICE_X9Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y105_SLICE_X9Y105_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y105_SLICE_X9Y105_AO5),
.O6(CLBLM_R_X7Y105_SLICE_X9Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y106_SLICE_X8Y106_DO5),
.O6(CLBLM_R_X7Y106_SLICE_X8Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y106_SLICE_X8Y106_CO5),
.O6(CLBLM_R_X7Y106_SLICE_X8Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y106_SLICE_X8Y106_BO5),
.O6(CLBLM_R_X7Y106_SLICE_X8Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y106_SLICE_X8Y106_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y106_SLICE_X8Y106_AO5),
.O6(CLBLM_R_X7Y106_SLICE_X8Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h39c69c63c639639c)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_DLUT (
.I0(CLBLM_L_X8Y106_SLICE_X10Y106_AO6),
.I1(CLBLM_R_X7Y104_SLICE_X9Y104_CO6),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_AO5),
.I3(CLBLM_R_X7Y106_SLICE_X9Y106_AO5),
.I4(CLBLM_L_X8Y106_SLICE_X11Y106_DO6),
.I5(CLBLM_L_X8Y106_SLICE_X10Y106_DO6),
.O5(CLBLM_R_X7Y106_SLICE_X9Y106_DO5),
.O6(CLBLM_R_X7Y106_SLICE_X9Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0b2b0bbb2fffbfff)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_CLUT (
.I0(CLBLM_L_X8Y106_SLICE_X10Y106_BO6),
.I1(CLBLM_L_X8Y105_SLICE_X10Y105_CO6),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(CLBLM_L_X8Y106_SLICE_X10Y106_AO6),
.O5(CLBLM_R_X7Y106_SLICE_X9Y106_CO5),
.O6(CLBLM_R_X7Y106_SLICE_X9Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd25ab49678f01e3c)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_BLUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(CLBLM_L_X8Y105_SLICE_X10Y105_CO6),
.I2(CLBLM_L_X8Y105_SLICE_X10Y105_BO6),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(CLBLM_L_X8Y106_SLICE_X10Y106_BO6),
.I5(RIOB33_X105Y101_IOB_X1Y102_I),
.O5(CLBLM_R_X7Y106_SLICE_X9Y106_BO5),
.O6(CLBLM_R_X7Y106_SLICE_X9Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff0f0fffff)
  ) CLBLM_R_X7Y106_SLICE_X9Y106_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y106_SLICE_X9Y106_AO5),
.O6(CLBLM_R_X7Y106_SLICE_X9Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y107_SLICE_X8Y107_DO5),
.O6(CLBLM_R_X7Y107_SLICE_X8Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1f5f7fff03135f7f)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_CLUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(CLBLM_R_X7Y107_SLICE_X9Y107_CO6),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(CLBLM_L_X8Y107_SLICE_X11Y107_BO6),
.I5(CLBLM_L_X8Y108_SLICE_X10Y108_BO6),
.O5(CLBLM_R_X7Y107_SLICE_X8Y107_CO5),
.O6(CLBLM_R_X7Y107_SLICE_X8Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h95aa6aaaa95a565a)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_BLUT (
.I0(CLBLM_L_X8Y107_SLICE_X11Y107_DO6),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_CO6),
.I3(LIOB33_X0Y109_IOB_X0Y109_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_L_X8Y108_SLICE_X10Y108_BO6),
.O5(CLBLM_R_X7Y107_SLICE_X8Y107_BO5),
.O6(CLBLM_R_X7Y107_SLICE_X8Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h93cc6cccc93c363c)
  ) CLBLM_R_X7Y107_SLICE_X8Y107_ALUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(CLBLM_L_X8Y107_SLICE_X11Y107_BO6),
.I2(CLBLM_R_X7Y107_SLICE_X9Y107_CO6),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLM_L_X8Y108_SLICE_X10Y108_BO6),
.O5(CLBLM_R_X7Y107_SLICE_X8Y107_AO5),
.O6(CLBLM_R_X7Y107_SLICE_X8Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h59a69a65a659659a)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_DLUT (
.I0(CLBLM_R_X7Y107_SLICE_X9Y107_AO6),
.I1(CLBLM_L_X8Y107_SLICE_X11Y107_BO6),
.I2(CLBLM_L_X8Y108_SLICE_X10Y108_CO6),
.I3(CLBLM_L_X8Y107_SLICE_X11Y107_CO6),
.I4(CLBLM_R_X7Y108_SLICE_X9Y108_BO5),
.I5(CLBLM_L_X8Y106_SLICE_X11Y106_AO6),
.O5(CLBLM_R_X7Y107_SLICE_X9Y107_DO5),
.O6(CLBLM_R_X7Y107_SLICE_X9Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69969696c33c3c3c)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_R_X11Y107_SLICE_X14Y107_BO6),
.I2(CLBLM_L_X10Y108_SLICE_X12Y108_AO6),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(RIOB33_X105Y101_IOB_X1Y101_I),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLM_R_X7Y107_SLICE_X9Y107_CO5),
.O6(CLBLM_R_X7Y107_SLICE_X9Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a55555cc333333)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_BLUT (
.I0(CLBLM_L_X8Y102_SLICE_X10Y102_CO6),
.I1(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I2(RIOB33_X105Y109_IOB_X1Y109_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y107_SLICE_X9Y107_BO5),
.O6(CLBLM_R_X7Y107_SLICE_X9Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff3f3f3f3f)
  ) CLBLM_R_X7Y107_SLICE_X9Y107_ALUT (
.I0(1'b1),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(1'b1),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y107_SLICE_X9Y107_AO5),
.O6(CLBLM_R_X7Y107_SLICE_X9Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_DO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd278b41e5af0963c)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_CLUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(CLBLM_L_X8Y109_SLICE_X10Y109_CO6),
.I2(CLBLM_L_X8Y108_SLICE_X10Y108_DO6),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(CLBLM_R_X7Y109_SLICE_X8Y109_DO6),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_CO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc399699969cc3ccc)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_BLUT (
.I0(CLBLM_R_X7Y109_SLICE_X8Y109_DO6),
.I1(CLBLM_L_X8Y108_SLICE_X10Y108_AO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(CLBLM_L_X8Y109_SLICE_X10Y109_CO6),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_BO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h03bb2bbb2bff3fff)
  ) CLBLM_R_X7Y108_SLICE_X8Y108_ALUT (
.I0(CLBLM_R_X7Y109_SLICE_X8Y109_DO6),
.I1(CLBLM_L_X8Y108_SLICE_X10Y108_AO6),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(CLBLM_L_X8Y109_SLICE_X10Y109_CO6),
.O5(CLBLM_R_X7Y108_SLICE_X8Y108_AO5),
.O6(CLBLM_R_X7Y108_SLICE_X8Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_DO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2dd2d22db44b4bb4)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_CLUT (
.I0(CLBLM_L_X8Y108_SLICE_X10Y108_AO6),
.I1(CLBLM_R_X7Y109_SLICE_X9Y109_CO6),
.I2(CLBLM_L_X8Y108_SLICE_X10Y108_CO6),
.I3(CLBLM_L_X8Y107_SLICE_X11Y107_BO6),
.I4(CLBLM_R_X7Y108_SLICE_X9Y108_BO5),
.I5(CLBLM_R_X7Y108_SLICE_X9Y108_BO6),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_CO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fff0fff3f3f3f3f)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_X0Y109_IOB_X0Y110_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_BO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3f3f3f3f0fff0fff)
  ) CLBLM_R_X7Y108_SLICE_X9Y108_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y115_IOB_X0Y116_I),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y108_SLICE_X9Y108_AO5),
.O6(CLBLM_R_X7Y108_SLICE_X9Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff07778fff0888)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_DLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I5(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_DO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6696969999696966)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_CLUT (
.I0(CLBLM_L_X8Y108_SLICE_X10Y108_AO6),
.I1(CLBLM_R_X7Y109_SLICE_X9Y109_CO6),
.I2(CLBLM_R_X7Y109_SLICE_X9Y109_DO6),
.I3(CLBLM_R_X5Y110_SLICE_X7Y110_DO6),
.I4(CLBLM_R_X3Y110_SLICE_X3Y110_AO5),
.I5(CLBLM_R_X7Y108_SLICE_X9Y108_BO6),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_CO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h6999a55596665aaa)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_BLUT (
.I0(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I1(LIOB33_X0Y107_IOB_X0Y107_I),
.I2(LIOB33_X0Y107_IOB_X0Y108_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLM_L_X8Y111_SLICE_X11Y111_CO6),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_BO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc96c399c693c99cc)
  ) CLBLM_R_X7Y109_SLICE_X8Y109_ALUT (
.I0(CLBLM_R_X7Y110_SLICE_X8Y110_DO6),
.I1(CLBLM_R_X7Y109_SLICE_X9Y109_BO6),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(CLBLM_R_X7Y109_SLICE_X8Y109_BO6),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(LIOB33_X0Y103_IOB_X0Y103_I),
.O5(CLBLM_R_X7Y109_SLICE_X8Y109_AO5),
.O6(CLBLM_R_X7Y109_SLICE_X8Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93936c36c9c936)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_DLUT (
.I0(CLBLM_R_X7Y109_SLICE_X9Y109_AO6),
.I1(CLBLM_L_X8Y109_SLICE_X11Y109_BO6),
.I2(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I3(CLBLM_R_X7Y109_SLICE_X9Y109_AO5),
.I4(CLBLM_R_X7Y108_SLICE_X9Y108_AO5),
.I5(CLBLM_L_X8Y109_SLICE_X10Y109_AO6),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_DO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hecb38020fefbc832)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_CLUT (
.I0(CLBLM_R_X7Y109_SLICE_X9Y109_AO6),
.I1(CLBLM_L_X8Y109_SLICE_X11Y109_BO6),
.I2(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I3(CLBLM_R_X7Y109_SLICE_X9Y109_AO5),
.I4(CLBLM_R_X7Y108_SLICE_X9Y108_AO5),
.I5(CLBLM_L_X8Y109_SLICE_X10Y109_AO6),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_CO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd5b97f132a4680ec)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(CLBLM_L_X8Y109_SLICE_X10Y109_AO6),
.I2(LIOB33_X0Y113_IOB_X0Y114_I),
.I3(CLBLM_R_X7Y110_SLICE_X8Y110_CO6),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLM_L_X8Y109_SLICE_X11Y109_BO6),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_BO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff00ffffff)
  ) CLBLM_R_X7Y109_SLICE_X9Y109_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(1'b1),
.I3(LIOB33_X0Y107_IOB_X0Y108_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(1'b1),
.O5(CLBLM_R_X7Y109_SLICE_X9Y109_AO5),
.O6(CLBLM_R_X7Y109_SLICE_X9Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h70f7f770f7f77070)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_DLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(CLBLM_R_X7Y111_SLICE_X8Y111_CO6),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_DO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h48dec0fcdedefcfc)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_CLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(CLBLM_R_X5Y110_SLICE_X6Y110_CO6),
.I2(CLBLM_L_X8Y110_SLICE_X11Y110_BO6),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_CO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887878787787878)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(CLBLM_L_X8Y110_SLICE_X11Y110_BO6),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLM_R_X5Y110_SLICE_X6Y110_CO6),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_BO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff0fff0fff)
  ) CLBLM_R_X7Y110_SLICE_X8Y110_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y110_SLICE_X8Y110_AO5),
.O6(CLBLM_R_X7Y110_SLICE_X8Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_DO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_CO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h59a69a65a659659a)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_BLUT (
.I0(CLBLM_L_X8Y110_SLICE_X11Y110_CO6),
.I1(CLBLM_L_X8Y110_SLICE_X11Y110_AO6),
.I2(CLBLM_R_X5Y110_SLICE_X6Y110_CO6),
.I3(CLBLM_L_X10Y110_SLICE_X12Y110_AO6),
.I4(CLBLM_R_X7Y110_SLICE_X9Y110_AO6),
.I5(CLBLM_R_X7Y110_SLICE_X9Y110_AO5),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_BO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h777777775f5f5f5f)
  ) CLBLM_R_X7Y110_SLICE_X9Y110_ALUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y110_SLICE_X9Y110_AO5),
.O6(CLBLM_R_X7Y110_SLICE_X9Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996a55a96965a5a)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_DLUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_CO6),
.I1(LIOB33_X0Y103_IOB_X0Y103_I),
.I2(CLBLM_R_X5Y111_SLICE_X7Y111_DO6),
.I3(LIOB33_X0Y107_IOB_X0Y107_I),
.I4(LIOB33_X0Y107_IOB_X0Y108_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_DO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdb242bd44bb4bb44)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_CLUT (
.I0(CLBLM_R_X7Y111_SLICE_X8Y111_AO6),
.I1(CLBLM_L_X8Y111_SLICE_X10Y111_DO6),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_L_X8Y110_SLICE_X11Y110_BO6),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(LIOB33_X0Y113_IOB_X0Y114_I),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_CO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h47650ff000aaaa00)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_BLUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y115_IOB_X0Y116_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(RIOB33_X105Y113_IOB_X1Y113_I),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_BO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h77ff115566aa9955)
  ) CLBLM_R_X7Y111_SLICE_X8Y111_ALUT (
.I0(CLBLM_L_X8Y112_SLICE_X10Y112_AO6),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(1'b1),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(CLBLM_R_X7Y112_SLICE_X8Y112_AO6),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X8Y111_AO5),
.O6(CLBLM_R_X7Y111_SLICE_X8Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_DO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_CO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aaaa5665aaa9666)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_BLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_BO6),
.I1(CLBLM_R_X7Y111_SLICE_X8Y111_BO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(CLBLM_R_X7Y111_SLICE_X9Y111_AO6),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_BO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h404000406c60ac60)
  ) CLBLM_R_X7Y111_SLICE_X9Y111_ALUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(RIOB33_X105Y113_IOB_X1Y113_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(RIOB33_X105Y101_IOB_X1Y101_I),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(LIOB33_X0Y115_IOB_X0Y116_I),
.O5(CLBLM_R_X7Y111_SLICE_X9Y111_AO5),
.O6(CLBLM_R_X7Y111_SLICE_X9Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_DO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_CO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_BO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6cff006cffff6c6c)
  ) CLBLM_R_X7Y112_SLICE_X8Y112_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(CLBLM_R_X7Y111_SLICE_X9Y111_BO6),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(CLBLL_L_X4Y111_SLICE_X5Y111_CO6),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_R_X7Y112_SLICE_X8Y112_AO5),
.O6(CLBLM_R_X7Y112_SLICE_X8Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_DO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h78871ee18778e11e)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_CLUT (
.I0(CLBLM_R_X7Y112_SLICE_X9Y112_AO6),
.I1(CLBLL_L_X4Y111_SLICE_X5Y111_CO6),
.I2(CLBLM_L_X8Y112_SLICE_X11Y112_DO6),
.I3(CLBLM_R_X7Y112_SLICE_X9Y112_AO5),
.I4(CLBLM_L_X8Y111_SLICE_X10Y111_BO6),
.I5(CLBLM_L_X8Y111_SLICE_X10Y111_CO6),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_CO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h16348aa81eb402a8)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_BLUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_BO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33ff33ff3f3f3f3f)
  ) CLBLM_R_X7Y112_SLICE_X9Y112_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X7Y112_SLICE_X9Y112_AO5),
.O6(CLBLM_R_X7Y112_SLICE_X9Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y103_SLICE_X14Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y103_SLICE_X14Y103_DO5),
.O6(CLBLM_R_X11Y103_SLICE_X14Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y103_SLICE_X14Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y103_SLICE_X14Y103_CO5),
.O6(CLBLM_R_X11Y103_SLICE_X14Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffbf3f153f2a00)
  ) CLBLM_R_X11Y103_SLICE_X14Y103_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y104_SLICE_X15Y104_DO6),
.I5(CLBLM_R_X11Y104_SLICE_X15Y104_CO6),
.O5(CLBLM_R_X11Y103_SLICE_X14Y103_BO5),
.O6(CLBLM_R_X11Y103_SLICE_X14Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h2b8eaf0abbeeffaa)
  ) CLBLM_R_X11Y103_SLICE_X14Y103_ALUT (
.I0(CLBLM_R_X11Y104_SLICE_X14Y104_DO6),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(CLBLM_L_X10Y103_SLICE_X13Y103_CO6),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y103_SLICE_X14Y103_AO5),
.O6(CLBLM_R_X11Y103_SLICE_X14Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y103_SLICE_X15Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y103_SLICE_X15Y103_DO5),
.O6(CLBLM_R_X11Y103_SLICE_X15Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y103_SLICE_X15Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y103_SLICE_X15Y103_CO5),
.O6(CLBLM_R_X11Y103_SLICE_X15Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y103_SLICE_X15Y103_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y103_SLICE_X15Y103_BO5),
.O6(CLBLM_R_X11Y103_SLICE_X15Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y103_SLICE_X15Y103_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y103_SLICE_X15Y103_AO5),
.O6(CLBLM_R_X11Y103_SLICE_X15Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfccffccfd44dc00c)
  ) CLBLM_R_X11Y104_SLICE_X14Y104_DLUT (
.I0(CLBLM_R_X11Y105_SLICE_X15Y105_AO6),
.I1(CLBLM_R_X11Y104_SLICE_X15Y104_AO5),
.I2(CLBLL_L_X4Y103_SLICE_X4Y103_BO6),
.I3(CLBLM_L_X12Y104_SLICE_X16Y104_BO6),
.I4(CLBLM_R_X11Y104_SLICE_X15Y104_AO6),
.I5(CLBLM_L_X12Y104_SLICE_X16Y104_CO6),
.O5(CLBLM_R_X11Y104_SLICE_X14Y104_DO5),
.O6(CLBLM_R_X11Y104_SLICE_X14Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3cc33cc39669c33c)
  ) CLBLM_R_X11Y104_SLICE_X14Y104_CLUT (
.I0(CLBLM_R_X11Y105_SLICE_X15Y105_AO6),
.I1(CLBLM_R_X11Y104_SLICE_X15Y104_AO5),
.I2(CLBLL_L_X4Y103_SLICE_X4Y103_BO6),
.I3(CLBLM_L_X12Y104_SLICE_X16Y104_BO6),
.I4(CLBLM_R_X11Y104_SLICE_X15Y104_AO6),
.I5(CLBLM_L_X12Y104_SLICE_X16Y104_CO6),
.O5(CLBLM_R_X11Y104_SLICE_X14Y104_CO5),
.O6(CLBLM_R_X11Y104_SLICE_X14Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h69969966a55a55aa)
  ) CLBLM_R_X11Y104_SLICE_X14Y104_BLUT (
.I0(CLBLM_R_X11Y104_SLICE_X14Y104_DO6),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_L_X10Y103_SLICE_X13Y103_CO6),
.I4(LIOB33_X0Y103_IOB_X0Y104_I),
.I5(LIOB33_X0Y101_IOB_X0Y102_I),
.O5(CLBLM_R_X11Y104_SLICE_X14Y104_BO5),
.O6(CLBLM_R_X11Y104_SLICE_X14Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h6c93936c936c936c)
  ) CLBLM_R_X11Y104_SLICE_X14Y104_ALUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(CLBLM_R_X11Y104_SLICE_X15Y104_DO6),
.I2(RIOB33_X105Y105_IOB_X1Y105_I),
.I3(CLBLM_R_X11Y104_SLICE_X15Y104_CO6),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_R_X11Y104_SLICE_X14Y104_AO5),
.O6(CLBLM_R_X11Y104_SLICE_X14Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h9c3cc39c6ccc336c)
  ) CLBLM_R_X11Y104_SLICE_X15Y104_DLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(CLBLM_L_X10Y103_SLICE_X13Y103_CO6),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(CLBLM_L_X10Y103_SLICE_X13Y103_AO6),
.I4(CLBLM_R_X11Y104_SLICE_X15Y104_BO5),
.I5(RIOB33_X105Y107_IOB_X1Y107_I),
.O5(CLBLM_R_X11Y104_SLICE_X15Y104_DO5),
.O6(CLBLM_R_X11Y104_SLICE_X15Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h70f7f7f780f8f8f8)
  ) CLBLM_R_X11Y104_SLICE_X15Y104_CLUT (
.I0(RIOB33_X105Y105_IOB_X1Y105_I),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(CLBLM_L_X10Y106_SLICE_X12Y106_CO6),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(CLBLM_L_X12Y104_SLICE_X16Y104_AO6),
.O5(CLBLM_R_X11Y104_SLICE_X15Y104_CO5),
.O6(CLBLM_R_X11Y104_SLICE_X15Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0000fffcccccfff)
  ) CLBLM_R_X11Y104_SLICE_X15Y104_BLUT (
.I0(1'b1),
.I1(CLBLM_L_X12Y104_SLICE_X16Y104_CO6),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(CLBLM_R_X11Y105_SLICE_X15Y105_AO6),
.I5(1'b1),
.O5(CLBLM_R_X11Y104_SLICE_X15Y104_BO5),
.O6(CLBLM_R_X11Y104_SLICE_X15Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fffff3333ffff)
  ) CLBLM_R_X11Y104_SLICE_X15Y104_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(1'b1),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y104_SLICE_X15Y104_AO5),
.O6(CLBLM_R_X11Y104_SLICE_X15Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h965aa596aaaa6666)
  ) CLBLM_R_X11Y105_SLICE_X14Y105_DLUT (
.I0(CLBLM_L_X10Y104_SLICE_X13Y104_DO6),
.I1(CLBLM_R_X11Y105_SLICE_X15Y105_CO6),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(CLBLM_R_X11Y106_SLICE_X15Y106_DO6),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_R_X11Y105_SLICE_X14Y105_DO5),
.O6(CLBLM_R_X11Y105_SLICE_X14Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4bb4d22db44b2dd2)
  ) CLBLM_R_X11Y105_SLICE_X14Y105_CLUT (
.I0(CLBLM_R_X11Y105_SLICE_X14Y105_AO6),
.I1(CLBLM_R_X11Y105_SLICE_X15Y105_CO6),
.I2(CLBLM_L_X10Y104_SLICE_X13Y104_DO6),
.I3(CLBLM_R_X11Y105_SLICE_X14Y105_AO5),
.I4(CLBLM_R_X11Y106_SLICE_X15Y106_DO6),
.I5(CLBLM_L_X10Y105_SLICE_X13Y105_AO6),
.O5(CLBLM_R_X11Y105_SLICE_X14Y105_CO5),
.O6(CLBLM_R_X11Y105_SLICE_X14Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hefbfce3b8c230802)
  ) CLBLM_R_X11Y105_SLICE_X14Y105_BLUT (
.I0(CLBLM_R_X11Y106_SLICE_X15Y106_DO6),
.I1(CLBLM_L_X10Y104_SLICE_X13Y104_DO6),
.I2(CLBLM_R_X11Y105_SLICE_X15Y105_CO6),
.I3(CLBLM_L_X10Y105_SLICE_X13Y105_AO6),
.I4(CLBLM_R_X11Y105_SLICE_X14Y105_AO6),
.I5(CLBLM_R_X11Y105_SLICE_X14Y105_AO5),
.O5(CLBLM_R_X11Y105_SLICE_X14Y105_BO5),
.O6(CLBLM_R_X11Y105_SLICE_X14Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffffff0fff0fff)
  ) CLBLM_R_X11Y105_SLICE_X14Y105_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(LIOB33_X0Y105_IOB_X0Y105_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y105_SLICE_X14Y105_AO5),
.O6(CLBLM_R_X11Y105_SLICE_X14Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha6996a5566a6aa6a)
  ) CLBLM_R_X11Y105_SLICE_X15Y105_DLUT (
.I0(CLBLM_L_X12Y104_SLICE_X16Y104_AO6),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(CLBLM_R_X11Y106_SLICE_X15Y106_AO5),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_R_X11Y104_SLICE_X15Y104_BO6),
.O5(CLBLM_R_X11Y105_SLICE_X15Y105_DO5),
.O6(CLBLM_R_X11Y105_SLICE_X15Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h7887878787787878)
  ) CLBLM_R_X11Y105_SLICE_X15Y105_CLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(CLBLM_L_X10Y106_SLICE_X12Y106_CO6),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(RIOB33_X105Y105_IOB_X1Y105_I),
.I5(CLBLM_L_X12Y104_SLICE_X16Y104_AO6),
.O5(CLBLM_R_X11Y105_SLICE_X15Y105_CO5),
.O6(CLBLM_R_X11Y105_SLICE_X15Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0455f30044004400)
  ) CLBLM_R_X11Y105_SLICE_X15Y105_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y105_SLICE_X15Y105_BO5),
.O6(CLBLM_R_X11Y105_SLICE_X15Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h113b80aa6e44a288)
  ) CLBLM_R_X11Y105_SLICE_X15Y105_ALUT (
.I0(RIOB33_X105Y113_IOB_X1Y113_I),
.I1(RIOB33_X105Y107_IOB_X1Y107_I),
.I2(RIOB33_X105Y111_IOB_X1Y112_I),
.I3(RIOB33_X105Y107_IOB_X1Y108_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y105_SLICE_X15Y105_AO5),
.O6(CLBLM_R_X11Y105_SLICE_X15Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h669c639c999c9c9c)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_DLUT (
.I0(CLBLM_R_X11Y105_SLICE_X15Y105_BO6),
.I1(CLBLM_R_X11Y105_SLICE_X15Y105_AO6),
.I2(CLBLM_R_X11Y106_SLICE_X15Y106_BO6),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(RIOB33_X105Y105_IOB_X1Y105_I),
.O5(CLBLM_R_X11Y106_SLICE_X14Y106_DO5),
.O6(CLBLM_R_X11Y106_SLICE_X14Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hd7b1284e5f93a06c)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_CLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(CLBLM_R_X11Y106_SLICE_X15Y106_AO6),
.I2(RIOB33_X105Y103_IOB_X1Y104_I),
.I3(CLBLM_R_X11Y107_SLICE_X14Y107_AO5),
.I4(CLBLM_R_X11Y106_SLICE_X14Y106_DO6),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_R_X11Y106_SLICE_X14Y106_CO5),
.O6(CLBLM_R_X11Y106_SLICE_X14Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f13ff5fb320ffa0)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y104_I),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(CLBLM_R_X11Y108_SLICE_X15Y108_BO6),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(CLBLM_R_X11Y106_SLICE_X14Y106_CO6),
.O5(CLBLM_R_X11Y106_SLICE_X14Y106_BO5),
.O6(CLBLM_R_X11Y106_SLICE_X14Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h07708dfa5a5a0000)
  ) CLBLM_R_X11Y106_SLICE_X14Y106_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(RIOB33_X105Y105_IOB_X1Y105_I),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(RIOB33_X105Y113_IOB_X1Y113_I),
.O5(CLBLM_R_X11Y106_SLICE_X14Y106_AO5),
.O6(CLBLM_R_X11Y106_SLICE_X14Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7b12f330ff5afff0)
  ) CLBLM_R_X11Y106_SLICE_X15Y106_DLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(CLBLM_R_X11Y106_SLICE_X14Y106_DO6),
.I3(CLBLM_L_X10Y107_SLICE_X13Y107_CO6),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_R_X11Y106_SLICE_X15Y106_DO5),
.O6(CLBLM_R_X11Y106_SLICE_X15Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996a55ac33c0ff0)
  ) CLBLM_R_X11Y106_SLICE_X15Y106_CLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(CLBLM_R_X11Y106_SLICE_X14Y106_DO6),
.I3(CLBLM_L_X10Y107_SLICE_X13Y107_CO6),
.I4(RIOB33_X105Y103_IOB_X1Y104_I),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_R_X11Y106_SLICE_X15Y106_CO5),
.O6(CLBLM_R_X11Y106_SLICE_X15Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h1d602e605160ae60)
  ) CLBLM_R_X11Y106_SLICE_X15Y106_BLUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(RIOB33_X105Y105_IOB_X1Y105_I),
.I2(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(RIOB33_X105Y107_IOB_X1Y107_I),
.I5(RIOB33_X105Y111_IOB_X1Y112_I),
.O5(CLBLM_R_X11Y106_SLICE_X15Y106_BO5),
.O6(CLBLM_R_X11Y106_SLICE_X15Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88778877f0f7f0f7)
  ) CLBLM_R_X11Y106_SLICE_X15Y106_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(CLBLM_R_X11Y105_SLICE_X15Y105_BO6),
.I3(CLBLM_R_X11Y106_SLICE_X15Y106_BO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y106_SLICE_X15Y106_AO5),
.O6(CLBLM_R_X11Y106_SLICE_X15Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3fc03f9fc03fc060)
  ) CLBLM_R_X11Y107_SLICE_X14Y107_DLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(RIOB33_X105Y103_IOB_X1Y104_I),
.I2(LIOB33_X0Y101_IOB_X0Y101_I),
.I3(CLBLM_L_X10Y107_SLICE_X13Y107_BO6),
.I4(CLBLM_R_X11Y106_SLICE_X14Y106_AO6),
.I5(CLBLM_R_X11Y106_SLICE_X15Y106_BO6),
.O5(CLBLM_R_X11Y107_SLICE_X14Y107_DO5),
.O6(CLBLM_R_X11Y107_SLICE_X14Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c39933963c66cc)
  ) CLBLM_R_X11Y107_SLICE_X14Y107_CLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(CLBLM_R_X11Y106_SLICE_X14Y106_CO6),
.I2(LIOB33_X0Y105_IOB_X0Y105_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(CLBLM_R_X11Y108_SLICE_X15Y108_BO6),
.O5(CLBLM_R_X11Y107_SLICE_X14Y107_CO5),
.O6(CLBLM_R_X11Y107_SLICE_X14Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd2a5780f5ad2f078)
  ) CLBLM_R_X11Y107_SLICE_X14Y107_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(CLBLM_R_X11Y107_SLICE_X15Y107_CO6),
.I3(CLBLM_R_X11Y108_SLICE_X14Y108_AO6),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(CLBLM_R_X11Y107_SLICE_X14Y107_CO6),
.O5(CLBLM_R_X11Y107_SLICE_X14Y107_BO5),
.O6(CLBLM_R_X11Y107_SLICE_X14Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'ha5a50f0fcdcdcfcf)
  ) CLBLM_R_X11Y107_SLICE_X14Y107_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y101_I),
.I1(CLBLM_L_X10Y107_SLICE_X13Y107_BO6),
.I2(CLBLM_R_X11Y106_SLICE_X14Y106_AO6),
.I3(1'b1),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y107_SLICE_X14Y107_AO5),
.O6(CLBLM_R_X11Y107_SLICE_X14Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3963c3c69c396)
  ) CLBLM_R_X11Y107_SLICE_X15Y107_DLUT (
.I0(CLBLM_R_X11Y107_SLICE_X15Y107_AO6),
.I1(CLBLM_R_X11Y105_SLICE_X14Y105_AO6),
.I2(CLBLM_L_X10Y109_SLICE_X13Y109_AO5),
.I3(CLBLM_R_X11Y108_SLICE_X15Y108_BO6),
.I4(CLBLM_L_X10Y106_SLICE_X13Y106_AO6),
.I5(CLBLM_R_X11Y106_SLICE_X15Y106_CO6),
.O5(CLBLM_R_X11Y107_SLICE_X15Y107_DO5),
.O6(CLBLM_R_X11Y107_SLICE_X15Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h6996c33c3cc36996)
  ) CLBLM_R_X11Y107_SLICE_X15Y107_CLUT (
.I0(CLBLM_R_X11Y107_SLICE_X15Y107_AO6),
.I1(CLBLM_R_X11Y105_SLICE_X14Y105_AO6),
.I2(CLBLM_R_X11Y106_SLICE_X15Y106_DO6),
.I3(CLBLM_R_X11Y105_SLICE_X15Y105_CO6),
.I4(CLBLM_R_X11Y108_SLICE_X15Y108_BO6),
.I5(CLBLM_R_X11Y106_SLICE_X15Y106_CO6),
.O5(CLBLM_R_X11Y107_SLICE_X15Y107_CO5),
.O6(CLBLM_R_X11Y107_SLICE_X15Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hedffa5ed84a50084)
  ) CLBLM_R_X11Y107_SLICE_X15Y107_BLUT (
.I0(CLBLM_L_X10Y106_SLICE_X13Y106_AO6),
.I1(CLBLM_R_X11Y108_SLICE_X15Y108_BO6),
.I2(CLBLM_R_X11Y105_SLICE_X14Y105_AO6),
.I3(CLBLM_R_X11Y106_SLICE_X15Y106_CO6),
.I4(CLBLM_R_X11Y107_SLICE_X15Y107_AO6),
.I5(CLBLM_L_X10Y109_SLICE_X13Y109_AO5),
.O5(CLBLM_R_X11Y107_SLICE_X15Y107_BO5),
.O6(CLBLM_R_X11Y107_SLICE_X15Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffffff0f0fffff)
  ) CLBLM_R_X11Y107_SLICE_X15Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y103_IOB_X0Y104_I),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(1'b1),
.O5(CLBLM_R_X11Y107_SLICE_X15Y107_AO5),
.O6(CLBLM_R_X11Y107_SLICE_X15Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb42ddddd4bd22222)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_DLUT (
.I0(CLBLM_R_X11Y107_SLICE_X14Y107_AO6),
.I1(CLBLM_R_X11Y109_SLICE_X14Y109_AO5),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLM_R_X11Y107_SLICE_X14Y107_DO6),
.O5(CLBLM_R_X11Y108_SLICE_X14Y108_DO5),
.O6(CLBLM_R_X11Y108_SLICE_X14Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3963ca50f5af0)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(CLBLM_R_X11Y109_SLICE_X14Y109_BO6),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLM_R_X11Y108_SLICE_X14Y108_DO6),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLM_R_X11Y108_SLICE_X14Y108_CO5),
.O6(CLBLM_R_X11Y108_SLICE_X14Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h93cc6cccc93c363c)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_BLUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(CLBLM_L_X10Y108_SLICE_X13Y108_CO6),
.I2(CLBLM_R_X11Y108_SLICE_X15Y108_CO6),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(CLBLM_R_X11Y109_SLICE_X14Y109_BO6),
.O5(CLBLM_R_X11Y108_SLICE_X14Y108_BO5),
.O6(CLBLM_R_X11Y108_SLICE_X14Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7dfff5ff143c50f0)
  ) CLBLM_R_X11Y108_SLICE_X14Y108_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(LIOB33_X0Y103_IOB_X0Y104_I),
.I2(CLBLM_R_X11Y108_SLICE_X14Y108_DO6),
.I3(LIOB33_X0Y105_IOB_X0Y105_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(CLBLM_R_X11Y109_SLICE_X14Y109_BO6),
.O5(CLBLM_R_X11Y108_SLICE_X14Y108_AO5),
.O6(CLBLM_R_X11Y108_SLICE_X14Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y108_SLICE_X15Y108_DO5),
.O6(CLBLM_R_X11Y108_SLICE_X15Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h69c3963c993366cc)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_CLUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(CLBLM_R_X11Y107_SLICE_X14Y107_DO6),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(CLBLM_L_X10Y109_SLICE_X13Y109_DO6),
.I5(RIOB33_X105Y103_IOB_X1Y103_I),
.O5(CLBLM_R_X11Y108_SLICE_X15Y108_CO5),
.O6(CLBLM_R_X11Y108_SLICE_X15Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2b8e8e8ebbeeeeee)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_BLUT (
.I0(CLBLM_L_X10Y109_SLICE_X13Y109_DO6),
.I1(CLBLM_R_X11Y107_SLICE_X14Y107_DO6),
.I2(RIOB33_X105Y101_IOB_X1Y102_I),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(RIOB33_X105Y103_IOB_X1Y103_I),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_R_X11Y108_SLICE_X15Y108_BO5),
.O6(CLBLM_R_X11Y108_SLICE_X15Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00002fa0d000d0a0)
  ) CLBLM_R_X11Y108_SLICE_X15Y108_ALUT (
.I0(RIOB33_X105Y103_IOB_X1Y104_I),
.I1(RIOB33_X105Y111_IOB_X1Y112_I),
.I2(RIOB33_X105Y113_IOB_X1Y113_I),
.I3(RIOB33_X105Y103_IOB_X1Y103_I),
.I4(RIOB33_X105Y101_IOB_X1Y102_I),
.I5(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O5(CLBLM_R_X11Y108_SLICE_X15Y108_AO5),
.O6(CLBLM_R_X11Y108_SLICE_X15Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y109_SLICE_X14Y109_DO5),
.O6(CLBLM_R_X11Y109_SLICE_X14Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55a9aa56ff0f00f0)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_CLUT (
.I0(RIOB33_X105Y103_IOB_X1Y103_I),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I3(CLBLM_R_X11Y108_SLICE_X15Y108_AO6),
.I4(CLBLM_R_X11Y106_SLICE_X14Y106_AO6),
.I5(LIOB33_X0Y101_IOB_X0Y101_I),
.O5(CLBLM_R_X11Y109_SLICE_X14Y109_CO5),
.O6(CLBLM_R_X11Y109_SLICE_X14Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2bbbafff8eee0aaa)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_BLUT (
.I0(CLBLM_L_X10Y110_SLICE_X13Y110_DO6),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(RIOB33_X105Y101_IOB_X1Y101_I),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLM_R_X11Y109_SLICE_X14Y109_CO6),
.O5(CLBLM_R_X11Y109_SLICE_X14Y109_BO5),
.O6(CLBLM_R_X11Y109_SLICE_X14Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h99559955f1f5f1f5)
  ) CLBLM_R_X11Y109_SLICE_X14Y109_ALUT (
.I0(CLBLM_L_X10Y106_SLICE_X12Y106_BO6),
.I1(RIOB33_X105Y101_IOB_X1Y102_I),
.I2(CLBLM_R_X11Y108_SLICE_X15Y108_AO6),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y109_SLICE_X14Y109_AO5),
.O6(CLBLM_R_X11Y109_SLICE_X14Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y109_SLICE_X15Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y109_SLICE_X15Y109_DO5),
.O6(CLBLM_R_X11Y109_SLICE_X15Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y109_SLICE_X15Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y109_SLICE_X15Y109_CO5),
.O6(CLBLM_R_X11Y109_SLICE_X15Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y109_SLICE_X15Y109_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y109_SLICE_X15Y109_BO5),
.O6(CLBLM_R_X11Y109_SLICE_X15Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h10223022ba001a00)
  ) CLBLM_R_X11Y109_SLICE_X15Y109_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y102_I),
.I1(RIOB33_X105Y101_IOB_X1Y101_I),
.I2(RIOB33_X105Y103_IOB_X1Y103_I),
.I3(RIOB33_X105Y113_IOB_X1Y113_I),
.I4(RIOB33_X105Y111_IOB_X1Y112_I),
.I5(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O5(CLBLM_R_X11Y109_SLICE_X15Y109_AO5),
.O6(CLBLM_R_X11Y109_SLICE_X15Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y110_SLICE_X14Y110_DO5),
.O6(CLBLM_R_X11Y110_SLICE_X14Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y110_SLICE_X14Y110_CO5),
.O6(CLBLM_R_X11Y110_SLICE_X14Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he12d78b469a53cf0)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_BLUT (
.I0(CLBLM_L_X10Y110_SLICE_X13Y110_AO5),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(CLBLM_R_X11Y109_SLICE_X14Y109_CO6),
.I3(RIOB33_X105Y101_IOB_X1Y102_I),
.I4(CLBLM_R_X11Y109_SLICE_X14Y109_AO6),
.I5(RIOB33_X105Y101_IOB_X1Y101_I),
.O5(CLBLM_R_X11Y110_SLICE_X14Y110_BO5),
.O6(CLBLM_R_X11Y110_SLICE_X14Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7777777755ff55ff)
  ) CLBLM_R_X11Y110_SLICE_X14Y110_ALUT (
.I0(RIOB33_X105Y101_IOB_X1Y101_I),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(1'b1),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y110_SLICE_X14Y110_AO5),
.O6(CLBLM_R_X11Y110_SLICE_X14Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y110_SLICE_X15Y110_DO5),
.O6(CLBLM_R_X11Y110_SLICE_X15Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y110_SLICE_X15Y110_CO5),
.O6(CLBLM_R_X11Y110_SLICE_X15Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y110_SLICE_X15Y110_BO5),
.O6(CLBLM_R_X11Y110_SLICE_X15Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y110_SLICE_X15Y110_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y110_SLICE_X15Y110_AO5),
.O6(CLBLM_R_X11Y110_SLICE_X15Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y101_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y101_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y102_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y102_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y103_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y103_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y104_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y104_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y105_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y105_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y106_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y106_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y107_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y107_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y108_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y108_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y109_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y109_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y110_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y110_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y111_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y111_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y112_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y112_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y113_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y113_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y114_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y114_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y115_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y115_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y116_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y116_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y117_IOB_X0Y117_IBUF (
.I(LIOB33_X0Y117_IOB_X0Y117_IPAD),
.O(LIOB33_X0Y117_IOB_X0Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y117_IOB_X0Y118_OBUF (
.I(CLBLL_L_X2Y113_SLICE_X0Y113_AO5),
.O(LIOB33_X0Y117_IOB_X0Y118_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUF (
.I(CLBLM_R_X3Y109_SLICE_X2Y109_BO5),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUF (
.I(CLBLL_L_X2Y112_SLICE_X0Y112_AO5),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUF (
.I(CLBLL_L_X2Y112_SLICE_X0Y112_BO5),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUF (
.I(CLBLM_R_X3Y109_SLICE_X2Y109_AO6),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUF (
.I(CLBLL_L_X2Y112_SLICE_X1Y112_BO6),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(CLBLM_R_X3Y113_SLICE_X2Y113_AO6),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y125_OBUF (
.I(CLBLM_R_X3Y112_SLICE_X3Y112_AO6),
.O(LIOB33_X0Y125_IOB_X0Y125_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y125_IOB_X0Y126_OBUF (
.I(CLBLM_R_X3Y113_SLICE_X3Y113_AO6),
.O(LIOB33_X0Y125_IOB_X0Y126_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y127_OBUF (
.I(CLBLM_R_X3Y111_SLICE_X3Y111_BO5),
.O(LIOB33_X0Y127_IOB_X0Y127_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y127_IOB_X0Y128_OBUF (
.I(CLBLM_R_X3Y110_SLICE_X3Y110_AO6),
.O(LIOB33_X0Y127_IOB_X0Y128_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y129_OBUF (
.I(CLBLM_R_X3Y110_SLICE_X2Y110_DO6),
.O(LIOB33_X0Y129_IOB_X0Y129_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y129_IOB_X0Y130_OBUF (
.I(CLBLL_L_X2Y113_SLICE_X0Y113_AO6),
.O(LIOB33_X0Y129_IOB_X0Y130_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y131_OBUF (
.I(CLBLM_R_X3Y109_SLICE_X3Y109_AO6),
.O(LIOB33_X0Y131_IOB_X0Y131_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y131_IOB_X0Y132_OBUF (
.I(CLBLM_R_X3Y107_SLICE_X2Y107_AO6),
.O(LIOB33_X0Y131_IOB_X0Y132_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y133_OBUF (
.I(CLBLL_L_X4Y109_SLICE_X5Y109_AO6),
.O(LIOB33_X0Y133_IOB_X0Y133_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y133_IOB_X0Y134_OBUF (
.I(1'b0),
.O(LIOB33_X0Y133_IOB_X0Y134_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y135_OBUF (
.I(CLBLM_R_X3Y107_SLICE_X3Y107_AO6),
.O(LIOB33_X0Y135_IOB_X0Y135_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y135_IOB_X0Y136_OBUF (
.I(CLBLM_R_X3Y108_SLICE_X3Y108_AO6),
.O(LIOB33_X0Y135_IOB_X0Y136_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y137_OBUF (
.I(CLBLL_L_X4Y107_SLICE_X4Y107_AO5),
.O(LIOB33_X0Y137_IOB_X0Y137_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y137_IOB_X0Y138_OBUF (
.I(CLBLL_L_X4Y107_SLICE_X4Y107_AO6),
.O(LIOB33_X0Y137_IOB_X0Y138_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y139_OBUF (
.I(CLBLL_L_X4Y106_SLICE_X4Y106_BO6),
.O(LIOB33_X0Y139_IOB_X0Y139_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y139_IOB_X0Y140_OBUF (
.I(CLBLL_L_X4Y106_SLICE_X4Y106_BO5),
.O(LIOB33_X0Y139_IOB_X0Y140_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y141_OBUF (
.I(CLBLM_R_X3Y104_SLICE_X3Y104_AO6),
.O(LIOB33_X0Y141_IOB_X0Y141_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y141_IOB_X0Y142_OBUF (
.I(CLBLM_R_X3Y104_SLICE_X3Y104_AO5),
.O(LIOB33_X0Y141_IOB_X0Y142_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y143_IOB_X0Y143_OBUF (
.I(CLBLM_R_X3Y104_SLICE_X2Y104_DO6),
.O(LIOB33_X0Y143_IOB_X0Y143_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y145_OBUF (
.I(CLBLM_R_X3Y103_SLICE_X2Y103_DO6),
.O(LIOB33_X0Y145_IOB_X0Y145_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y145_IOB_X0Y146_OBUF (
.I(CLBLM_R_X3Y103_SLICE_X2Y103_AO6),
.O(LIOB33_X0Y145_IOB_X0Y146_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y147_OBUF (
.I(CLBLL_L_X2Y106_SLICE_X0Y106_AO6),
.O(LIOB33_X0Y147_IOB_X0Y147_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y147_IOB_X0Y148_OBUF (
.I(CLBLL_L_X2Y106_SLICE_X0Y106_CO6),
.O(LIOB33_X0Y147_IOB_X0Y148_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y100_IOB_X0Y100_IBUF (
.I(LIOB33_SING_X0Y100_IOB_X0Y100_IPAD),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y149_IOB_X0Y149_OBUF (
.I(CLBLL_L_X2Y106_SLICE_X0Y106_AO5),
.O(LIOB33_SING_X0Y149_IOB_X0Y149_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y101_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y101_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y101_IOB_X1Y102_IBUF (
.I(RIOB33_X105Y101_IOB_X1Y102_IPAD),
.O(RIOB33_X105Y101_IOB_X1Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y103_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y103_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y103_IOB_X1Y104_IBUF (
.I(RIOB33_X105Y103_IOB_X1Y104_IPAD),
.O(RIOB33_X105Y103_IOB_X1Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y105_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y105_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y105_IOB_X1Y106_IBUF (
.I(RIOB33_X105Y105_IOB_X1Y106_IPAD),
.O(RIOB33_X105Y105_IOB_X1Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y107_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y107_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y107_IOB_X1Y108_IBUF (
.I(RIOB33_X105Y107_IOB_X1Y108_IPAD),
.O(RIOB33_X105Y107_IOB_X1Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y109_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y109_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y109_IOB_X1Y110_IBUF (
.I(RIOB33_X105Y109_IOB_X1Y110_IPAD),
.O(RIOB33_X105Y109_IOB_X1Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y111_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y111_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y111_IOB_X1Y112_IBUF (
.I(RIOB33_X105Y111_IOB_X1Y112_IPAD),
.O(RIOB33_X105Y111_IOB_X1Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_X105Y113_IOB_X1Y113_IBUF (
.I(RIOB33_X105Y113_IOB_X1Y113_IPAD),
.O(RIOB33_X105Y113_IOB_X1Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) RIOB33_SING_X105Y100_IOB_X1Y100_IBUF (
.I(RIOB33_SING_X105Y100_IOB_X1Y100_IPAD),
.O(RIOB33_SING_X105Y100_IOB_X1Y100_I)
  );
  assign CLBLL_L_X2Y103_SLICE_X0Y103_A = CLBLL_L_X2Y103_SLICE_X0Y103_AO6;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_B = CLBLL_L_X2Y103_SLICE_X0Y103_BO6;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_C = CLBLL_L_X2Y103_SLICE_X0Y103_CO6;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_D = CLBLL_L_X2Y103_SLICE_X0Y103_DO6;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_AMUX = CLBLL_L_X2Y103_SLICE_X0Y103_AO5;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_A = CLBLL_L_X2Y103_SLICE_X1Y103_AO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_B = CLBLL_L_X2Y103_SLICE_X1Y103_BO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_C = CLBLL_L_X2Y103_SLICE_X1Y103_CO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_D = CLBLL_L_X2Y103_SLICE_X1Y103_DO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_CMUX = CLBLL_L_X2Y103_SLICE_X1Y103_CO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A = CLBLL_L_X2Y104_SLICE_X0Y104_AO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B = CLBLL_L_X2Y104_SLICE_X0Y104_BO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C = CLBLL_L_X2Y104_SLICE_X0Y104_CO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D = CLBLL_L_X2Y104_SLICE_X0Y104_DO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A = CLBLL_L_X2Y104_SLICE_X1Y104_AO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B = CLBLL_L_X2Y104_SLICE_X1Y104_BO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C = CLBLL_L_X2Y104_SLICE_X1Y104_CO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D = CLBLL_L_X2Y104_SLICE_X1Y104_DO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A = CLBLL_L_X2Y105_SLICE_X0Y105_AO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B = CLBLL_L_X2Y105_SLICE_X0Y105_BO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C = CLBLL_L_X2Y105_SLICE_X0Y105_CO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D = CLBLL_L_X2Y105_SLICE_X0Y105_DO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A = CLBLL_L_X2Y105_SLICE_X1Y105_AO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B = CLBLL_L_X2Y105_SLICE_X1Y105_BO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C = CLBLL_L_X2Y105_SLICE_X1Y105_CO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D = CLBLL_L_X2Y105_SLICE_X1Y105_DO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A = CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B = CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C = CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D = CLBLL_L_X2Y106_SLICE_X0Y106_DO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_AMUX = CLBLL_L_X2Y106_SLICE_X0Y106_AO5;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A = CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B = CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C = CLBLL_L_X2Y106_SLICE_X1Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D = CLBLL_L_X2Y106_SLICE_X1Y106_DO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A = CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B = CLBLL_L_X2Y110_SLICE_X0Y110_BO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C = CLBLL_L_X2Y110_SLICE_X0Y110_CO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D = CLBLL_L_X2Y110_SLICE_X0Y110_DO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A = CLBLL_L_X2Y110_SLICE_X1Y110_AO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B = CLBLL_L_X2Y110_SLICE_X1Y110_BO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C = CLBLL_L_X2Y110_SLICE_X1Y110_CO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D = CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A = CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B = CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C = CLBLL_L_X2Y111_SLICE_X0Y111_CO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D = CLBLL_L_X2Y111_SLICE_X0Y111_DO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_AMUX = CLBLL_L_X2Y111_SLICE_X0Y111_AO5;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_CMUX = CLBLL_L_X2Y111_SLICE_X0Y111_CO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A = CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B = CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C = CLBLL_L_X2Y111_SLICE_X1Y111_CO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D = CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_AMUX = CLBLL_L_X2Y111_SLICE_X1Y111_AO5;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_BMUX = CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B = CLBLL_L_X2Y112_SLICE_X0Y112_BO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C = CLBLL_L_X2Y112_SLICE_X0Y112_CO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D = CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_AMUX = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_BMUX = CLBLL_L_X2Y112_SLICE_X0Y112_BO5;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_CMUX = CLBLL_L_X2Y112_SLICE_X0Y112_CO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A = CLBLL_L_X2Y112_SLICE_X1Y112_AO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B = CLBLL_L_X2Y112_SLICE_X1Y112_BO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C = CLBLL_L_X2Y112_SLICE_X1Y112_CO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D = CLBLL_L_X2Y112_SLICE_X1Y112_DO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_AMUX = CLBLL_L_X2Y112_SLICE_X1Y112_AO5;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A = CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B = CLBLL_L_X2Y113_SLICE_X0Y113_BO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C = CLBLL_L_X2Y113_SLICE_X0Y113_CO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D = CLBLL_L_X2Y113_SLICE_X0Y113_DO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_AMUX = CLBLL_L_X2Y113_SLICE_X0Y113_AO5;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A = CLBLL_L_X2Y113_SLICE_X1Y113_AO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B = CLBLL_L_X2Y113_SLICE_X1Y113_BO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C = CLBLL_L_X2Y113_SLICE_X1Y113_CO6;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D = CLBLL_L_X2Y113_SLICE_X1Y113_DO6;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_A = CLBLL_L_X4Y101_SLICE_X4Y101_AO6;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_B = CLBLL_L_X4Y101_SLICE_X4Y101_BO6;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_C = CLBLL_L_X4Y101_SLICE_X4Y101_CO6;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_D = CLBLL_L_X4Y101_SLICE_X4Y101_DO6;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_AMUX = CLBLL_L_X4Y101_SLICE_X4Y101_AO5;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_A = CLBLL_L_X4Y101_SLICE_X5Y101_AO6;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_B = CLBLL_L_X4Y101_SLICE_X5Y101_BO6;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_C = CLBLL_L_X4Y101_SLICE_X5Y101_CO6;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_D = CLBLL_L_X4Y101_SLICE_X5Y101_DO6;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_A = CLBLL_L_X4Y102_SLICE_X4Y102_AO6;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_B = CLBLL_L_X4Y102_SLICE_X4Y102_BO6;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_C = CLBLL_L_X4Y102_SLICE_X4Y102_CO6;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_D = CLBLL_L_X4Y102_SLICE_X4Y102_DO6;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_AMUX = CLBLL_L_X4Y102_SLICE_X4Y102_AO5;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_A = CLBLL_L_X4Y102_SLICE_X5Y102_AO6;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_B = CLBLL_L_X4Y102_SLICE_X5Y102_BO6;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_C = CLBLL_L_X4Y102_SLICE_X5Y102_CO6;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_D = CLBLL_L_X4Y102_SLICE_X5Y102_DO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A = CLBLL_L_X4Y103_SLICE_X4Y103_AO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B = CLBLL_L_X4Y103_SLICE_X4Y103_BO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C = CLBLL_L_X4Y103_SLICE_X4Y103_CO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D = CLBLL_L_X4Y103_SLICE_X4Y103_DO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_AMUX = CLBLL_L_X4Y103_SLICE_X4Y103_AO5;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_BMUX = CLBLL_L_X4Y103_SLICE_X4Y103_BO5;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A = CLBLL_L_X4Y103_SLICE_X5Y103_AO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B = CLBLL_L_X4Y103_SLICE_X5Y103_BO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C = CLBLL_L_X4Y103_SLICE_X5Y103_CO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D = CLBLL_L_X4Y103_SLICE_X5Y103_DO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_AMUX = CLBLL_L_X4Y103_SLICE_X5Y103_AO5;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_BMUX = CLBLL_L_X4Y103_SLICE_X5Y103_BO5;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A = CLBLL_L_X4Y104_SLICE_X4Y104_AO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B = CLBLL_L_X4Y104_SLICE_X4Y104_BO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C = CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D = CLBLL_L_X4Y104_SLICE_X4Y104_DO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_AMUX = CLBLL_L_X4Y104_SLICE_X4Y104_AO5;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_BMUX = CLBLL_L_X4Y104_SLICE_X4Y104_BO5;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_CMUX = CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_DMUX = CLBLL_L_X4Y104_SLICE_X4Y104_DO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A = CLBLL_L_X4Y104_SLICE_X5Y104_AO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B = CLBLL_L_X4Y104_SLICE_X5Y104_BO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C = CLBLL_L_X4Y104_SLICE_X5Y104_CO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D = CLBLL_L_X4Y104_SLICE_X5Y104_DO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_AMUX = CLBLL_L_X4Y104_SLICE_X5Y104_AO5;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A = CLBLL_L_X4Y105_SLICE_X4Y105_AO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B = CLBLL_L_X4Y105_SLICE_X4Y105_BO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C = CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D = CLBLL_L_X4Y105_SLICE_X4Y105_DO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A = CLBLL_L_X4Y105_SLICE_X5Y105_AO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C = CLBLL_L_X4Y105_SLICE_X5Y105_CO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D = CLBLL_L_X4Y105_SLICE_X5Y105_DO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_AMUX = CLBLL_L_X4Y105_SLICE_X5Y105_AO5;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_BMUX = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A = CLBLL_L_X4Y106_SLICE_X4Y106_AO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B = CLBLL_L_X4Y106_SLICE_X4Y106_BO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C = CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D = CLBLL_L_X4Y106_SLICE_X4Y106_DO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_AMUX = CLBLL_L_X4Y106_SLICE_X4Y106_AO5;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_BMUX = CLBLL_L_X4Y106_SLICE_X4Y106_BO5;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A = CLBLL_L_X4Y106_SLICE_X5Y106_AO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B = CLBLL_L_X4Y106_SLICE_X5Y106_BO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C = CLBLL_L_X4Y106_SLICE_X5Y106_CO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D = CLBLL_L_X4Y106_SLICE_X5Y106_DO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_AMUX = CLBLL_L_X4Y106_SLICE_X5Y106_AO5;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A = CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B = CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C = CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D = CLBLL_L_X4Y107_SLICE_X4Y107_DO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_AMUX = CLBLL_L_X4Y107_SLICE_X4Y107_AO5;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_BMUX = CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A = CLBLL_L_X4Y107_SLICE_X5Y107_AO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B = CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C = CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D = CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_AMUX = CLBLL_L_X4Y107_SLICE_X5Y107_AO5;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B = CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D = CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_AMUX = CLBLL_L_X4Y108_SLICE_X4Y108_AO5;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_CMUX = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A = CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B = CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C = CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D = CLBLL_L_X4Y108_SLICE_X5Y108_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A = CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B = CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_DMUX = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A = CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B = CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C = CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D = CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A = CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B = CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C = CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_AMUX = CLBLL_L_X4Y111_SLICE_X4Y111_AO5;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_BMUX = CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A = CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B = CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D = CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_AMUX = CLBLL_L_X4Y111_SLICE_X5Y111_AO5;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A = CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B = CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D = CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_AMUX = CLBLL_L_X4Y112_SLICE_X4Y112_AO5;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_BMUX = CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A = CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C = CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D = CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_AMUX = CLBLL_L_X4Y112_SLICE_X5Y112_AO5;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_BMUX = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A = CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C = CLBLL_L_X4Y113_SLICE_X4Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D = CLBLL_L_X4Y113_SLICE_X4Y113_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A = CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C = CLBLL_L_X4Y113_SLICE_X5Y113_CO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D = CLBLL_L_X4Y113_SLICE_X5Y113_DO6;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_A = CLBLM_L_X8Y101_SLICE_X10Y101_AO6;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_B = CLBLM_L_X8Y101_SLICE_X10Y101_BO6;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_C = CLBLM_L_X8Y101_SLICE_X10Y101_CO6;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_D = CLBLM_L_X8Y101_SLICE_X10Y101_DO6;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_A = CLBLM_L_X8Y101_SLICE_X11Y101_AO6;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_B = CLBLM_L_X8Y101_SLICE_X11Y101_BO6;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_C = CLBLM_L_X8Y101_SLICE_X11Y101_CO6;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_D = CLBLM_L_X8Y101_SLICE_X11Y101_DO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_A = CLBLM_L_X8Y102_SLICE_X10Y102_AO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_B = CLBLM_L_X8Y102_SLICE_X10Y102_BO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_C = CLBLM_L_X8Y102_SLICE_X10Y102_CO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_D = CLBLM_L_X8Y102_SLICE_X10Y102_DO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_AMUX = CLBLM_L_X8Y102_SLICE_X10Y102_AO5;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_A = CLBLM_L_X8Y102_SLICE_X11Y102_AO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_B = CLBLM_L_X8Y102_SLICE_X11Y102_BO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_C = CLBLM_L_X8Y102_SLICE_X11Y102_CO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_D = CLBLM_L_X8Y102_SLICE_X11Y102_DO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_AMUX = CLBLM_L_X8Y102_SLICE_X11Y102_AO5;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A = CLBLM_L_X8Y103_SLICE_X10Y103_AO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B = CLBLM_L_X8Y103_SLICE_X10Y103_BO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C = CLBLM_L_X8Y103_SLICE_X10Y103_CO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D = CLBLM_L_X8Y103_SLICE_X10Y103_DO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A = CLBLM_L_X8Y103_SLICE_X11Y103_AO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B = CLBLM_L_X8Y103_SLICE_X11Y103_BO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C = CLBLM_L_X8Y103_SLICE_X11Y103_CO6;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D = CLBLM_L_X8Y103_SLICE_X11Y103_DO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A = CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B = CLBLM_L_X8Y104_SLICE_X10Y104_BO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C = CLBLM_L_X8Y104_SLICE_X10Y104_CO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D = CLBLM_L_X8Y104_SLICE_X10Y104_DO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A = CLBLM_L_X8Y104_SLICE_X11Y104_AO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B = CLBLM_L_X8Y104_SLICE_X11Y104_BO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C = CLBLM_L_X8Y104_SLICE_X11Y104_CO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D = CLBLM_L_X8Y104_SLICE_X11Y104_DO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A = CLBLM_L_X8Y105_SLICE_X10Y105_AO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B = CLBLM_L_X8Y105_SLICE_X10Y105_BO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C = CLBLM_L_X8Y105_SLICE_X10Y105_CO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D = CLBLM_L_X8Y105_SLICE_X10Y105_DO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_AMUX = CLBLM_L_X8Y105_SLICE_X10Y105_AO5;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A = CLBLM_L_X8Y105_SLICE_X11Y105_AO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B = CLBLM_L_X8Y105_SLICE_X11Y105_BO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C = CLBLM_L_X8Y105_SLICE_X11Y105_CO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D = CLBLM_L_X8Y105_SLICE_X11Y105_DO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A = CLBLM_L_X8Y106_SLICE_X10Y106_AO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B = CLBLM_L_X8Y106_SLICE_X10Y106_BO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C = CLBLM_L_X8Y106_SLICE_X10Y106_CO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D = CLBLM_L_X8Y106_SLICE_X10Y106_DO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A = CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B = CLBLM_L_X8Y106_SLICE_X11Y106_BO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C = CLBLM_L_X8Y106_SLICE_X11Y106_CO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D = CLBLM_L_X8Y106_SLICE_X11Y106_DO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A = CLBLM_L_X8Y107_SLICE_X10Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B = CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C = CLBLM_L_X8Y107_SLICE_X10Y107_CO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D = CLBLM_L_X8Y107_SLICE_X10Y107_DO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_AMUX = CLBLM_L_X8Y107_SLICE_X10Y107_AO5;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A = CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B = CLBLM_L_X8Y107_SLICE_X11Y107_BO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C = CLBLM_L_X8Y107_SLICE_X11Y107_CO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D = CLBLM_L_X8Y107_SLICE_X11Y107_DO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_AMUX = CLBLM_L_X8Y107_SLICE_X11Y107_AO5;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A = CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B = CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C = CLBLM_L_X8Y108_SLICE_X10Y108_CO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D = CLBLM_L_X8Y108_SLICE_X10Y108_DO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A = CLBLM_L_X8Y108_SLICE_X11Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B = CLBLM_L_X8Y108_SLICE_X11Y108_BO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C = CLBLM_L_X8Y108_SLICE_X11Y108_CO6;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D = CLBLM_L_X8Y108_SLICE_X11Y108_DO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A = CLBLM_L_X8Y109_SLICE_X10Y109_AO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B = CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C = CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D = CLBLM_L_X8Y109_SLICE_X10Y109_DO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A = CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B = CLBLM_L_X8Y109_SLICE_X11Y109_BO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C = CLBLM_L_X8Y109_SLICE_X11Y109_CO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D = CLBLM_L_X8Y109_SLICE_X11Y109_DO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_AMUX = CLBLM_L_X8Y109_SLICE_X11Y109_AO5;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A = CLBLM_L_X8Y110_SLICE_X10Y110_AO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B = CLBLM_L_X8Y110_SLICE_X10Y110_BO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C = CLBLM_L_X8Y110_SLICE_X10Y110_CO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D = CLBLM_L_X8Y110_SLICE_X10Y110_DO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A = CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B = CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D = CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A = CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B = CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D = CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_AMUX = CLBLM_L_X8Y111_SLICE_X10Y111_AO5;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_BMUX = CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_CMUX = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A = CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B = CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D = CLBLM_L_X8Y111_SLICE_X11Y111_DO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A = CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B = CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C = CLBLM_L_X8Y112_SLICE_X10Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D = CLBLM_L_X8Y112_SLICE_X10Y112_DO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A = CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B = CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C = CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D = CLBLM_L_X8Y112_SLICE_X11Y112_DO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_AMUX = CLBLM_L_X8Y112_SLICE_X11Y112_AO5;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_CMUX = CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_A = CLBLM_L_X10Y101_SLICE_X12Y101_AO6;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_B = CLBLM_L_X10Y101_SLICE_X12Y101_BO6;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_C = CLBLM_L_X10Y101_SLICE_X12Y101_CO6;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_D = CLBLM_L_X10Y101_SLICE_X12Y101_DO6;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_A = CLBLM_L_X10Y101_SLICE_X13Y101_AO6;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_B = CLBLM_L_X10Y101_SLICE_X13Y101_BO6;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_C = CLBLM_L_X10Y101_SLICE_X13Y101_CO6;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_D = CLBLM_L_X10Y101_SLICE_X13Y101_DO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_A = CLBLM_L_X10Y102_SLICE_X12Y102_AO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_B = CLBLM_L_X10Y102_SLICE_X12Y102_BO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_C = CLBLM_L_X10Y102_SLICE_X12Y102_CO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_D = CLBLM_L_X10Y102_SLICE_X12Y102_DO6;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_A = CLBLM_L_X10Y102_SLICE_X13Y102_AO6;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_B = CLBLM_L_X10Y102_SLICE_X13Y102_BO6;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_C = CLBLM_L_X10Y102_SLICE_X13Y102_CO6;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_D = CLBLM_L_X10Y102_SLICE_X13Y102_DO6;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_AMUX = CLBLM_L_X10Y102_SLICE_X13Y102_AO5;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_BMUX = CLBLM_L_X10Y102_SLICE_X13Y102_BO5;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_CMUX = CLBLM_L_X10Y102_SLICE_X13Y102_CO5;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A = CLBLM_L_X10Y103_SLICE_X12Y103_AO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B = CLBLM_L_X10Y103_SLICE_X12Y103_BO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C = CLBLM_L_X10Y103_SLICE_X12Y103_CO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D = CLBLM_L_X10Y103_SLICE_X12Y103_DO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A = CLBLM_L_X10Y103_SLICE_X13Y103_AO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B = CLBLM_L_X10Y103_SLICE_X13Y103_BO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C = CLBLM_L_X10Y103_SLICE_X13Y103_CO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D = CLBLM_L_X10Y103_SLICE_X13Y103_DO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_AMUX = CLBLM_L_X10Y103_SLICE_X13Y103_AO5;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A = CLBLM_L_X10Y104_SLICE_X12Y104_AO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C = CLBLM_L_X10Y104_SLICE_X12Y104_CO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D = CLBLM_L_X10Y104_SLICE_X12Y104_DO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A = CLBLM_L_X10Y104_SLICE_X13Y104_AO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B = CLBLM_L_X10Y104_SLICE_X13Y104_BO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C = CLBLM_L_X10Y104_SLICE_X13Y104_CO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D = CLBLM_L_X10Y104_SLICE_X13Y104_DO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_BMUX = CLBLM_L_X10Y104_SLICE_X13Y104_BO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A = CLBLM_L_X10Y105_SLICE_X12Y105_AO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B = CLBLM_L_X10Y105_SLICE_X12Y105_BO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C = CLBLM_L_X10Y105_SLICE_X12Y105_CO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D = CLBLM_L_X10Y105_SLICE_X12Y105_DO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_AMUX = CLBLM_L_X10Y105_SLICE_X12Y105_AO5;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_BMUX = CLBLM_L_X10Y105_SLICE_X12Y105_BO5;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A = CLBLM_L_X10Y105_SLICE_X13Y105_AO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B = CLBLM_L_X10Y105_SLICE_X13Y105_BO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C = CLBLM_L_X10Y105_SLICE_X13Y105_CO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D = CLBLM_L_X10Y105_SLICE_X13Y105_DO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_AMUX = CLBLM_L_X10Y105_SLICE_X13Y105_AO5;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A = CLBLM_L_X10Y106_SLICE_X12Y106_AO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C = CLBLM_L_X10Y106_SLICE_X12Y106_CO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D = CLBLM_L_X10Y106_SLICE_X12Y106_DO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_AMUX = CLBLM_L_X10Y106_SLICE_X12Y106_AO5;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_CMUX = CLBLM_L_X10Y106_SLICE_X12Y106_CO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_DMUX = CLBLM_L_X10Y106_SLICE_X12Y106_DO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A = CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B = CLBLM_L_X10Y106_SLICE_X13Y106_BO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C = CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D = CLBLM_L_X10Y106_SLICE_X13Y106_DO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A = CLBLM_L_X10Y107_SLICE_X12Y107_AO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B = CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C = CLBLM_L_X10Y107_SLICE_X12Y107_CO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D = CLBLM_L_X10Y107_SLICE_X12Y107_DO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_AMUX = CLBLM_L_X10Y107_SLICE_X12Y107_AO5;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A = CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B = CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C = CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D = CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_AMUX = CLBLM_L_X10Y107_SLICE_X13Y107_AO5;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A = CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B = CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C = CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D = CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A = CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B = CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C = CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D = CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A = CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C = CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_AMUX = CLBLM_L_X10Y109_SLICE_X12Y109_AO5;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A = CLBLM_L_X10Y109_SLICE_X13Y109_AO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B = CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D = CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_AMUX = CLBLM_L_X10Y109_SLICE_X13Y109_AO5;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_BMUX = CLBLM_L_X10Y109_SLICE_X13Y109_BO5;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A = CLBLM_L_X10Y110_SLICE_X12Y110_AO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B = CLBLM_L_X10Y110_SLICE_X12Y110_BO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C = CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D = CLBLM_L_X10Y110_SLICE_X12Y110_DO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_DMUX = CLBLM_L_X10Y110_SLICE_X12Y110_DO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A = CLBLM_L_X10Y110_SLICE_X13Y110_AO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B = CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C = CLBLM_L_X10Y110_SLICE_X13Y110_CO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D = CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_AMUX = CLBLM_L_X10Y110_SLICE_X13Y110_AO5;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_BMUX = CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A = CLBLM_L_X10Y111_SLICE_X12Y111_AO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B = CLBLM_L_X10Y111_SLICE_X12Y111_BO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C = CLBLM_L_X10Y111_SLICE_X12Y111_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D = CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_AMUX = CLBLM_L_X10Y111_SLICE_X12Y111_AO5;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A = CLBLM_L_X10Y111_SLICE_X13Y111_AO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B = CLBLM_L_X10Y111_SLICE_X13Y111_BO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C = CLBLM_L_X10Y111_SLICE_X13Y111_CO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D = CLBLM_L_X10Y111_SLICE_X13Y111_DO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_A = CLBLM_L_X12Y104_SLICE_X16Y104_AO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_B = CLBLM_L_X12Y104_SLICE_X16Y104_BO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_C = CLBLM_L_X12Y104_SLICE_X16Y104_CO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_D = CLBLM_L_X12Y104_SLICE_X16Y104_DO6;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_A = CLBLM_L_X12Y104_SLICE_X17Y104_AO6;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_B = CLBLM_L_X12Y104_SLICE_X17Y104_BO6;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_C = CLBLM_L_X12Y104_SLICE_X17Y104_CO6;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_D = CLBLM_L_X12Y104_SLICE_X17Y104_DO6;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_A = CLBLM_R_X3Y102_SLICE_X2Y102_AO6;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_B = CLBLM_R_X3Y102_SLICE_X2Y102_BO6;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_C = CLBLM_R_X3Y102_SLICE_X2Y102_CO6;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_D = CLBLM_R_X3Y102_SLICE_X2Y102_DO6;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_AMUX = CLBLM_R_X3Y102_SLICE_X2Y102_AO6;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_BMUX = CLBLM_R_X3Y102_SLICE_X2Y102_BO6;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_A = CLBLM_R_X3Y102_SLICE_X3Y102_AO6;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_B = CLBLM_R_X3Y102_SLICE_X3Y102_BO6;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_C = CLBLM_R_X3Y102_SLICE_X3Y102_CO6;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_D = CLBLM_R_X3Y102_SLICE_X3Y102_DO6;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_AMUX = CLBLM_R_X3Y102_SLICE_X3Y102_AO5;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A = CLBLM_R_X3Y103_SLICE_X2Y103_AO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B = CLBLM_R_X3Y103_SLICE_X2Y103_BO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C = CLBLM_R_X3Y103_SLICE_X2Y103_CO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D = CLBLM_R_X3Y103_SLICE_X2Y103_DO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A = CLBLM_R_X3Y103_SLICE_X3Y103_AO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B = CLBLM_R_X3Y103_SLICE_X3Y103_BO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C = CLBLM_R_X3Y103_SLICE_X3Y103_CO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D = CLBLM_R_X3Y103_SLICE_X3Y103_DO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_AMUX = CLBLM_R_X3Y103_SLICE_X3Y103_AO5;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_CMUX = CLBLM_R_X3Y103_SLICE_X3Y103_CO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A = CLBLM_R_X3Y104_SLICE_X2Y104_AO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B = CLBLM_R_X3Y104_SLICE_X2Y104_BO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C = CLBLM_R_X3Y104_SLICE_X2Y104_CO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D = CLBLM_R_X3Y104_SLICE_X2Y104_DO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_AMUX = CLBLM_R_X3Y104_SLICE_X2Y104_AO5;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A = CLBLM_R_X3Y104_SLICE_X3Y104_AO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B = CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C = CLBLM_R_X3Y104_SLICE_X3Y104_CO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D = CLBLM_R_X3Y104_SLICE_X3Y104_DO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_AMUX = CLBLM_R_X3Y104_SLICE_X3Y104_AO5;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_BMUX = CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A = CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B = CLBLM_R_X3Y105_SLICE_X2Y105_BO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C = CLBLM_R_X3Y105_SLICE_X2Y105_CO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D = CLBLM_R_X3Y105_SLICE_X2Y105_DO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A = CLBLM_R_X3Y105_SLICE_X3Y105_AO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B = CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C = CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D = CLBLM_R_X3Y105_SLICE_X3Y105_DO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_AMUX = CLBLM_R_X3Y105_SLICE_X3Y105_AO5;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_BMUX = CLBLM_R_X3Y105_SLICE_X3Y105_BO5;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_CMUX = CLBLM_R_X3Y105_SLICE_X3Y105_CO5;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A = CLBLM_R_X3Y106_SLICE_X2Y106_AO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B = CLBLM_R_X3Y106_SLICE_X2Y106_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C = CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D = CLBLM_R_X3Y106_SLICE_X2Y106_DO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A = CLBLM_R_X3Y106_SLICE_X3Y106_AO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B = CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C = CLBLM_R_X3Y106_SLICE_X3Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D = CLBLM_R_X3Y106_SLICE_X3Y106_DO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_AMUX = CLBLM_R_X3Y106_SLICE_X3Y106_AO5;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A = CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B = CLBLM_R_X3Y107_SLICE_X2Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C = CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D = CLBLM_R_X3Y107_SLICE_X2Y107_DO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_AMUX = CLBLM_R_X3Y107_SLICE_X2Y107_AO5;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_CMUX = CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A = CLBLM_R_X3Y107_SLICE_X3Y107_AO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B = CLBLM_R_X3Y107_SLICE_X3Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C = CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D = CLBLM_R_X3Y107_SLICE_X3Y107_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_DMUX = CLBLM_R_X3Y107_SLICE_X3Y107_DO5;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A = CLBLM_R_X3Y108_SLICE_X2Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B = CLBLM_R_X3Y108_SLICE_X2Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C = CLBLM_R_X3Y108_SLICE_X2Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D = CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A = CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B = CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C = CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A = CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B = CLBLM_R_X3Y109_SLICE_X2Y109_BO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D = CLBLM_R_X3Y109_SLICE_X2Y109_DO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_AMUX = CLBLM_R_X3Y109_SLICE_X2Y109_AO5;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_BMUX = CLBLM_R_X3Y109_SLICE_X2Y109_BO5;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A = CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B = CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C = CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D = CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_AMUX = CLBLM_R_X3Y109_SLICE_X3Y109_AO5;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A = CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C = CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_AMUX = CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B = CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C = CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_AMUX = CLBLM_R_X3Y110_SLICE_X3Y110_AO5;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A = CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B = CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D = CLBLM_R_X3Y111_SLICE_X2Y111_DO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_AMUX = CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A = CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B = CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C = CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_AMUX = CLBLM_R_X3Y111_SLICE_X3Y111_AO5;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_BMUX = CLBLM_R_X3Y111_SLICE_X3Y111_BO5;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_CMUX = CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A = CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B = CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C = CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D = CLBLM_R_X3Y112_SLICE_X2Y112_DO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A = CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C = CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D = CLBLM_R_X3Y112_SLICE_X3Y112_DO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_AMUX = CLBLM_R_X3Y112_SLICE_X3Y112_AO5;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B = CLBLM_R_X3Y113_SLICE_X2Y113_BO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C = CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D = CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_AMUX = CLBLM_R_X3Y113_SLICE_X2Y113_AO5;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_BMUX = CLBLM_R_X3Y113_SLICE_X2Y113_BO5;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_CMUX = CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A = CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B = CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C = CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D = CLBLM_R_X3Y113_SLICE_X3Y113_DO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_BMUX = CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_A = CLBLM_R_X5Y100_SLICE_X6Y100_AO6;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_B = CLBLM_R_X5Y100_SLICE_X6Y100_BO6;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_C = CLBLM_R_X5Y100_SLICE_X6Y100_CO6;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_D = CLBLM_R_X5Y100_SLICE_X6Y100_DO6;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_A = CLBLM_R_X5Y100_SLICE_X7Y100_AO6;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_B = CLBLM_R_X5Y100_SLICE_X7Y100_BO6;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_C = CLBLM_R_X5Y100_SLICE_X7Y100_CO6;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_D = CLBLM_R_X5Y100_SLICE_X7Y100_DO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_A = CLBLM_R_X5Y101_SLICE_X6Y101_AO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_B = CLBLM_R_X5Y101_SLICE_X6Y101_BO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_C = CLBLM_R_X5Y101_SLICE_X6Y101_CO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_D = CLBLM_R_X5Y101_SLICE_X6Y101_DO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_AMUX = CLBLM_R_X5Y101_SLICE_X6Y101_AO5;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_A = CLBLM_R_X5Y101_SLICE_X7Y101_AO6;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_B = CLBLM_R_X5Y101_SLICE_X7Y101_BO6;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_C = CLBLM_R_X5Y101_SLICE_X7Y101_CO6;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_D = CLBLM_R_X5Y101_SLICE_X7Y101_DO6;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_AMUX = CLBLM_R_X5Y101_SLICE_X7Y101_AO5;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_A = CLBLM_R_X5Y102_SLICE_X6Y102_AO6;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_B = CLBLM_R_X5Y102_SLICE_X6Y102_BO6;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_C = CLBLM_R_X5Y102_SLICE_X6Y102_CO6;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_D = CLBLM_R_X5Y102_SLICE_X6Y102_DO6;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_CMUX = CLBLM_R_X5Y102_SLICE_X6Y102_CO6;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_A = CLBLM_R_X5Y102_SLICE_X7Y102_AO6;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_B = CLBLM_R_X5Y102_SLICE_X7Y102_BO6;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_C = CLBLM_R_X5Y102_SLICE_X7Y102_CO6;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_D = CLBLM_R_X5Y102_SLICE_X7Y102_DO6;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_AMUX = CLBLM_R_X5Y102_SLICE_X7Y102_AO5;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_BMUX = CLBLM_R_X5Y102_SLICE_X7Y102_BO5;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_A = CLBLM_R_X5Y103_SLICE_X6Y103_AO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_B = CLBLM_R_X5Y103_SLICE_X6Y103_BO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_C = CLBLM_R_X5Y103_SLICE_X6Y103_CO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_D = CLBLM_R_X5Y103_SLICE_X6Y103_DO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_AMUX = CLBLM_R_X5Y103_SLICE_X6Y103_AO5;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_A = CLBLM_R_X5Y103_SLICE_X7Y103_AO6;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_B = CLBLM_R_X5Y103_SLICE_X7Y103_BO6;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_C = CLBLM_R_X5Y103_SLICE_X7Y103_CO6;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_D = CLBLM_R_X5Y103_SLICE_X7Y103_DO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A = CLBLM_R_X5Y104_SLICE_X6Y104_AO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B = CLBLM_R_X5Y104_SLICE_X6Y104_BO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C = CLBLM_R_X5Y104_SLICE_X6Y104_CO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D = CLBLM_R_X5Y104_SLICE_X6Y104_DO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_AMUX = CLBLM_R_X5Y104_SLICE_X6Y104_AO5;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A = CLBLM_R_X5Y104_SLICE_X7Y104_AO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B = CLBLM_R_X5Y104_SLICE_X7Y104_BO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C = CLBLM_R_X5Y104_SLICE_X7Y104_CO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D = CLBLM_R_X5Y104_SLICE_X7Y104_DO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_AMUX = CLBLM_R_X5Y104_SLICE_X7Y104_AO5;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A = CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B = CLBLM_R_X5Y105_SLICE_X6Y105_BO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C = CLBLM_R_X5Y105_SLICE_X6Y105_CO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D = CLBLM_R_X5Y105_SLICE_X6Y105_DO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_AMUX = CLBLM_R_X5Y105_SLICE_X6Y105_AO5;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A = CLBLM_R_X5Y105_SLICE_X7Y105_AO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B = CLBLM_R_X5Y105_SLICE_X7Y105_BO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C = CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D = CLBLM_R_X5Y105_SLICE_X7Y105_DO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_AMUX = CLBLM_R_X5Y105_SLICE_X7Y105_AO5;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_BMUX = CLBLM_R_X5Y105_SLICE_X7Y105_BO5;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A = CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B = CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C = CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D = CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_AMUX = CLBLM_R_X5Y106_SLICE_X6Y106_AO5;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A = CLBLM_R_X5Y106_SLICE_X7Y106_AO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B = CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C = CLBLM_R_X5Y106_SLICE_X7Y106_CO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D = CLBLM_R_X5Y106_SLICE_X7Y106_DO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_AMUX = CLBLM_R_X5Y106_SLICE_X7Y106_AO5;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_BMUX = CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A = CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C = CLBLM_R_X5Y107_SLICE_X6Y107_CO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D = CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_DMUX = CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A = CLBLM_R_X5Y107_SLICE_X7Y107_AO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C = CLBLM_R_X5Y107_SLICE_X7Y107_CO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D = CLBLM_R_X5Y107_SLICE_X7Y107_DO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_AMUX = CLBLM_R_X5Y107_SLICE_X7Y107_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A = CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B = CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C = CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D = CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A = CLBLM_R_X5Y108_SLICE_X7Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B = CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C = CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D = CLBLM_R_X5Y108_SLICE_X7Y108_DO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_CMUX = CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A = CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B = CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C = CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D = CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_AMUX = CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A = CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B = CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C = CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D = CLBLM_R_X5Y109_SLICE_X7Y109_DO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_AMUX = CLBLM_R_X5Y109_SLICE_X7Y109_AO5;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B = CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D = CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A = CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B = CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C = CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D = CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_AMUX = CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B = CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C = CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_AMUX = CLBLM_R_X5Y111_SLICE_X6Y111_AO5;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A = CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B = CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C = CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_AMUX = CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_BMUX = CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A = CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B = CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C = CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D = CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_AMUX = CLBLM_R_X5Y112_SLICE_X6Y112_AO5;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A = CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B = CLBLM_R_X5Y112_SLICE_X7Y112_BO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C = CLBLM_R_X5Y112_SLICE_X7Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D = CLBLM_R_X5Y112_SLICE_X7Y112_DO6;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_A = CLBLM_R_X7Y100_SLICE_X8Y100_AO6;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_B = CLBLM_R_X7Y100_SLICE_X8Y100_BO6;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_C = CLBLM_R_X7Y100_SLICE_X8Y100_CO6;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_D = CLBLM_R_X7Y100_SLICE_X8Y100_DO6;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_AMUX = CLBLM_R_X7Y100_SLICE_X8Y100_AO5;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_BMUX = CLBLM_R_X7Y100_SLICE_X8Y100_BO5;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_A = CLBLM_R_X7Y100_SLICE_X9Y100_AO6;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_B = CLBLM_R_X7Y100_SLICE_X9Y100_BO6;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_C = CLBLM_R_X7Y100_SLICE_X9Y100_CO6;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_D = CLBLM_R_X7Y100_SLICE_X9Y100_DO6;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_A = CLBLM_R_X7Y101_SLICE_X8Y101_AO6;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_B = CLBLM_R_X7Y101_SLICE_X8Y101_BO6;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_C = CLBLM_R_X7Y101_SLICE_X8Y101_CO6;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_D = CLBLM_R_X7Y101_SLICE_X8Y101_DO6;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_AMUX = CLBLM_R_X7Y101_SLICE_X8Y101_AO5;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_BMUX = CLBLM_R_X7Y101_SLICE_X8Y101_BO5;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_CMUX = CLBLM_R_X7Y101_SLICE_X8Y101_CO5;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_A = CLBLM_R_X7Y101_SLICE_X9Y101_AO6;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_B = CLBLM_R_X7Y101_SLICE_X9Y101_BO6;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_C = CLBLM_R_X7Y101_SLICE_X9Y101_CO6;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_D = CLBLM_R_X7Y101_SLICE_X9Y101_DO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_A = CLBLM_R_X7Y102_SLICE_X8Y102_AO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_B = CLBLM_R_X7Y102_SLICE_X8Y102_BO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_C = CLBLM_R_X7Y102_SLICE_X8Y102_CO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_D = CLBLM_R_X7Y102_SLICE_X8Y102_DO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_AMUX = CLBLM_R_X7Y102_SLICE_X8Y102_AO5;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_A = CLBLM_R_X7Y102_SLICE_X9Y102_AO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_B = CLBLM_R_X7Y102_SLICE_X9Y102_BO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_C = CLBLM_R_X7Y102_SLICE_X9Y102_CO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_D = CLBLM_R_X7Y102_SLICE_X9Y102_DO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A = CLBLM_R_X7Y103_SLICE_X8Y103_AO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B = CLBLM_R_X7Y103_SLICE_X8Y103_BO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C = CLBLM_R_X7Y103_SLICE_X8Y103_CO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D = CLBLM_R_X7Y103_SLICE_X8Y103_DO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_AMUX = CLBLM_R_X7Y103_SLICE_X8Y103_AO5;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A = CLBLM_R_X7Y103_SLICE_X9Y103_AO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B = CLBLM_R_X7Y103_SLICE_X9Y103_BO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C = CLBLM_R_X7Y103_SLICE_X9Y103_CO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D = CLBLM_R_X7Y103_SLICE_X9Y103_DO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_AMUX = CLBLM_R_X7Y103_SLICE_X9Y103_AO5;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_CMUX = CLBLM_R_X7Y103_SLICE_X9Y103_CO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A = CLBLM_R_X7Y104_SLICE_X8Y104_AO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B = CLBLM_R_X7Y104_SLICE_X8Y104_BO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C = CLBLM_R_X7Y104_SLICE_X8Y104_CO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D = CLBLM_R_X7Y104_SLICE_X8Y104_DO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_AMUX = CLBLM_R_X7Y104_SLICE_X8Y104_AO5;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_BMUX = CLBLM_R_X7Y104_SLICE_X8Y104_BO5;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_DMUX = CLBLM_R_X7Y104_SLICE_X8Y104_DO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A = CLBLM_R_X7Y104_SLICE_X9Y104_AO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B = CLBLM_R_X7Y104_SLICE_X9Y104_BO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C = CLBLM_R_X7Y104_SLICE_X9Y104_CO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D = CLBLM_R_X7Y104_SLICE_X9Y104_DO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_AMUX = CLBLM_R_X7Y104_SLICE_X9Y104_AO5;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A = CLBLM_R_X7Y105_SLICE_X8Y105_AO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B = CLBLM_R_X7Y105_SLICE_X8Y105_BO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C = CLBLM_R_X7Y105_SLICE_X8Y105_CO6;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D = CLBLM_R_X7Y105_SLICE_X8Y105_DO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A = CLBLM_R_X7Y105_SLICE_X9Y105_AO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B = CLBLM_R_X7Y105_SLICE_X9Y105_BO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C = CLBLM_R_X7Y105_SLICE_X9Y105_CO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D = CLBLM_R_X7Y105_SLICE_X9Y105_DO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A = CLBLM_R_X7Y106_SLICE_X8Y106_AO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B = CLBLM_R_X7Y106_SLICE_X8Y106_BO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C = CLBLM_R_X7Y106_SLICE_X8Y106_CO6;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D = CLBLM_R_X7Y106_SLICE_X8Y106_DO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A = CLBLM_R_X7Y106_SLICE_X9Y106_AO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B = CLBLM_R_X7Y106_SLICE_X9Y106_BO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C = CLBLM_R_X7Y106_SLICE_X9Y106_CO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D = CLBLM_R_X7Y106_SLICE_X9Y106_DO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_AMUX = CLBLM_R_X7Y106_SLICE_X9Y106_AO5;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A = CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B = CLBLM_R_X7Y107_SLICE_X8Y107_BO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C = CLBLM_R_X7Y107_SLICE_X8Y107_CO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D = CLBLM_R_X7Y107_SLICE_X8Y107_DO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A = CLBLM_R_X7Y107_SLICE_X9Y107_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B = CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C = CLBLM_R_X7Y107_SLICE_X9Y107_CO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D = CLBLM_R_X7Y107_SLICE_X9Y107_DO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_AMUX = CLBLM_R_X7Y107_SLICE_X9Y107_AO5;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_BMUX = CLBLM_R_X7Y107_SLICE_X9Y107_BO5;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_CMUX = CLBLM_R_X7Y107_SLICE_X9Y107_CO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B = CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C = CLBLM_R_X7Y108_SLICE_X8Y108_CO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D = CLBLM_R_X7Y108_SLICE_X8Y108_DO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A = CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B = CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C = CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D = CLBLM_R_X7Y108_SLICE_X9Y108_DO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_AMUX = CLBLM_R_X7Y108_SLICE_X9Y108_AO5;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_BMUX = CLBLM_R_X7Y108_SLICE_X9Y108_BO5;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A = CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B = CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C = CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D = CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A = CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B = CLBLM_R_X7Y109_SLICE_X9Y109_BO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C = CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D = CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_AMUX = CLBLM_R_X7Y109_SLICE_X9Y109_AO5;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A = CLBLM_R_X7Y110_SLICE_X8Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B = CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D = CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_AMUX = CLBLM_R_X7Y110_SLICE_X8Y110_AO5;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A = CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B = CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C = CLBLM_R_X7Y110_SLICE_X9Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D = CLBLM_R_X7Y110_SLICE_X9Y110_DO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_AMUX = CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A = CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C = CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_AMUX = CLBLM_R_X7Y111_SLICE_X8Y111_AO5;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B = CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C = CLBLM_R_X7Y111_SLICE_X9Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D = CLBLM_R_X7Y111_SLICE_X9Y111_DO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B = CLBLM_R_X7Y112_SLICE_X8Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C = CLBLM_R_X7Y112_SLICE_X8Y112_CO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D = CLBLM_R_X7Y112_SLICE_X8Y112_DO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A = CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D = CLBLM_R_X7Y112_SLICE_X9Y112_DO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_AMUX = CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_A = CLBLM_R_X11Y103_SLICE_X14Y103_AO6;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_B = CLBLM_R_X11Y103_SLICE_X14Y103_BO6;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_C = CLBLM_R_X11Y103_SLICE_X14Y103_CO6;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_D = CLBLM_R_X11Y103_SLICE_X14Y103_DO6;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_AMUX = CLBLM_R_X11Y103_SLICE_X14Y103_AO6;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_A = CLBLM_R_X11Y103_SLICE_X15Y103_AO6;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_B = CLBLM_R_X11Y103_SLICE_X15Y103_BO6;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_C = CLBLM_R_X11Y103_SLICE_X15Y103_CO6;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_D = CLBLM_R_X11Y103_SLICE_X15Y103_DO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_A = CLBLM_R_X11Y104_SLICE_X14Y104_AO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_B = CLBLM_R_X11Y104_SLICE_X14Y104_BO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_C = CLBLM_R_X11Y104_SLICE_X14Y104_CO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_D = CLBLM_R_X11Y104_SLICE_X14Y104_DO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_AMUX = CLBLM_R_X11Y104_SLICE_X14Y104_AO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_A = CLBLM_R_X11Y104_SLICE_X15Y104_AO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_B = CLBLM_R_X11Y104_SLICE_X15Y104_BO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_C = CLBLM_R_X11Y104_SLICE_X15Y104_CO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_D = CLBLM_R_X11Y104_SLICE_X15Y104_DO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_AMUX = CLBLM_R_X11Y104_SLICE_X15Y104_AO5;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_BMUX = CLBLM_R_X11Y104_SLICE_X15Y104_BO5;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A = CLBLM_R_X11Y105_SLICE_X14Y105_AO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B = CLBLM_R_X11Y105_SLICE_X14Y105_BO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C = CLBLM_R_X11Y105_SLICE_X14Y105_CO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D = CLBLM_R_X11Y105_SLICE_X14Y105_DO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_AMUX = CLBLM_R_X11Y105_SLICE_X14Y105_AO5;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A = CLBLM_R_X11Y105_SLICE_X15Y105_AO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B = CLBLM_R_X11Y105_SLICE_X15Y105_BO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C = CLBLM_R_X11Y105_SLICE_X15Y105_CO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D = CLBLM_R_X11Y105_SLICE_X15Y105_DO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_CMUX = CLBLM_R_X11Y105_SLICE_X15Y105_CO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A = CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B = CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C = CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D = CLBLM_R_X11Y106_SLICE_X14Y106_DO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A = CLBLM_R_X11Y106_SLICE_X15Y106_AO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B = CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C = CLBLM_R_X11Y106_SLICE_X15Y106_CO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D = CLBLM_R_X11Y106_SLICE_X15Y106_DO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_AMUX = CLBLM_R_X11Y106_SLICE_X15Y106_AO5;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_BMUX = CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A = CLBLM_R_X11Y107_SLICE_X14Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B = CLBLM_R_X11Y107_SLICE_X14Y107_BO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C = CLBLM_R_X11Y107_SLICE_X14Y107_CO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D = CLBLM_R_X11Y107_SLICE_X14Y107_DO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_AMUX = CLBLM_R_X11Y107_SLICE_X14Y107_AO5;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A = CLBLM_R_X11Y107_SLICE_X15Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B = CLBLM_R_X11Y107_SLICE_X15Y107_BO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C = CLBLM_R_X11Y107_SLICE_X15Y107_CO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D = CLBLM_R_X11Y107_SLICE_X15Y107_DO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_AMUX = CLBLM_R_X11Y107_SLICE_X15Y107_AO5;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_CMUX = CLBLM_R_X11Y107_SLICE_X15Y107_CO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A = CLBLM_R_X11Y108_SLICE_X14Y108_AO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B = CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C = CLBLM_R_X11Y108_SLICE_X14Y108_CO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D = CLBLM_R_X11Y108_SLICE_X14Y108_DO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A = CLBLM_R_X11Y108_SLICE_X15Y108_AO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B = CLBLM_R_X11Y108_SLICE_X15Y108_BO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C = CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D = CLBLM_R_X11Y108_SLICE_X15Y108_DO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_AMUX = CLBLM_R_X11Y108_SLICE_X15Y108_AO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_CMUX = CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A = CLBLM_R_X11Y109_SLICE_X14Y109_AO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B = CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C = CLBLM_R_X11Y109_SLICE_X14Y109_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D = CLBLM_R_X11Y109_SLICE_X14Y109_DO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_AMUX = CLBLM_R_X11Y109_SLICE_X14Y109_AO5;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A = CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B = CLBLM_R_X11Y109_SLICE_X15Y109_BO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C = CLBLM_R_X11Y109_SLICE_X15Y109_CO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D = CLBLM_R_X11Y109_SLICE_X15Y109_DO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A = CLBLM_R_X11Y110_SLICE_X14Y110_AO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B = CLBLM_R_X11Y110_SLICE_X14Y110_BO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C = CLBLM_R_X11Y110_SLICE_X14Y110_CO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D = CLBLM_R_X11Y110_SLICE_X14Y110_DO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_AMUX = CLBLM_R_X11Y110_SLICE_X14Y110_AO5;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A = CLBLM_R_X11Y110_SLICE_X15Y110_AO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B = CLBLM_R_X11Y110_SLICE_X15Y110_BO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C = CLBLM_R_X11Y110_SLICE_X15Y110_CO6;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D = CLBLM_R_X11Y110_SLICE_X15Y110_DO6;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_O = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_O = LIOB33_X0Y101_IOB_X0Y101_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_O = LIOB33_X0Y103_IOB_X0Y104_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_O = LIOB33_X0Y103_IOB_X0Y103_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_O = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_O = LIOB33_X0Y105_IOB_X0Y105_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_O = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_O = LIOB33_X0Y109_IOB_X0Y109_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_O = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_O = LIOB33_X0Y111_IOB_X0Y111_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_O = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_O = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_O = LIOB33_X0Y117_IOB_X0Y117_I;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_OQ = CLBLL_L_X2Y113_SLICE_X0Y113_AO5;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = CLBLL_L_X2Y112_SLICE_X0Y112_BO5;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = CLBLL_L_X2Y112_SLICE_X1Y112_BO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_OQ = CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_TQ = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_OQ = CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_OQ = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_TQ = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_OQ = CLBLM_R_X3Y111_SLICE_X3Y111_BO5;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_OQ = CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_TQ = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_OQ = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_OQ = 1'b0;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_TQ = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_OQ = CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_OQ = CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_TQ = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_OQ = CLBLM_R_X3Y107_SLICE_X3Y107_AO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_OQ = CLBLL_L_X4Y106_SLICE_X4Y106_BO5;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_TQ = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_OQ = CLBLL_L_X4Y106_SLICE_X4Y106_BO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_OQ = CLBLM_R_X3Y104_SLICE_X3Y104_AO5;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_TQ = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_OQ = CLBLM_R_X3Y104_SLICE_X3Y104_AO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_OQ = CLBLM_R_X3Y103_SLICE_X2Y103_AO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_TQ = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_OQ = CLBLM_R_X3Y103_SLICE_X2Y103_DO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_OQ = CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_TQ = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_OQ = CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_TQ = 1'b1;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_O = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_OQ = CLBLL_L_X2Y106_SLICE_X0Y106_AO5;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O = LIOB33_X0Y107_IOB_X0Y107_I;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = CLBLM_R_X3Y109_SLICE_X2Y109_BO5;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_OQ = CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_OQ = CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_OQ = CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_OQ = CLBLM_R_X3Y104_SLICE_X2Y104_DO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O = LIOB33_X0Y113_IOB_X0Y113_I;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_OQ = CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_OQ = CLBLL_L_X4Y107_SLICE_X4Y107_AO5;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_TQ = 1'b1;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_O = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_O = RIOB33_X105Y101_IOB_X1Y101_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_O = RIOB33_X105Y103_IOB_X1Y104_I;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_O = RIOB33_X105Y103_IOB_X1Y103_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_O = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_O = RIOB33_X105Y105_IOB_X1Y105_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_O = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_O = RIOB33_X105Y109_IOB_X1Y109_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_O = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_O = RIOB33_X105Y111_IOB_X1Y111_I;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_O = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_O = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_O = RIOB33_X105Y107_IOB_X1Y107_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_O = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D1 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D2 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D3 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D4 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D5 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_D6 = 1'b1;
  assign LIOB33_X0Y147_IOB_X0Y147_O = CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  assign LIOB33_X0Y147_IOB_X0Y148_O = CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B5 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B6 = 1'b1;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_A1 = CLBLM_R_X5Y102_SLICE_X7Y102_DO6;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_A3 = CLBLL_L_X4Y102_SLICE_X5Y102_DO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A1 = CLBLM_L_X10Y105_SLICE_X12Y105_BO5;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A2 = CLBLM_L_X10Y105_SLICE_X13Y105_AO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A3 = CLBLM_L_X10Y102_SLICE_X13Y102_DO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A4 = CLBLM_L_X10Y102_SLICE_X13Y102_BO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A5 = CLBLM_R_X11Y104_SLICE_X14Y104_BO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_A6 = CLBLM_R_X11Y104_SLICE_X15Y104_CO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B1 = CLBLM_L_X10Y105_SLICE_X12Y105_BO5;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B2 = CLBLM_L_X10Y102_SLICE_X13Y102_BO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B3 = CLBLM_L_X10Y105_SLICE_X13Y105_AO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B4 = CLBLM_L_X10Y102_SLICE_X13Y102_DO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B5 = CLBLM_R_X11Y104_SLICE_X14Y104_BO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_B6 = CLBLM_R_X11Y104_SLICE_X15Y104_CO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C1 = CLBLM_R_X11Y104_SLICE_X14Y104_BO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C5 = CLBLM_R_X11Y104_SLICE_X15Y104_CO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_C6 = CLBLM_L_X10Y102_SLICE_X13Y102_DO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D1 = CLBLM_L_X10Y106_SLICE_X12Y106_CO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D2 = CLBLM_R_X11Y104_SLICE_X14Y104_DO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D3 = CLBLM_L_X10Y103_SLICE_X13Y103_DO6;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D4 = CLBLM_L_X10Y105_SLICE_X13Y105_AO5;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D5 = CLBLM_L_X10Y102_SLICE_X13Y102_BO5;
  assign CLBLM_L_X10Y104_SLICE_X13Y104_D6 = CLBLM_R_X11Y104_SLICE_X14Y104_CO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A1 = CLBLM_L_X10Y104_SLICE_X13Y104_CO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_A6 = CLBLM_R_X11Y105_SLICE_X14Y105_BO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B1 = CLBLM_L_X10Y105_SLICE_X12Y105_AO5;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B2 = CLBLM_L_X8Y102_SLICE_X11Y102_BO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B3 = CLBLM_L_X10Y104_SLICE_X13Y104_AO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B4 = CLBLM_L_X10Y105_SLICE_X12Y105_BO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B5 = CLBLM_L_X10Y102_SLICE_X12Y102_AO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_B6 = CLBLM_L_X10Y102_SLICE_X12Y102_CO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C2 = CLBLM_L_X10Y104_SLICE_X13Y104_AO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C5 = CLBLM_L_X10Y102_SLICE_X12Y102_DO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_C6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D1 = CLBLM_L_X10Y102_SLICE_X12Y102_AO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D2 = CLBLM_L_X10Y104_SLICE_X13Y104_AO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D3 = CLBLM_L_X10Y104_SLICE_X13Y104_BO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D4 = CLBLM_R_X11Y105_SLICE_X14Y105_BO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D5 = CLBLM_L_X8Y105_SLICE_X10Y105_AO6;
  assign CLBLM_L_X10Y104_SLICE_X12Y104_D6 = CLBLM_L_X10Y105_SLICE_X12Y105_BO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A1 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A2 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_A6 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B5 = CLBLM_R_X11Y106_SLICE_X15Y106_DO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_B6 = CLBLM_R_X11Y105_SLICE_X15Y105_DO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C2 = CLBLM_L_X8Y102_SLICE_X10Y102_CO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C3 = CLBLM_R_X11Y106_SLICE_X15Y106_DO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C4 = CLBLM_R_X11Y105_SLICE_X15Y105_DO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_C6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D2 = CLBLM_L_X10Y104_SLICE_X13Y104_CO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D3 = CLBLM_R_X11Y104_SLICE_X14Y104_AO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D4 = CLBLM_L_X10Y105_SLICE_X13Y105_CO6;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y105_SLICE_X13Y105_D6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A1 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A5 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_A6 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B1 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B4 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_B6 = 1'b1;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C1 = CLBLM_L_X10Y105_SLICE_X12Y105_AO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C2 = CLBLM_L_X8Y105_SLICE_X10Y105_AO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C3 = CLBLM_R_X11Y105_SLICE_X14Y105_CO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C4 = CLBLM_L_X10Y104_SLICE_X13Y104_BO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C5 = CLBLM_R_X11Y107_SLICE_X15Y107_BO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_C6 = CLBLM_R_X11Y105_SLICE_X14Y105_BO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D2 = CLBLM_L_X10Y104_SLICE_X13Y104_CO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D4 = CLBLM_R_X11Y105_SLICE_X14Y105_BO6;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y105_SLICE_X12Y105_D6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_A1 = CLBLM_R_X5Y101_SLICE_X7Y101_CO6;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_A2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_A3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_A4 = CLBLM_R_X5Y101_SLICE_X7Y101_AO5;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_A5 = CLBLM_R_X5Y100_SLICE_X6Y100_AO6;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_A6 = 1'b1;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_B1 = CLBLM_R_X5Y101_SLICE_X7Y101_CO6;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_B3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_B4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_B5 = CLBLL_L_X4Y101_SLICE_X5Y101_BO6;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_B6 = CLBLL_L_X4Y101_SLICE_X4Y101_AO5;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_C1 = CLBLL_L_X4Y101_SLICE_X5Y101_BO6;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_C2 = CLBLM_R_X5Y101_SLICE_X7Y101_CO6;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_C3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_C4 = CLBLL_L_X4Y101_SLICE_X4Y101_AO5;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_C6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_D1 = 1'b1;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_D2 = 1'b1;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_D3 = 1'b1;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_D4 = 1'b1;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_D5 = 1'b1;
  assign CLBLL_L_X4Y101_SLICE_X4Y101_D6 = 1'b1;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_A1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_A2 = CLBLM_R_X5Y101_SLICE_X7Y101_AO5;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_A3 = CLBLM_R_X5Y100_SLICE_X6Y100_AO6;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_A4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_A5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_A6 = CLBLL_L_X4Y101_SLICE_X5Y101_CO6;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_B1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_B2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_B3 = CLBLM_R_X5Y100_SLICE_X6Y100_AO6;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_B4 = CLBLM_R_X5Y101_SLICE_X7Y101_AO5;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_B5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_B6 = CLBLL_L_X4Y101_SLICE_X5Y101_CO6;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_C1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_C2 = CLBLM_R_X5Y101_SLICE_X6Y101_BO6;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_C3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_C4 = CLBLM_R_X5Y101_SLICE_X7Y101_DO6;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_C5 = CLBLM_R_X5Y101_SLICE_X6Y101_CO6;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_C6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_D1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_D2 = CLBLM_R_X5Y101_SLICE_X6Y101_BO6;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_D3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_D4 = CLBLM_R_X5Y101_SLICE_X7Y101_DO6;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_D5 = CLBLM_R_X5Y101_SLICE_X6Y101_CO6;
  assign CLBLL_L_X4Y101_SLICE_X5Y101_D6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A1 = CLBLM_L_X10Y107_SLICE_X13Y107_AO5;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A2 = CLBLM_L_X10Y106_SLICE_X12Y106_DO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A3 = CLBLM_L_X10Y106_SLICE_X12Y106_CO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A4 = CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A5 = CLBLM_L_X10Y105_SLICE_X13Y105_AO5;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_A6 = CLBLM_R_X11Y104_SLICE_X14Y104_CO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B2 = CLBLM_R_X11Y105_SLICE_X14Y105_CO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B5 = CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_B6 = CLBLM_L_X10Y105_SLICE_X13Y105_BO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C1 = CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C2 = CLBLM_R_X11Y105_SLICE_X14Y105_CO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_C6 = CLBLM_L_X10Y105_SLICE_X13Y105_BO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D1 = CLBLM_R_X11Y106_SLICE_X14Y106_BO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D5 = CLBLM_R_X11Y105_SLICE_X14Y105_DO6;
  assign CLBLM_L_X10Y106_SLICE_X13Y106_D6 = CLBLM_L_X10Y105_SLICE_X13Y105_BO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A2 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A4 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_A6 = 1'b1;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_B6 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C1 = CLBLM_L_X10Y106_SLICE_X12Y106_AO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C2 = CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C3 = CLBLM_R_X11Y105_SLICE_X15Y105_AO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C4 = CLBLM_L_X10Y106_SLICE_X12Y106_AO5;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C5 = CLBLM_R_X11Y104_SLICE_X15Y104_AO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_C6 = CLBLM_R_X11Y105_SLICE_X15Y105_BO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D1 = CLBLM_L_X10Y106_SLICE_X12Y106_AO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D2 = CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D3 = CLBLM_R_X11Y105_SLICE_X15Y105_AO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D4 = CLBLM_L_X10Y106_SLICE_X12Y106_AO5;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D5 = CLBLM_R_X11Y104_SLICE_X15Y104_AO6;
  assign CLBLM_L_X10Y106_SLICE_X12Y106_D6 = CLBLM_R_X11Y105_SLICE_X15Y105_BO6;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_A1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_A2 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_A3 = CLBLL_L_X4Y102_SLICE_X5Y102_AO6;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_A4 = CLBLL_L_X4Y101_SLICE_X5Y101_DO6;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_A5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_A6 = 1'b1;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_B1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_B2 = CLBLL_L_X4Y103_SLICE_X5Y103_BO6;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_B3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_B4 = CLBLM_R_X3Y102_SLICE_X2Y102_BO6;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_B5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_B6 = CLBLM_R_X5Y101_SLICE_X6Y101_AO5;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_C1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_C2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_C3 = CLBLL_L_X4Y103_SLICE_X5Y103_BO6;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_C4 = CLBLM_R_X5Y101_SLICE_X6Y101_AO5;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_C5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_C6 = CLBLM_R_X3Y102_SLICE_X2Y102_BO6;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_D1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_D2 = CLBLL_L_X4Y102_SLICE_X5Y102_AO6;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_D3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_D4 = CLBLL_L_X4Y102_SLICE_X4Y102_CO6;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_D5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y102_SLICE_X4Y102_D6 = CLBLL_L_X4Y101_SLICE_X5Y101_DO6;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_A1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_A2 = CLBLM_R_X5Y101_SLICE_X6Y101_AO5;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_A3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_A4 = CLBLL_L_X4Y102_SLICE_X5Y102_BO6;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_A5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_A6 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_B1 = CLBLM_R_X3Y102_SLICE_X3Y102_BO6;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_B2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_B3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_B4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_B5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_B6 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_C1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_C2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_C3 = CLBLM_R_X3Y102_SLICE_X3Y102_BO6;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_C4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_C5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_C6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_D1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_D2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_D3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_D4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_D5 = CLBLM_R_X5Y102_SLICE_X6Y102_CO6;
  assign CLBLL_L_X4Y102_SLICE_X5Y102_D6 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A1 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A3 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_A6 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_B6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C1 = CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C2 = CLBLM_L_X10Y106_SLICE_X12Y106_AO5;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C3 = CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C4 = CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C5 = CLBLM_R_X5Y109_SLICE_X7Y109_AO5;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_C6 = CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D1 = CLBLM_L_X10Y107_SLICE_X13Y107_AO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D2 = CLBLM_L_X10Y106_SLICE_X12Y106_AO5;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D3 = CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D4 = CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D5 = CLBLM_R_X5Y109_SLICE_X7Y109_AO5;
  assign CLBLM_L_X10Y107_SLICE_X13Y107_D6 = CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A2 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A5 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_A6 = 1'b1;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B1 = CLBLM_R_X11Y105_SLICE_X14Y105_CO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B2 = CLBLM_R_X11Y107_SLICE_X15Y107_DO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B3 = CLBLM_L_X10Y105_SLICE_X12Y105_AO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B4 = CLBLM_R_X11Y107_SLICE_X15Y107_BO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B5 = CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_B6 = CLBLM_L_X10Y107_SLICE_X12Y107_AO5;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C1 = CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C2 = CLBLM_R_X11Y107_SLICE_X15Y107_CO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_C6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D1 = CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D2 = CLBLM_R_X11Y107_SLICE_X15Y107_CO6;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y107_SLICE_X12Y107_D6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A1 = CLBLL_L_X2Y103_SLICE_X1Y103_BO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A2 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A4 = CLBLL_L_X4Y102_SLICE_X4Y102_DO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A6 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B2 = CLBLL_L_X4Y102_SLICE_X4Y102_AO5;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B5 = CLBLL_L_X4Y101_SLICE_X5Y101_AO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B6 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C1 = CLBLL_L_X4Y104_SLICE_X5Y104_AO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C4 = CLBLM_R_X5Y104_SLICE_X6Y104_AO5;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C6 = CLBLL_L_X4Y104_SLICE_X5Y104_BO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D2 = CLBLL_L_X4Y101_SLICE_X5Y101_DO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D4 = CLBLL_L_X4Y102_SLICE_X4Y102_CO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D5 = CLBLL_L_X4Y102_SLICE_X5Y102_AO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A1 = CLBLM_R_X5Y104_SLICE_X6Y104_AO5;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A3 = CLBLL_L_X4Y104_SLICE_X5Y104_AO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A5 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A6 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B1 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B2 = CLBLL_L_X4Y102_SLICE_X5Y102_BO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B6 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C4 = CLBLL_L_X4Y103_SLICE_X5Y103_AO5;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C6 = CLBLL_L_X4Y104_SLICE_X5Y104_BO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D1 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D2 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D3 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D4 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D5 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D6 = 1'b1;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A1 = CLBLM_L_X10Y109_SLICE_X12Y109_AO5;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A2 = CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A3 = CLBLM_R_X11Y107_SLICE_X15Y107_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A4 = CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A5 = CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_A6 = CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B1 = CLBLM_L_X10Y109_SLICE_X12Y109_AO5;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B2 = CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B3 = CLBLM_R_X11Y107_SLICE_X15Y107_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B4 = CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B5 = CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_B6 = CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C1 = CLBLM_L_X10Y107_SLICE_X13Y107_AO5;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C2 = CLBLM_R_X11Y107_SLICE_X15Y107_AO5;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C3 = CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C4 = CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C5 = CLBLM_L_X10Y106_SLICE_X12Y106_DO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_C6 = CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D1 = CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D2 = CLBLM_L_X10Y109_SLICE_X12Y109_AO5;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D3 = CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D4 = CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D5 = CLBLM_R_X11Y107_SLICE_X15Y107_AO6;
  assign CLBLM_L_X10Y108_SLICE_X13Y108_D6 = CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A4 = CLBLM_L_X10Y110_SLICE_X12Y110_BO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_A6 = CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B1 = CLBLM_R_X11Y107_SLICE_X15Y107_DO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B2 = CLBLM_L_X10Y108_SLICE_X13Y108_DO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B3 = CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B4 = CLBLM_L_X10Y110_SLICE_X12Y110_BO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B5 = CLBLM_L_X10Y107_SLICE_X12Y107_AO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_B6 = CLBLM_L_X10Y107_SLICE_X12Y107_AO5;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C4 = CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_C6 = CLBLM_L_X10Y110_SLICE_X12Y110_BO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D3 = CLBLM_R_X11Y108_SLICE_X14Y108_CO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D4 = CLBLM_R_X11Y108_SLICE_X14Y108_BO6;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y108_SLICE_X12Y108_D6 = CLBLM_L_X10Y111_SLICE_X13Y111_AO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A1 = CLBLM_R_X5Y105_SLICE_X7Y105_BO5;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A3 = CLBLL_L_X4Y101_SLICE_X4Y101_AO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A5 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A6 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B1 = CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B2 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B5 = CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B6 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C1 = CLBLL_L_X4Y101_SLICE_X4Y101_BO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C2 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C4 = CLBLL_L_X4Y104_SLICE_X4Y104_AO5;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C5 = CLBLM_R_X5Y105_SLICE_X7Y105_BO5;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D1 = CLBLL_L_X4Y101_SLICE_X4Y101_BO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D2 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D4 = CLBLL_L_X4Y104_SLICE_X4Y104_AO5;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D5 = CLBLM_R_X5Y105_SLICE_X7Y105_BO5;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A1 = CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A2 = CLBLM_R_X5Y103_SLICE_X6Y103_AO5;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A5 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A6 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B1 = CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B2 = CLBLM_R_X5Y103_SLICE_X6Y103_AO5;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B4 = CLBLM_R_X5Y102_SLICE_X6Y102_AO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C1 = CLBLL_L_X4Y106_SLICE_X5Y106_AO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C2 = CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C3 = CLBLM_R_X5Y103_SLICE_X6Y103_AO5;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C4 = CLBLL_L_X4Y104_SLICE_X5Y104_AO5;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C5 = CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C6 = CLBLM_R_X5Y102_SLICE_X6Y102_AO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C3 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D1 = CLBLL_L_X4Y104_SLICE_X5Y104_AO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D2 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D4 = CLBLL_L_X4Y104_SLICE_X5Y104_CO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D6 = CLBLM_R_X5Y104_SLICE_X6Y104_AO5;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D3 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D4 = 1'b1;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_D = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_D = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A1 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A2 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_A6 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B1 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B3 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_B6 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C1 = CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C2 = CLBLM_R_X11Y108_SLICE_X15Y108_AO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C3 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C4 = CLBLM_R_X5Y109_SLICE_X7Y109_AO5;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C5 = CLBLM_L_X10Y109_SLICE_X13Y109_BO5;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_C6 = CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D1 = CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D2 = CLBLM_R_X11Y108_SLICE_X15Y108_AO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D3 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D4 = CLBLM_R_X5Y109_SLICE_X7Y109_AO5;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D5 = CLBLM_L_X10Y109_SLICE_X13Y109_BO5;
  assign CLBLM_L_X10Y109_SLICE_X13Y109_D6 = CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A4 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A5 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_A6 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C3 = 1'b1;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_B6 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C1 = CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C2 = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C3 = CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C4 = CLBLM_R_X11Y107_SLICE_X15Y107_AO5;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C5 = CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_C6 = CLBLM_L_X10Y107_SLICE_X13Y107_DO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D3 = CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y109_SLICE_X12Y109_D6 = CLBLM_R_X11Y109_SLICE_X14Y109_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A2 = CLBLM_R_X5Y103_SLICE_X6Y103_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A6 = CLBLL_L_X4Y103_SLICE_X4Y103_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B2 = CLBLM_R_X3Y105_SLICE_X3Y105_AO5;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B6 = CLBLL_L_X4Y103_SLICE_X5Y103_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C1 = CLBLL_L_X4Y104_SLICE_X4Y104_AO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C3 = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D1 = CLBLL_L_X4Y105_SLICE_X4Y105_AO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D2 = CLBLL_L_X4Y105_SLICE_X5Y105_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D3 = CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D4 = CLBLM_R_X3Y105_SLICE_X3Y105_DO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D5 = CLBLL_L_X4Y104_SLICE_X4Y104_BO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D6 = CLBLL_L_X4Y105_SLICE_X4Y105_BO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D3 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D4 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_A1 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_A2 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_A3 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_A4 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_A5 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_A6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_D1 = CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_B1 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_B2 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_B3 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_B4 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_B5 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A2 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_C1 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_C2 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_C3 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A5 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_C5 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A6 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B1 = CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B4 = CLBLM_R_X5Y103_SLICE_X6Y103_AO5;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B6 = CLBLM_R_X5Y105_SLICE_X7Y105_BO6;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_D1 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_D2 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_D3 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_D4 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_D5 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_D6 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C1 = CLBLM_R_X3Y106_SLICE_X3Y106_AO5;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C2 = CLBLM_R_X5Y103_SLICE_X6Y103_DO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C3 = CLBLL_L_X4Y104_SLICE_X5Y104_DO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C4 = CLBLL_L_X4Y105_SLICE_X5Y105_AO5;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C5 = CLBLL_L_X4Y105_SLICE_X5Y105_AO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C6 = CLBLM_R_X5Y103_SLICE_X6Y103_CO6;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_A1 = CLBLM_R_X11Y104_SLICE_X14Y104_DO6;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_A2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_A3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_A4 = CLBLM_L_X10Y103_SLICE_X13Y103_CO6;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_A5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D1 = CLBLM_R_X3Y106_SLICE_X3Y106_AO5;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D2 = CLBLM_R_X5Y103_SLICE_X6Y103_DO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D3 = CLBLL_L_X4Y104_SLICE_X5Y104_DO6;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_B1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_B2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_B3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D5 = CLBLL_L_X4Y105_SLICE_X5Y105_AO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D6 = CLBLM_R_X5Y103_SLICE_X6Y103_CO6;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_B5 = CLBLM_R_X11Y104_SLICE_X15Y104_DO6;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_B6 = CLBLM_R_X11Y104_SLICE_X15Y104_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_C1 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_C2 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_C3 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_C4 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_C5 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_C6 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D5 = CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_D1 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_D2 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_D3 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_D4 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_D5 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X14Y103_D6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_D1 = CLBLL_L_X4Y107_SLICE_X4Y107_AO5;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C1 = CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C2 = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C3 = CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A2 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A3 = CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A5 = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_A6 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B1 = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B2 = CLBLM_R_X11Y110_SLICE_X14Y110_AO5;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B3 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B4 = CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B5 = CLBLM_R_X11Y110_SLICE_X14Y110_AO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_B6 = CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C2 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C3 = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C5 = CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_C6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D1 = CLBLM_R_X11Y110_SLICE_X14Y110_AO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D2 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D3 = CLBLM_R_X11Y110_SLICE_X14Y110_AO5;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D4 = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D5 = CLBLM_R_X11Y109_SLICE_X15Y109_AO6;
  assign CLBLM_L_X10Y110_SLICE_X13Y110_D6 = CLBLM_L_X10Y109_SLICE_X13Y109_BO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A1 = CLBLM_L_X10Y111_SLICE_X12Y111_AO5;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A2 = CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A3 = CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A4 = CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A5 = CLBLM_L_X10Y109_SLICE_X13Y109_AO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_A6 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B1 = CLBLM_L_X10Y111_SLICE_X12Y111_AO5;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B2 = CLBLM_L_X8Y109_SLICE_X11Y109_AO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B3 = CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B4 = CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B5 = CLBLM_L_X10Y109_SLICE_X13Y109_AO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_B6 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C2 = CLBLM_L_X10Y109_SLICE_X12Y109_CO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C5 = CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_C6 = CLBLM_L_X10Y109_SLICE_X12Y109_DO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D4 = CLBLM_R_X5Y112_SLICE_X6Y112_AO5;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A1 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A3 = CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A4 = CLBLM_R_X5Y105_SLICE_X6Y105_CO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A6 = 1'b1;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D1 = CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D2 = CLBLM_L_X10Y109_SLICE_X13Y109_CO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D3 = CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B1 = CLBLL_L_X4Y107_SLICE_X4Y107_DO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B2 = CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B3 = CLBLL_L_X4Y106_SLICE_X5Y106_DO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B4 = CLBLM_R_X3Y105_SLICE_X3Y105_DO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B5 = CLBLL_L_X4Y105_SLICE_X4Y105_AO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B6 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C2 = CLBLM_R_X5Y103_SLICE_X6Y103_CO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C6 = CLBLL_L_X4Y103_SLICE_X4Y103_CO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D1 = CLBLM_R_X5Y103_SLICE_X6Y103_CO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D2 = CLBLM_R_X3Y105_SLICE_X3Y105_DO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D3 = CLBLL_L_X4Y106_SLICE_X5Y106_DO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D4 = CLBLL_L_X4Y104_SLICE_X5Y104_DO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D5 = CLBLL_L_X4Y107_SLICE_X4Y107_DO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D6 = CLBLL_L_X4Y105_SLICE_X5Y105_AO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_A1 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_A2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_A4 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_A6 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A1 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A2 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A6 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_B1 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_B2 = CLBLM_L_X12Y104_SLICE_X16Y104_CO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_B3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B4 = CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B6 = CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_C2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C3 = CLBLM_R_X3Y106_SLICE_X3Y106_AO5;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C6 = CLBLM_R_X5Y104_SLICE_X6Y104_BO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_D2 = CLBLM_L_X10Y103_SLICE_X13Y103_CO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_D3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_D4 = CLBLM_L_X10Y103_SLICE_X13Y103_AO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_D5 = CLBLM_R_X11Y104_SLICE_X15Y104_BO5;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_D6 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D3 = CLBLM_R_X3Y106_SLICE_X3Y106_AO5;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D6 = CLBLM_R_X5Y104_SLICE_X6Y104_BO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_A1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_A2 = CLBLM_R_X11Y104_SLICE_X15Y104_DO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_A4 = CLBLM_R_X11Y104_SLICE_X15Y104_CO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_A5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_A6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_B1 = CLBLM_R_X11Y104_SLICE_X14Y104_DO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_B2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_B4 = CLBLM_L_X10Y103_SLICE_X13Y103_CO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_B5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_B6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_C1 = CLBLM_R_X11Y105_SLICE_X15Y105_AO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_C2 = CLBLM_R_X11Y104_SLICE_X15Y104_AO5;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_C3 = CLBLL_L_X4Y103_SLICE_X4Y103_BO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_C4 = CLBLM_L_X12Y104_SLICE_X16Y104_BO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_C5 = CLBLM_R_X11Y104_SLICE_X15Y104_AO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_C6 = CLBLM_L_X12Y104_SLICE_X16Y104_CO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_D1 = CLBLM_R_X11Y105_SLICE_X15Y105_AO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_D2 = CLBLM_R_X11Y104_SLICE_X15Y104_AO5;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_D3 = CLBLL_L_X4Y103_SLICE_X4Y103_BO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_D4 = CLBLM_L_X12Y104_SLICE_X16Y104_BO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_D5 = CLBLM_R_X11Y104_SLICE_X15Y104_AO6;
  assign CLBLM_R_X11Y104_SLICE_X14Y104_D6 = CLBLM_L_X12Y104_SLICE_X16Y104_CO6;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_B5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A4 = CLBLM_R_X11Y110_SLICE_X14Y110_BO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A5 = CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_A6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B1 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B2 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B3 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B4 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B5 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_B6 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_A1 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_A2 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_A3 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_A4 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_A5 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C6 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_A6 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C1 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C2 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_B1 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_B2 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_B3 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_B4 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_B5 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_B6 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D2 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D3 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D5 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D6 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_C1 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_C2 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_C3 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_C4 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_C5 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_C6 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A1 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A4 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_A6 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_D1 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_D2 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_D3 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_D4 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_D5 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X11Y101_D6 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B2 = CLBLM_L_X8Y112_SLICE_X11Y112_AO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B5 = CLBLM_L_X10Y110_SLICE_X13Y110_AO6;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_A1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_A2 = CLBLM_L_X8Y103_SLICE_X10Y103_BO6;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_A3 = CLBLM_R_X7Y101_SLICE_X9Y101_BO6;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_A4 = CLBLM_L_X10Y101_SLICE_X12Y101_BO6;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_A5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_A6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C2 = CLBLM_R_X11Y110_SLICE_X14Y110_BO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_B1 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_B2 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A1 = CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A2 = CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A3 = CLBLM_R_X3Y107_SLICE_X3Y107_BO6;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_B6 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A4 = CLBLL_L_X4Y106_SLICE_X5Y106_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A5 = CLBLL_L_X4Y106_SLICE_X5Y106_BO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A6 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_B3 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_C1 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_C2 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_C3 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_C4 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_C5 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_C6 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B1 = CLBLM_R_X5Y107_SLICE_X6Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B4 = CLBLM_R_X3Y107_SLICE_X3Y107_DO5;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C2 = CLBLM_R_X5Y107_SLICE_X6Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C3 = CLBLM_R_X3Y107_SLICE_X3Y107_DO5;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_D1 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_D2 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_D3 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_D4 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_D5 = 1'b1;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_D6 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D1 = CLBLL_L_X4Y106_SLICE_X5Y106_BO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D2 = CLBLL_L_X4Y107_SLICE_X5Y107_AO5;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D3 = CLBLM_R_X5Y107_SLICE_X6Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D4 = CLBLM_R_X3Y107_SLICE_X3Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D5 = CLBLM_R_X3Y107_SLICE_X2Y107_AO5;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D6 = CLBLL_L_X4Y106_SLICE_X5Y106_CO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A1 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A3 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A6 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_A6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B2 = CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B6 = CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C2 = CLBLM_R_X5Y107_SLICE_X7Y107_AO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C3 = CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C6 = CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C3 = CLBLM_L_X10Y106_SLICE_X12Y106_CO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C6 = CLBLM_L_X12Y104_SLICE_X16Y104_AO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D1 = CLBLM_L_X12Y104_SLICE_X16Y104_AO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D1 = CLBLL_L_X4Y106_SLICE_X5Y106_CO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D2 = CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D3 = CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D4 = CLBLL_L_X4Y105_SLICE_X5Y105_DO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D5 = CLBLL_L_X4Y106_SLICE_X5Y106_BO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D6 = CLBLM_R_X3Y107_SLICE_X3Y107_BO6;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D4 = CLBLM_R_X11Y106_SLICE_X15Y106_AO5;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_D6 = CLBLM_R_X11Y104_SLICE_X15Y104_BO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A1 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A2 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_A6 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B1 = CLBLM_R_X11Y106_SLICE_X15Y106_DO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B2 = CLBLM_L_X10Y104_SLICE_X13Y104_DO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B3 = CLBLM_R_X11Y105_SLICE_X15Y105_CO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B4 = CLBLM_L_X10Y105_SLICE_X13Y105_AO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B5 = CLBLM_R_X11Y105_SLICE_X14Y105_AO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_B6 = CLBLM_R_X11Y105_SLICE_X14Y105_AO5;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C1 = CLBLM_R_X11Y105_SLICE_X14Y105_AO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C2 = CLBLM_R_X11Y105_SLICE_X15Y105_CO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C3 = CLBLM_L_X10Y104_SLICE_X13Y104_DO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C4 = CLBLM_R_X11Y105_SLICE_X14Y105_AO5;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C5 = CLBLM_R_X11Y106_SLICE_X15Y106_DO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_C6 = CLBLM_L_X10Y105_SLICE_X13Y105_AO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D1 = CLBLM_L_X10Y104_SLICE_X13Y104_DO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D2 = CLBLM_R_X11Y105_SLICE_X15Y105_CO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D5 = CLBLM_R_X11Y106_SLICE_X15Y106_DO6;
  assign CLBLM_R_X11Y105_SLICE_X14Y105_D6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_A1 = CLBLM_R_X7Y101_SLICE_X9Y101_CO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_A2 = CLBLM_L_X10Y101_SLICE_X13Y101_AO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_A4 = 1'b1;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_A5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_A6 = 1'b1;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_B1 = CLBLM_L_X8Y102_SLICE_X11Y102_DO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_B2 = CLBLM_L_X8Y103_SLICE_X10Y103_BO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_B3 = CLBLM_L_X8Y102_SLICE_X10Y102_AO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_B4 = CLBLM_R_X7Y102_SLICE_X9Y102_CO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_B5 = CLBLM_L_X10Y101_SLICE_X12Y101_BO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_B6 = CLBLM_L_X10Y102_SLICE_X13Y102_AO5;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_C1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_C2 = CLBLM_L_X8Y102_SLICE_X10Y102_CO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_C3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_C4 = CLBLM_L_X10Y101_SLICE_X13Y101_AO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_C5 = CLBLM_R_X7Y101_SLICE_X9Y101_CO6;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_C6 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_D1 = 1'b1;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_D2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_D3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_D4 = 1'b1;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_D5 = 1'b1;
  assign CLBLM_L_X8Y102_SLICE_X11Y102_D6 = 1'b1;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_A1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_A2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_A3 = CLBLM_L_X10Y101_SLICE_X12Y101_BO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_A4 = CLBLM_L_X8Y103_SLICE_X10Y103_BO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_A5 = 1'b1;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_A6 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A3 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A5 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A6 = 1'b1;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_B1 = CLBLM_L_X8Y102_SLICE_X10Y102_DO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_B2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B1 = CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B2 = CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B3 = CLBLM_R_X3Y105_SLICE_X3Y105_AO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B4 = CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B5 = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B6 = CLBLL_L_X4Y108_SLICE_X4Y108_AO5;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_B5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_B6 = CLBLM_L_X8Y102_SLICE_X10Y102_AO5;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C4 = CLBLM_R_X7Y108_SLICE_X8Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C5 = CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_C4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_C5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_C6 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_D1 = CLBLM_R_X7Y102_SLICE_X9Y102_CO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_D2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_D3 = CLBLM_L_X10Y101_SLICE_X12Y101_BO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_D4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D3 = CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D4 = CLBLM_R_X7Y108_SLICE_X8Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_D6 = CLBLM_L_X8Y103_SLICE_X10Y103_BO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A3 = CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A4 = CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A5 = CLBLM_R_X5Y107_SLICE_X7Y107_AO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A3 = CLBLM_R_X11Y105_SLICE_X15Y105_BO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B1 = CLBLM_R_X3Y102_SLICE_X3Y102_AO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B2 = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B3 = CLBLL_L_X4Y107_SLICE_X5Y107_AO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B4 = CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B5 = CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B6 = CLBLM_R_X5Y108_SLICE_X6Y108_BO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C5 = CLBLL_L_X4Y108_SLICE_X5Y108_DO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C6 = CLBLM_R_X5Y108_SLICE_X6Y108_CO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C3 = CLBLM_R_X11Y106_SLICE_X14Y106_DO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C4 = CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_C6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D2 = CLBLM_R_X5Y107_SLICE_X7Y107_CO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D5 = CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D6 = CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D3 = CLBLM_R_X11Y106_SLICE_X14Y106_DO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D4 = CLBLM_L_X10Y107_SLICE_X13Y107_CO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_D6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_A6 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B4 = CLBLM_R_X11Y108_SLICE_X15Y108_BO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_B6 = CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C2 = CLBLM_R_X11Y106_SLICE_X15Y106_AO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C3 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C4 = CLBLM_R_X11Y107_SLICE_X14Y107_AO5;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C5 = CLBLM_R_X11Y106_SLICE_X14Y106_DO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_C6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D1 = CLBLM_R_X11Y105_SLICE_X15Y105_BO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D2 = CLBLM_R_X11Y105_SLICE_X15Y105_AO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D3 = CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y106_SLICE_X14Y106_D6 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B5 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B6 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A1 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A2 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A3 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A4 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A5 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_A6 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B1 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B2 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B3 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B4 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B5 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_B6 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C1 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C2 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C3 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C4 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C5 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_C6 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D1 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D2 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D3 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D4 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D5 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X11Y103_D6 = 1'b1;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A1 = CLBLM_L_X8Y102_SLICE_X10Y102_DO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A3 = CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A4 = CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_A4 = CLBLM_L_X10Y102_SLICE_X12Y102_CO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B3 = CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B5 = CLBLM_L_X8Y102_SLICE_X11Y102_AO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_B6 = CLBLM_L_X8Y103_SLICE_X10Y103_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B1 = CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B5 = CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B6 = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C3 = CLBLM_R_X5Y109_SLICE_X6Y109_AO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C4 = CLBLM_R_X7Y109_SLICE_X8Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C6 = CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C3 = CLBLM_L_X8Y104_SLICE_X10Y104_DO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C4 = CLBLM_L_X8Y104_SLICE_X10Y104_CO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_C5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D1 = CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D5 = CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D6 = CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D1 = CLBLM_R_X7Y107_SLICE_X9Y107_BO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D2 = CLBLM_L_X8Y102_SLICE_X11Y102_AO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D4 = CLBLM_L_X8Y103_SLICE_X10Y103_CO6;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y103_SLICE_X10Y103_D6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A2 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A5 = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A6 = CLBLM_R_X5Y109_SLICE_X6Y109_BO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A1 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A2 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B2 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B3 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B4 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B5 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B6 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_A6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C2 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C3 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C4 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C5 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C6 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B3 = CLBLM_R_X11Y105_SLICE_X14Y105_AO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B4 = CLBLM_R_X11Y106_SLICE_X15Y106_CO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B5 = CLBLM_R_X11Y107_SLICE_X15Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B6 = CLBLM_L_X10Y109_SLICE_X13Y109_AO5;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C1 = CLBLM_R_X11Y107_SLICE_X15Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C2 = CLBLM_R_X11Y105_SLICE_X14Y105_AO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C3 = CLBLM_R_X11Y106_SLICE_X15Y106_DO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D2 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D3 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D4 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D5 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D6 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D1 = CLBLM_R_X11Y107_SLICE_X15Y107_AO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D2 = CLBLM_R_X11Y105_SLICE_X14Y105_AO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D3 = CLBLM_L_X10Y109_SLICE_X13Y109_AO5;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D4 = CLBLM_R_X11Y108_SLICE_X15Y108_BO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D5 = CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_D6 = CLBLM_R_X11Y106_SLICE_X15Y106_CO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A2 = CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A3 = CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A4 = 1'b1;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_A6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C3 = 1'b1;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_D = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B3 = CLBLM_R_X11Y107_SLICE_X15Y107_CO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B4 = CLBLM_R_X11Y108_SLICE_X14Y108_AO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_B6 = CLBLM_R_X11Y107_SLICE_X14Y107_CO6;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_D = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C2 = CLBLM_R_X11Y106_SLICE_X14Y106_CO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_C6 = CLBLM_R_X11Y108_SLICE_X15Y108_BO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D2 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D4 = CLBLM_L_X10Y107_SLICE_X13Y107_BO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D5 = CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  assign CLBLM_R_X11Y107_SLICE_X14Y107_D6 = CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D3 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D4 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A2 = CLBLM_L_X10Y103_SLICE_X12Y103_BO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A4 = CLBLM_L_X10Y104_SLICE_X12Y104_AO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_A6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B2 = CLBLM_L_X10Y103_SLICE_X12Y103_BO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B5 = CLBLM_L_X10Y104_SLICE_X12Y104_AO6;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_B6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C1 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C2 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C3 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C4 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C5 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_C6 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D1 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D2 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D3 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D4 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D5 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X11Y104_D6 = 1'b1;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A1 = CLBLM_L_X8Y104_SLICE_X10Y104_DO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A2 = CLBLM_L_X8Y102_SLICE_X10Y102_CO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_A6 = CLBLM_L_X8Y104_SLICE_X10Y104_CO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B3 = CLBLM_L_X10Y104_SLICE_X12Y104_AO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B5 = CLBLM_L_X10Y104_SLICE_X12Y104_CO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_B6 = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_C6 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X8Y104_SLICE_X10Y104_D6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C1 = CLBLM_R_X7Y111_SLICE_X8Y111_AO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C2 = CLBLM_L_X8Y111_SLICE_X10Y111_DO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A3 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_A6 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B1 = CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B2 = CLBLM_R_X11Y107_SLICE_X14Y107_DO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B5 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_B6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C2 = CLBLM_R_X11Y107_SLICE_X14Y107_DO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C5 = CLBLM_L_X10Y109_SLICE_X13Y109_DO6;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_C6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D1 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D2 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D3 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D4 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D5 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X15Y108_D6 = 1'b1;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A3 = CLBLM_R_X11Y108_SLICE_X14Y108_DO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_A6 = CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B2 = CLBLM_L_X10Y108_SLICE_X13Y108_CO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B3 = CLBLM_R_X11Y108_SLICE_X15Y108_CO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_B6 = CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C3 = CLBLM_R_X11Y109_SLICE_X14Y109_BO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C5 = CLBLM_R_X11Y108_SLICE_X14Y108_DO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_C6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D1 = CLBLM_R_X11Y107_SLICE_X14Y107_AO6;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D2 = CLBLM_R_X11Y109_SLICE_X14Y109_AO5;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y108_SLICE_X14Y108_D6 = CLBLM_R_X11Y107_SLICE_X14Y107_DO6;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A1 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A2 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A3 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A4 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A5 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_A6 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B1 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B2 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B3 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B4 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B5 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_B6 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C1 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C2 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C3 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C4 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C5 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_C6 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D1 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D2 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D3 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D4 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D5 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X11Y105_D6 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A1 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A2 = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A4 = CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_A6 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A3 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A5 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A6 = 1'b1;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_A2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B6 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B1 = CLBLM_L_X10Y105_SLICE_X12Y105_DO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B2 = CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B3 = CLBLM_L_X10Y104_SLICE_X12Y104_DO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C3 = CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_B6 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C1 = CLBLL_L_X4Y111_SLICE_X4Y111_AO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C2 = CLBLM_L_X10Y105_SLICE_X13Y105_DO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C5 = CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_C6 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D2 = CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_D6 = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign RIOI3_SING_X105Y100_ILOGIC_X1Y100_D = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D2 = CLBLM_L_X10Y105_SLICE_X13Y105_DO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D5 = CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  assign CLBLM_L_X8Y105_SLICE_X10Y105_D6 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A2 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A4 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_A6 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B1 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B2 = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B3 = CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B4 = CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B5 = CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_B6 = CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C1 = CLBLL_L_X4Y111_SLICE_X5Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C2 = CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C3 = CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C4 = CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C5 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_C6 = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_A6 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B1 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B2 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B3 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_B4 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D1 = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D3 = CLBLL_L_X4Y111_SLICE_X4Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D4 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X4Y111_SLICE_X5Y111_D6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C1 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C2 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C3 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C4 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C5 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_C6 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D1 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D2 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D3 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D4 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D5 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X15Y109_D6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y137_T1 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A1 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A3 = CLBLM_R_X11Y108_SLICE_X15Y108_AO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A5 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_A6 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B1 = CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_B6 = CLBLM_R_X11Y109_SLICE_X14Y109_CO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C1 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C3 = CLBLM_L_X10Y106_SLICE_X12Y106_BO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C4 = CLBLM_R_X11Y108_SLICE_X15Y108_AO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C5 = CLBLM_R_X11Y106_SLICE_X14Y106_AO6;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_C6 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D1 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D2 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D3 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D4 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D5 = 1'b1;
  assign CLBLM_R_X11Y109_SLICE_X14Y109_D6 = 1'b1;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_D = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_D = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A1 = CLBLM_L_X10Y107_SLICE_X12Y107_DO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A2 = CLBLM_L_X8Y107_SLICE_X11Y107_AO5;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A3 = CLBLM_R_X7Y104_SLICE_X8Y104_BO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A4 = CLBLM_R_X7Y106_SLICE_X9Y106_AO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A5 = CLBLM_L_X10Y105_SLICE_X12Y105_CO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_A6 = CLBLM_L_X10Y106_SLICE_X13Y106_BO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B2 = CLBLM_L_X10Y107_SLICE_X12Y107_DO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_B6 = CLBLM_L_X10Y106_SLICE_X13Y106_DO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C1 = CLBLM_L_X10Y105_SLICE_X12Y105_CO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C4 = CLBLM_L_X10Y106_SLICE_X13Y106_BO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C5 = CLBLM_L_X10Y107_SLICE_X12Y107_DO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_C6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D1 = CLBLM_L_X10Y105_SLICE_X12Y105_CO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D5 = CLBLM_R_X7Y104_SLICE_X8Y104_BO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D6 = CLBLM_R_X7Y106_SLICE_X9Y106_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A4 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A5 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_A6 = 1'b1;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D2 = CLBLM_L_X10Y107_SLICE_X12Y107_DO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D3 = CLBLM_L_X10Y106_SLICE_X13Y106_BO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A1 = CLBLM_L_X8Y107_SLICE_X10Y107_AO5;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A2 = CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A3 = CLBLM_L_X8Y105_SLICE_X10Y105_AO5;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A4 = CLBLM_R_X7Y106_SLICE_X9Y106_AO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A5 = CLBLM_L_X10Y105_SLICE_X12Y105_DO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_A6 = CLBLM_L_X10Y104_SLICE_X12Y104_DO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B1 = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B2 = CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C1 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C3 = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C5 = CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B4 = CLBLM_L_X10Y106_SLICE_X13Y106_DO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B5 = CLBLM_L_X10Y107_SLICE_X12Y107_DO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_B6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C1 = CLBLM_L_X8Y106_SLICE_X11Y106_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D3 = CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_D6 = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C2 = CLBLM_L_X8Y106_SLICE_X11Y106_CO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C3 = CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_C5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D1 = CLBLM_L_X10Y105_SLICE_X12Y105_DO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D2 = CLBLM_L_X8Y105_SLICE_X10Y105_AO5;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D3 = CLBLM_L_X10Y106_SLICE_X13Y106_CO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D4 = CLBLM_L_X10Y104_SLICE_X12Y104_DO6;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D5 = CLBLM_L_X8Y107_SLICE_X10Y107_AO5;
  assign CLBLM_L_X8Y106_SLICE_X10Y106_D6 = CLBLM_R_X7Y106_SLICE_X9Y106_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A1 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A2 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_A6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B1 = CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B2 = CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B3 = CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B4 = CLBLL_L_X4Y111_SLICE_X5Y111_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B5 = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_B6 = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C3 = CLBLL_L_X4Y111_SLICE_X5Y111_DO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C4 = CLBLM_R_X3Y111_SLICE_X2Y111_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_C6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_B5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A1 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A2 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A3 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A4 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A5 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_A6 = 1'b1;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D1 = CLBLL_L_X4Y112_SLICE_X5Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D2 = CLBLM_R_X3Y113_SLICE_X2Y113_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D3 = CLBLL_L_X4Y112_SLICE_X4Y112_DO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D4 = CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D5 = CLBLL_L_X4Y112_SLICE_X5Y112_BO6;
  assign CLBLL_L_X4Y112_SLICE_X5Y112_D6 = CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_A1 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_A2 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_A3 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_A4 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_A5 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_A6 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C1 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_B1 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_B2 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_B3 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_B4 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_B5 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_B6 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D1 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D2 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_C1 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_C2 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_C3 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_C4 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_C5 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_C6 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D3 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D4 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A1 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A3 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A5 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C5 = CLBLM_R_X3Y111_SLICE_X2Y111_AO5;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_D1 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_D3 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_D2 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_D4 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_D6 = 1'b1;
  assign CLBLL_L_X4Y111_SLICE_X4Y111_C6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y100_SLICE_X9Y100_D5 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B1 = CLBLM_L_X10Y110_SLICE_X13Y110_AO5;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B3 = CLBLM_R_X11Y109_SLICE_X14Y109_CO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_A1 = CLBLM_R_X7Y102_SLICE_X9Y102_DO6;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_A2 = CLBLM_R_X7Y101_SLICE_X8Y101_AO5;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_A3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_A4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_A5 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_A6 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C1 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C2 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C3 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_B1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_B2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_B3 = CLBLM_R_X7Y101_SLICE_X8Y101_AO6;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_B4 = CLBLM_L_X8Y101_SLICE_X10Y101_AO6;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_B5 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_B6 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D1 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D2 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D3 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_C1 = CLBLM_R_X7Y101_SLICE_X8Y101_AO6;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_C2 = CLBLM_R_X7Y101_SLICE_X8Y101_AO5;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_C3 = CLBLM_R_X7Y102_SLICE_X9Y102_DO6;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_C4 = CLBLM_R_X7Y100_SLICE_X8Y100_AO5;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_C5 = CLBLM_R_X7Y100_SLICE_X8Y100_BO5;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_C6 = CLBLM_L_X8Y101_SLICE_X10Y101_AO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D4 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D5 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_D6 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_D1 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_D2 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_D3 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_D4 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_D5 = 1'b1;
  assign CLBLM_R_X7Y100_SLICE_X8Y100_D6 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A1 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A3 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_A6 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B1 = CLBLM_L_X10Y107_SLICE_X12Y107_CO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B2 = CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B3 = CLBLM_L_X8Y107_SLICE_X10Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B4 = CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B5 = CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_B6 = CLBLM_L_X8Y107_SLICE_X11Y107_AO5;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C1 = CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C2 = CLBLM_L_X10Y107_SLICE_X12Y107_BO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C3 = CLBLM_L_X8Y107_SLICE_X11Y107_AO5;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C4 = CLBLM_L_X10Y107_SLICE_X12Y107_CO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C5 = CLBLM_L_X8Y107_SLICE_X10Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_C6 = CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A3 = CLBLL_L_X4Y113_SLICE_X5Y113_AO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A4 = CLBLL_L_X4Y113_SLICE_X4Y113_BO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_A6 = CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D1 = CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D2 = CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B4 = CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B5 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_B6 = CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D4 = CLBLM_L_X8Y107_SLICE_X11Y107_AO5;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D5 = CLBLM_L_X10Y107_SLICE_X12Y107_CO6;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D6 = CLBLM_L_X10Y106_SLICE_X13Y106_BO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C3 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C5 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_A6 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B3 = CLBLM_R_X11Y107_SLICE_X14Y107_BO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_D6 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C1 = CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B6 = CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C4 = CLBLM_L_X8Y106_SLICE_X11Y106_BO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_C6 = CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D1 = CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D4 = CLBLM_L_X8Y106_SLICE_X11Y106_BO6;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_D6 = CLBLM_L_X8Y107_SLICE_X10Y107_BO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A3 = CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_A6 = CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B2 = CLBLL_L_X4Y112_SLICE_X5Y112_DO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B4 = CLBLM_R_X5Y112_SLICE_X6Y112_CO6;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_B6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_C6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D2 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D3 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D4 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D5 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X5Y113_D6 = 1'b1;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_A1 = CLBLM_L_X8Y103_SLICE_X10Y103_DO6;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_A2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_A3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_A4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_A5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_A6 = CLBLM_R_X7Y103_SLICE_X9Y103_AO5;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_B1 = CLBLM_L_X8Y103_SLICE_X10Y103_DO6;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_B2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_B3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_B4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_B5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_B6 = CLBLM_R_X7Y103_SLICE_X9Y103_AO5;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_C1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_C2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_C3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_C4 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_C5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_C6 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_D1 = 1'b1;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_D2 = 1'b1;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_D3 = 1'b1;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_D4 = 1'b1;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_D5 = 1'b1;
  assign CLBLM_R_X7Y101_SLICE_X9Y101_D6 = 1'b1;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_A1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_A2 = CLBLM_R_X7Y103_SLICE_X8Y103_AO6;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_A3 = CLBLM_R_X7Y101_SLICE_X9Y101_AO6;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_A5 = 1'b1;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_A6 = 1'b1;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_B1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_B2 = CLBLM_L_X8Y101_SLICE_X10Y101_AO6;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_B3 = CLBLM_L_X8Y103_SLICE_X10Y103_AO6;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_B4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_B5 = CLBLM_R_X7Y101_SLICE_X8Y101_AO6;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_B6 = 1'b1;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_C1 = 1'b1;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_C2 = CLBLM_R_X7Y100_SLICE_X8Y100_CO6;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_C3 = 1'b1;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_C4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_C5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_C6 = 1'b1;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_D1 = 1'b1;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_D2 = 1'b1;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_D3 = 1'b1;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_D4 = 1'b1;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_D5 = 1'b1;
  assign CLBLM_R_X7Y101_SLICE_X8Y101_D6 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B1 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B2 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B3 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B4 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B5 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_B6 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A1 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A2 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A3 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A4 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A5 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_A6 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B1 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B2 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B3 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B4 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B5 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_B6 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C2 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C3 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C1 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C2 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C3 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C4 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C5 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_C6 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C4 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C5 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_C6 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D1 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D2 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D3 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D4 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D5 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X11Y108_D6 = 1'b1;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A1 = CLBLM_L_X8Y109_SLICE_X10Y109_DO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A2 = CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A3 = CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A4 = CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A5 = CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_A6 = CLBLM_R_X7Y109_SLICE_X9Y109_AO5;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B1 = CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B4 = CLBLM_L_X8Y109_SLICE_X10Y109_DO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_B6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C1 = CLBLM_L_X8Y107_SLICE_X11Y107_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C2 = CLBLM_R_X7Y109_SLICE_X9Y109_AO5;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C3 = CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C4 = CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C5 = CLBLM_L_X8Y109_SLICE_X10Y109_DO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_C6 = CLBLM_R_X7Y108_SLICE_X9Y108_AO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D2 = CLBLM_L_X10Y108_SLICE_X12Y108_CO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D4 = CLBLM_L_X10Y108_SLICE_X12Y108_BO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D5 = CLBLM_L_X8Y109_SLICE_X10Y109_DO6;
  assign CLBLM_L_X8Y108_SLICE_X10Y108_D6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_D = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_D = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D5 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A6 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X15Y110_D6 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_A1 = CLBLM_L_X8Y102_SLICE_X10Y102_CO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_A2 = CLBLM_R_X5Y101_SLICE_X7Y101_AO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_A3 = CLBLM_R_X5Y101_SLICE_X6Y101_AO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_A4 = CLBLM_R_X7Y101_SLICE_X9Y101_CO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_A5 = CLBLL_L_X4Y102_SLICE_X4Y102_AO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_A6 = CLBLM_L_X10Y101_SLICE_X13Y101_AO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_B1 = CLBLM_L_X8Y102_SLICE_X10Y102_CO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_B2 = CLBLL_L_X4Y102_SLICE_X4Y102_AO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_B3 = CLBLM_R_X5Y101_SLICE_X6Y101_AO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_B4 = CLBLM_R_X7Y101_SLICE_X9Y101_CO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_B5 = CLBLM_R_X5Y101_SLICE_X7Y101_AO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_B6 = CLBLM_L_X10Y101_SLICE_X13Y101_AO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_C1 = CLBLM_R_X7Y103_SLICE_X9Y103_AO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_C2 = CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_C3 = CLBLL_L_X4Y103_SLICE_X4Y103_AO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_C4 = CLBLM_L_X8Y103_SLICE_X10Y103_CO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_C5 = CLBLM_R_X7Y102_SLICE_X9Y102_AO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_C6 = CLBLM_R_X5Y102_SLICE_X7Y102_AO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_A6 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_D1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_D2 = CLBLM_R_X5Y103_SLICE_X7Y103_AO6;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_D3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_D4 = CLBLM_R_X7Y103_SLICE_X8Y103_AO5;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_D5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y102_SLICE_X9Y102_D6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C1 = CLBLM_R_X7Y112_SLICE_X9Y112_AO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_A1 = CLBLM_L_X8Y103_SLICE_X10Y103_AO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_A2 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_A3 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_A4 = CLBLM_R_X7Y101_SLICE_X8Y101_BO5;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_A5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_A6 = 1'b1;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_B1 = CLBLM_R_X7Y104_SLICE_X8Y104_BO5;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_B2 = CLBLM_L_X8Y103_SLICE_X10Y103_AO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_B3 = CLBLM_R_X7Y101_SLICE_X8Y101_CO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_B4 = CLBLM_R_X7Y101_SLICE_X8Y101_BO5;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_B5 = CLBLM_R_X7Y102_SLICE_X8Y102_AO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_B6 = CLBLM_R_X7Y100_SLICE_X8Y100_CO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C6 = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_C1 = CLBLM_R_X7Y102_SLICE_X8Y102_AO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_C2 = CLBLM_L_X8Y103_SLICE_X10Y103_AO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_C3 = CLBLM_R_X7Y101_SLICE_X8Y101_CO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_C4 = CLBLM_R_X7Y100_SLICE_X8Y100_CO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_C5 = CLBLM_R_X7Y104_SLICE_X8Y104_BO5;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_C6 = CLBLM_R_X7Y101_SLICE_X8Y101_BO5;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B5 = CLBLM_R_X11Y109_SLICE_X14Y109_AO6;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_B6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_D1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_D2 = CLBLM_R_X7Y100_SLICE_X8Y100_CO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_D3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_D5 = CLBLM_L_X8Y103_SLICE_X10Y103_AO6;
  assign CLBLM_R_X7Y102_SLICE_X8Y102_D6 = CLBLM_R_X7Y101_SLICE_X8Y101_BO5;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D1 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D3 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D4 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C4 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C5 = 1'b1;
  assign CLBLM_R_X11Y110_SLICE_X14Y110_C6 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A3 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A5 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_A6 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B1 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B2 = CLBLM_L_X10Y110_SLICE_X12Y110_BO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B3 = CLBLM_L_X10Y108_SLICE_X13Y108_AO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B4 = CLBLM_L_X10Y107_SLICE_X12Y107_AO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B5 = CLBLM_L_X10Y110_SLICE_X12Y110_AO6;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_B6 = CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C1 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C2 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C3 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C4 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C5 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_C6 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D1 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D2 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D3 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D4 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D5 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X11Y109_D6 = 1'b1;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A4 = CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_A6 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B4 = CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_B6 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C1 = CLBLM_L_X10Y108_SLICE_X12Y108_DO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C5 = CLBLM_L_X8Y109_SLICE_X10Y109_DO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_C6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D2 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y109_SLICE_X10Y109_D6 = CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C1 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C2 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A1 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A4 = CLBLM_R_X7Y103_SLICE_X9Y103_BO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A5 = CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_A6 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_B6 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C1 = CLBLM_L_X8Y104_SLICE_X10Y104_AO6;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_C6 = CLBLM_R_X7Y103_SLICE_X9Y103_BO6;
  assign CLBLM_L_X8Y106_SLICE_X11Y106_D4 = CLBLM_L_X8Y107_SLICE_X11Y107_AO5;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D1 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D2 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D3 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D4 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D5 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X9Y103_D6 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A1 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A3 = CLBLM_R_X7Y103_SLICE_X9Y103_CO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A4 = CLBLM_R_X7Y103_SLICE_X8Y103_BO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_A6 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B3 = CLBLM_R_X7Y105_SLICE_X8Y105_AO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_B6 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D3 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D4 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C1 = CLBLM_R_X7Y101_SLICE_X8Y101_BO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C2 = CLBLM_R_X7Y104_SLICE_X8Y104_CO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_C6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D5 = 1'b1;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D1 = CLBLM_R_X7Y101_SLICE_X8Y101_BO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D2 = CLBLM_R_X7Y104_SLICE_X8Y104_CO6;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y103_SLICE_X8Y103_D6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A1 = CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A2 = CLBLM_L_X10Y110_SLICE_X12Y110_DO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A3 = CLBLM_L_X8Y109_SLICE_X11Y109_AO5;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A4 = CLBLM_R_X7Y110_SLICE_X8Y110_AO5;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A5 = CLBLM_L_X10Y111_SLICE_X12Y111_AO5;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_A6 = CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B1 = CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B2 = CLBLM_L_X10Y110_SLICE_X12Y110_DO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_B6 = CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C1 = CLBLM_L_X8Y109_SLICE_X11Y109_AO5;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C2 = CLBLM_L_X10Y110_SLICE_X12Y110_DO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C3 = CLBLM_L_X10Y111_SLICE_X12Y111_AO5;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C4 = CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C5 = CLBLM_L_X8Y110_SLICE_X11Y110_DO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_C6 = CLBLM_R_X7Y110_SLICE_X8Y110_AO5;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D5 = CLBLM_L_X10Y110_SLICE_X13Y110_CO6;
  assign CLBLM_L_X8Y110_SLICE_X11Y110_D6 = CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A1 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A2 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A3 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A4 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_A6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B1 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B2 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B3 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B4 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_B6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C1 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C2 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C3 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C4 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_C6 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D1 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D2 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D3 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D4 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D5 = 1'b1;
  assign CLBLM_L_X8Y110_SLICE_X10Y110_D6 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A1 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A2 = CLBLM_R_X7Y104_SLICE_X8Y104_DO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A4 = CLBLM_L_X8Y104_SLICE_X11Y104_AO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_A6 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B2 = CLBLM_L_X8Y104_SLICE_X11Y104_BO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B5 = CLBLM_L_X8Y105_SLICE_X10Y105_DO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_B6 = CLBLM_R_X7Y104_SLICE_X9Y104_CO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C1 = CLBLM_R_X7Y104_SLICE_X9Y104_AO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C2 = CLBLM_L_X10Y104_SLICE_X12Y104_CO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C3 = CLBLM_L_X10Y104_SLICE_X12Y104_BO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C4 = CLBLM_L_X8Y105_SLICE_X10Y105_AO5;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C5 = CLBLM_R_X7Y104_SLICE_X8Y104_AO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_C6 = CLBLM_L_X10Y104_SLICE_X12Y104_AO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D2 = CLBLM_L_X8Y104_SLICE_X11Y104_BO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D4 = CLBLM_L_X8Y104_SLICE_X10Y104_BO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D5 = CLBLM_L_X8Y105_SLICE_X10Y105_DO6;
  assign CLBLM_R_X7Y104_SLICE_X9Y104_D6 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A2 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A4 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A5 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_A6 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B1 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B2 = 1'b1;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_B6 = 1'b1;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_D = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_D = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C1 = CLBLM_L_X8Y102_SLICE_X10Y102_BO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C3 = CLBLM_L_X10Y103_SLICE_X12Y103_AO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_C6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D1 = CLBLM_L_X8Y102_SLICE_X10Y102_BO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D3 = CLBLM_L_X10Y103_SLICE_X12Y103_AO6;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y104_SLICE_X8Y104_D6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A1 = CLBLM_L_X8Y112_SLICE_X11Y112_DO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A2 = CLBLM_L_X10Y110_SLICE_X13Y110_BO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A3 = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A4 = CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A5 = CLBLM_L_X10Y111_SLICE_X12Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_A6 = CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B1 = CLBLL_L_X4Y111_SLICE_X5Y111_AO5;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B2 = CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B3 = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B4 = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B5 = CLBLM_R_X11Y110_SLICE_X14Y110_AO5;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_B6 = CLBLM_L_X8Y112_SLICE_X11Y112_AO5;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C2 = CLBLM_L_X10Y110_SLICE_X12Y110_CO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C5 = CLBLM_L_X8Y111_SLICE_X11Y111_DO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_C6 = CLBLM_L_X10Y111_SLICE_X12Y111_CO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D2 = CLBLM_L_X10Y111_SLICE_X12Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D4 = CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y111_SLICE_X11Y111_D6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A2 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A4 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_A6 = 1'b1;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B1 = CLBLM_L_X8Y112_SLICE_X11Y112_AO5;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B2 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B3 = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B4 = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B5 = CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_B6 = CLBLM_L_X8Y111_SLICE_X10Y111_AO5;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C1 = CLBLM_L_X8Y111_SLICE_X10Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C2 = CLBLM_L_X8Y112_SLICE_X11Y112_AO5;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C3 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C4 = CLBLM_L_X8Y111_SLICE_X10Y111_AO5;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C5 = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_C6 = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D2 = CLBLM_L_X8Y112_SLICE_X10Y112_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D4 = CLBLM_L_X10Y111_SLICE_X12Y111_BO6;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y111_SLICE_X10Y111_D6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_A1 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_A2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_A3 = CLBLL_L_X2Y103_SLICE_X1Y103_AO6;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_A4 = CLBLL_L_X2Y103_SLICE_X0Y103_BO6;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_A5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_A6 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_B1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_B2 = CLBLL_L_X2Y103_SLICE_X1Y103_DO6;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_B4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_B5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_B6 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B3 = CLBLM_R_X3Y111_SLICE_X2Y111_DO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B4 = CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_C1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_C2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_C3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_C4 = CLBLL_L_X2Y103_SLICE_X0Y103_AO5;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_C5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_C6 = CLBLL_L_X2Y104_SLICE_X0Y104_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B5 = CLBLL_L_X4Y112_SLICE_X4Y112_AO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_B6 = CLBLL_L_X4Y112_SLICE_X4Y112_AO5;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_D1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_D2 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_D3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_D4 = CLBLL_L_X2Y103_SLICE_X0Y103_AO5;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_D5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_D6 = CLBLL_L_X2Y104_SLICE_X0Y104_AO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A1 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A2 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A3 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A4 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A5 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_A6 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B1 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B2 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B3 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B4 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B5 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_A1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_A2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_A3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_A4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_A5 = CLBLL_L_X2Y103_SLICE_X1Y103_CO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_A6 = CLBLL_L_X4Y102_SLICE_X4Y102_BO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C2 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C3 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_B6 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C5 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C1 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_B1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_B2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_B3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_B4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_B5 = CLBLL_L_X2Y103_SLICE_X1Y103_CO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_B6 = CLBLL_L_X4Y102_SLICE_X4Y102_BO6;
  assign CLBLL_L_X4Y112_SLICE_X4Y112_C6 = CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D1 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D2 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D3 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D4 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D5 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_D6 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_C1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_C2 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_C3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_C4 = CLBLM_R_X3Y102_SLICE_X2Y102_AO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_C5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_A6 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_D1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_D2 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_D3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B1 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_D4 = CLBLM_R_X3Y102_SLICE_X2Y102_AO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_D5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B4 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_D6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B6 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B2 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B3 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_B5 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C1 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C2 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C3 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C4 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C5 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_C6 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D1 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D2 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D3 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D4 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D5 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X8Y105_D6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A1 = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A2 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A5 = CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_A6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B1 = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B2 = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_B6 = CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_C6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D1 = CLBLM_L_X8Y112_SLICE_X11Y112_CO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D2 = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D3 = CLBLM_R_X11Y110_SLICE_X14Y110_AO5;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D4 = CLBLM_L_X8Y112_SLICE_X11Y112_AO5;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D5 = CLBLL_L_X4Y111_SLICE_X5Y111_AO5;
  assign CLBLM_L_X8Y112_SLICE_X11Y112_D6 = CLBLM_L_X10Y109_SLICE_X12Y109_BO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A2 = CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A3 = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_A6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B2 = CLBLM_L_X8Y112_SLICE_X11Y112_BO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B3 = CLBLM_L_X8Y111_SLICE_X10Y111_CO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_B6 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C1 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C2 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C3 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C4 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C5 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_C6 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A1 = CLBLL_L_X2Y103_SLICE_X1Y103_DO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D6 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D1 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B1 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B2 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B3 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B4 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B5 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B6 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C1 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C2 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C3 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C4 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C5 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C6 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_D1 = CLBLL_L_X2Y113_SLICE_X0Y113_AO5;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D1 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D2 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D3 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D4 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D5 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D6 = 1'b1;
  assign LIOI3_X0Y117_OLOGIC_X0Y118_T1 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A1 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A2 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_A6 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A1 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A2 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A3 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B5 = CLBLM_L_X8Y106_SLICE_X10Y106_BO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B6 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A4 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A5 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A6 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B2 = CLBLM_L_X8Y105_SLICE_X10Y105_CO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C6 = CLBLM_L_X8Y106_SLICE_X10Y106_AO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B1 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B2 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B3 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B4 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B5 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B6 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C1 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C2 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C3 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D2 = CLBLM_R_X7Y104_SLICE_X9Y104_CO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D3 = CLBLM_R_X7Y107_SLICE_X9Y107_AO5;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D4 = CLBLM_R_X7Y106_SLICE_X9Y106_AO5;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D5 = CLBLM_L_X8Y106_SLICE_X11Y106_DO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D6 = CLBLM_L_X8Y106_SLICE_X10Y106_DO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C4 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C5 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C6 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D1 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D2 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A1 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A2 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A3 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A4 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A5 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_A6 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D3 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D4 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D5 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D6 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B2 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B3 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B4 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B5 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B6 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_B1 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C1 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C2 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C3 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C4 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C5 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_C6 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D1 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D2 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D3 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D4 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D5 = 1'b1;
  assign CLBLM_R_X7Y106_SLICE_X8Y106_D6 = 1'b1;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_D = LIOB33_X0Y117_IOB_X0Y117_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y102_D = RIOB33_X105Y101_IOB_X1Y102_I;
  assign RIOI3_X105Y101_ILOGIC_X1Y101_D = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A1 = CLBLL_L_X2Y103_SLICE_X1Y103_DO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B5 = CLBLL_L_X2Y105_SLICE_X0Y105_AO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B6 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C1 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C2 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C3 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C4 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C5 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C6 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D1 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D2 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D3 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D4 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D5 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D6 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A1 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A4 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_A6 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A1 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A2 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A3 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A4 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A5 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A6 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B1 = CLBLM_L_X8Y102_SLICE_X10Y102_CO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B2 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B1 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B2 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C2 = CLBLM_R_X11Y107_SLICE_X14Y107_BO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B3 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B4 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B5 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B6 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C1 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C2 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C3 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C4 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C5 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C6 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D1 = CLBLM_R_X7Y107_SLICE_X9Y107_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D2 = CLBLM_L_X8Y107_SLICE_X11Y107_BO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D3 = CLBLM_L_X8Y108_SLICE_X10Y108_CO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D1 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D2 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D3 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D4 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D5 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D6 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D4 = CLBLM_L_X8Y107_SLICE_X11Y107_CO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A2 = CLBLM_L_X8Y107_SLICE_X11Y107_BO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A3 = CLBLM_R_X7Y107_SLICE_X9Y107_CO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_A6 = CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B1 = CLBLM_L_X8Y107_SLICE_X11Y107_DO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B3 = CLBLM_R_X7Y107_SLICE_X9Y107_CO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_B6 = CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C2 = CLBLM_R_X7Y107_SLICE_X9Y107_CO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C5 = CLBLM_L_X8Y107_SLICE_X11Y107_BO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_C6 = CLBLM_L_X8Y108_SLICE_X10Y108_BO6;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D1 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D2 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D3 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D4 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D5 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X8Y107_D6 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A1 = CLBLL_L_X2Y103_SLICE_X0Y103_DO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A2 = CLBLL_L_X2Y105_SLICE_X0Y105_BO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A3 = CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A4 = CLBLM_R_X3Y103_SLICE_X2Y103_CO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A5 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A6 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B2 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B6 = CLBLL_L_X2Y105_SLICE_X0Y105_AO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C1 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C3 = CLBLL_L_X2Y103_SLICE_X0Y103_DO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C4 = CLBLM_R_X3Y103_SLICE_X2Y103_CO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C5 = CLBLL_L_X2Y106_SLICE_X0Y106_DO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C6 = CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D3 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D4 = CLBLL_L_X2Y105_SLICE_X0Y105_AO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D6 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A1 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A2 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A3 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A5 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A6 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A4 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A5 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A6 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B5 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B6 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B1 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B2 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B3 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B4 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C3 = CLBLM_L_X8Y108_SLICE_X10Y108_CO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C4 = CLBLM_L_X8Y107_SLICE_X11Y107_BO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C5 = CLBLM_R_X7Y108_SLICE_X9Y108_BO5;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C1 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C2 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C3 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C4 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C5 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C6 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X11Y107_D3 = CLBLM_L_X10Y107_SLICE_X12Y107_DO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C6 = CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D1 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D2 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D3 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D4 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D5 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D6 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D1 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D2 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D3 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D4 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D5 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A1 = CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A2 = CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_A6 = CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B1 = CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B2 = CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_B6 = CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C2 = CLBLM_L_X8Y109_SLICE_X10Y109_CO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C3 = CLBLM_L_X8Y108_SLICE_X10Y108_DO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C5 = CLBLM_R_X7Y109_SLICE_X8Y109_DO6;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_C6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D1 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D2 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D3 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D4 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D5 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X8Y108_D6 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = CLBLL_L_X2Y112_SLICE_X0Y112_BO5;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign CLBLM_L_X8Y107_SLICE_X10Y107_B5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A1 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A3 = 1'b1;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_A6 = 1'b1;
  assign RIOI3_X105Y103_ILOGIC_X1Y104_D = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B2 = CLBLM_L_X8Y109_SLICE_X10Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B4 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_B6 = CLBLM_L_X8Y109_SLICE_X11Y109_BO6;
  assign RIOI3_X105Y103_ILOGIC_X1Y103_D = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C1 = CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C2 = CLBLM_L_X8Y109_SLICE_X11Y109_BO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C3 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C4 = CLBLM_R_X7Y109_SLICE_X9Y109_AO5;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C5 = CLBLM_R_X7Y108_SLICE_X9Y108_AO5;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_C6 = CLBLM_L_X8Y109_SLICE_X10Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D1 = CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D2 = CLBLM_L_X8Y109_SLICE_X11Y109_BO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D3 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D4 = CLBLM_R_X7Y109_SLICE_X9Y109_AO5;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D5 = CLBLM_R_X7Y108_SLICE_X9Y108_AO5;
  assign CLBLM_R_X7Y109_SLICE_X9Y109_D6 = CLBLM_L_X8Y109_SLICE_X10Y109_AO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A1 = CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A2 = CLBLM_R_X7Y109_SLICE_X9Y109_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A4 = CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_A6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B1 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_B6 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C1 = CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C2 = CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C3 = CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C4 = CLBLM_R_X5Y110_SLICE_X7Y110_DO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C5 = CLBLM_R_X3Y110_SLICE_X3Y110_AO5;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_C6 = CLBLM_R_X7Y108_SLICE_X9Y108_BO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D3 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D5 = CLBLM_R_X7Y110_SLICE_X8Y110_CO6;
  assign CLBLM_R_X7Y109_SLICE_X8Y109_D6 = CLBLM_L_X8Y111_SLICE_X11Y111_CO6;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C1 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C4 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A4 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A5 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_A6 = 1'b1;
  assign CLBLL_L_X4Y113_SLICE_X4Y113_C6 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B1 = CLBLM_L_X8Y110_SLICE_X11Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B2 = CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B3 = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B4 = CLBLM_L_X10Y110_SLICE_X12Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B5 = CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_B6 = CLBLM_R_X7Y110_SLICE_X9Y110_AO5;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_A1 = CLBLM_R_X5Y102_SLICE_X7Y102_CO6;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_A2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_A3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C4 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C5 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C6 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_A4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_A5 = CLBLM_R_X7Y102_SLICE_X9Y102_DO6;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_A6 = CLBLM_R_X7Y101_SLICE_X8Y101_AO5;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C1 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_C2 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_B1 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_B2 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_B3 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_B4 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_B5 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_B6 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D5 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D6 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D1 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X9Y110_D2 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_C1 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_C2 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_C3 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_C4 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_C5 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_C6 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A1 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A5 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_A6 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_D1 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_D2 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_D3 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_D4 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_D5 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X7Y100_D6 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B6 = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B3 = CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_B4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C2 = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C3 = CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_C6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_A1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_A2 = CLBLM_R_X7Y100_SLICE_X8Y100_AO6;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_A3 = CLBLM_R_X5Y100_SLICE_X7Y100_AO6;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_A4 = CLBLM_R_X7Y100_SLICE_X8Y100_BO6;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_A5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_A6 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_B1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_B2 = CLBLM_R_X7Y100_SLICE_X8Y100_AO6;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_B3 = CLBLM_R_X5Y100_SLICE_X7Y100_AO6;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_B4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_B5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_B6 = CLBLM_R_X7Y100_SLICE_X8Y100_BO6;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D3 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_C1 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_C2 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_C3 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_C4 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_C5 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_C6 = 1'b1;
  assign CLBLM_R_X7Y110_SLICE_X8Y110_D6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_D1 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_D2 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_D3 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_D4 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_D5 = 1'b1;
  assign CLBLM_R_X5Y100_SLICE_X6Y100_D6 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = CLBLL_L_X2Y112_SLICE_X1Y112_BO6;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_A6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B1 = CLBLM_R_X7Y112_SLICE_X9Y112_BO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B2 = CLBLM_R_X7Y111_SLICE_X8Y111_BO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B5 = CLBLM_R_X7Y111_SLICE_X9Y111_AO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_B6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_A1 = CLBLM_R_X5Y101_SLICE_X7Y101_DO6;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_A2 = CLBLM_R_X5Y101_SLICE_X6Y101_BO6;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_A3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C4 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C5 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C6 = 1'b1;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_A4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_A6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C1 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_C2 = 1'b1;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_B2 = CLBLM_R_X7Y102_SLICE_X8Y102_AO5;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_B3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_B4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_B5 = CLBLM_R_X7Y101_SLICE_X8Y101_CO5;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_B6 = CLBLM_R_X5Y100_SLICE_X6Y100_BO6;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D5 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D6 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D1 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X9Y111_D2 = 1'b1;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_C1 = CLBLM_R_X7Y101_SLICE_X8Y101_CO5;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_C2 = CLBLM_R_X7Y102_SLICE_X8Y102_AO5;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_C3 = CLBLM_R_X5Y100_SLICE_X6Y100_BO6;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_C5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_C6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A1 = CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A3 = 1'b1;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A5 = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_A6 = 1'b1;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_D1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_D2 = CLBLM_R_X5Y102_SLICE_X7Y102_CO6;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_D3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_D4 = CLBLM_R_X7Y101_SLICE_X8Y101_AO5;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_D5 = CLBLM_R_X7Y102_SLICE_X9Y102_DO6;
  assign CLBLM_R_X5Y101_SLICE_X7Y101_D6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B6 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_A1 = CLBLM_R_X5Y101_SLICE_X6Y101_DO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C4 = CLBLM_L_X8Y110_SLICE_X11Y110_BO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_C6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_A2 = CLBLL_L_X4Y102_SLICE_X5Y102_CO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_A3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_A5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_A6 = 1'b1;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_B1 = CLBLM_R_X5Y102_SLICE_X7Y102_AO5;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_B2 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_B3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_B4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_B5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_B6 = CLBLM_R_X5Y102_SLICE_X6Y102_BO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D1 = CLBLM_R_X7Y111_SLICE_X8Y111_CO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D3 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_C1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_C2 = CLBLL_L_X4Y102_SLICE_X5Y102_CO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_C3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_C4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_C5 = CLBLM_R_X5Y102_SLICE_X7Y102_AO5;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_C6 = CLBLM_R_X5Y102_SLICE_X7Y102_BO6;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X7Y111_SLICE_X8Y111_D6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_D1 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_D2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_D3 = CLBLM_R_X5Y102_SLICE_X6Y102_BO6;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_D4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_D5 = CLBLM_R_X5Y102_SLICE_X7Y102_AO5;
  assign CLBLM_R_X5Y101_SLICE_X6Y101_D6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y106_D = RIOB33_X105Y105_IOB_X1Y106_I;
  assign RIOI3_X105Y105_ILOGIC_X1Y105_D = RIOB33_X105Y105_IOB_X1Y105_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D = LIOB33_X0Y107_IOB_X0Y107_I;
  assign RIOI3_TBYTETERM_X105Y113_ILOGIC_X1Y113_D = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C6 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A1 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_A5 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_B1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D1 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C2 = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C3 = CLBLM_L_X8Y112_SLICE_X11Y112_DO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C4 = CLBLM_R_X7Y112_SLICE_X9Y112_AO5;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_C5 = CLBLM_L_X8Y111_SLICE_X10Y111_BO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D6 = 1'b1;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_A2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_A4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_A5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_A6 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D2 = 1'b1;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_B1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_B2 = CLBLM_R_X5Y102_SLICE_X6Y102_BO6;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D5 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X9Y112_D6 = 1'b1;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_B3 = CLBLM_R_X5Y103_SLICE_X7Y103_AO6;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_B4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_B6 = 1'b1;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_C1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_C2 = CLBLL_L_X4Y102_SLICE_X5Y102_DO6;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_C3 = CLBLM_R_X7Y103_SLICE_X8Y103_AO5;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_C4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_C5 = CLBLM_R_X5Y102_SLICE_X7Y102_BO5;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_C6 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A2 = CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_A5 = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_D1 = CLBLM_R_X5Y103_SLICE_X7Y103_AO6;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_D2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_D3 = CLBLM_R_X7Y103_SLICE_X8Y103_AO5;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_D4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_D5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B5 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B6 = 1'b1;
  assign CLBLM_R_X5Y102_SLICE_X7Y102_D6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B1 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B2 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B3 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_B4 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C3 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C4 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C5 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_C6 = 1'b1;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_A1 = CLBLM_R_X5Y102_SLICE_X6Y102_DO6;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_A2 = CLBLM_R_X7Y102_SLICE_X8Y102_CO6;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_A3 = CLBLM_R_X7Y104_SLICE_X8Y104_AO5;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_A4 = CLBLM_R_X7Y103_SLICE_X8Y103_DO6;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_A5 = CLBLM_R_X5Y100_SLICE_X6Y100_BO6;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_A6 = CLBLM_R_X7Y102_SLICE_X8Y102_BO6;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_B1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_B2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_B3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_B4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D2 = 1'b1;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_B5 = CLBLM_R_X5Y102_SLICE_X6Y102_CO6;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_B6 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D6 = 1'b1;
  assign CLBLM_R_X7Y112_SLICE_X8Y112_D1 = 1'b1;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_C1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_C2 = CLBLM_R_X7Y105_SLICE_X8Y105_AO6;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_C3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_C4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_C5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_C6 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_D1 = 1'b1;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_D2 = 1'b1;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_D3 = 1'b1;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_D5 = 1'b1;
  assign CLBLM_R_X5Y102_SLICE_X6Y102_D6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A4 = CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A5 = CLBLL_L_X2Y111_SLICE_X0Y111_CO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_A6 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_B6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_C6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D1 = CLBLL_L_X2Y111_SLICE_X0Y111_AO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D3 = CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y111_SLICE_X0Y111_D6 = CLBLL_L_X2Y112_SLICE_X0Y112_AO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A3 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A5 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_A6 = 1'b1;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B1 = CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B3 = CLBLL_L_X2Y111_SLICE_X0Y111_CO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B5 = CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_B6 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C1 = CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C2 = CLBLL_L_X2Y111_SLICE_X0Y111_AO5;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C3 = CLBLM_R_X3Y111_SLICE_X2Y111_AO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_C6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_D1 = CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D1 = CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D2 = CLBLL_L_X2Y111_SLICE_X0Y111_CO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D3 = CLBLL_L_X2Y112_SLICE_X1Y112_AO5;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D4 = CLBLL_L_X2Y111_SLICE_X1Y111_AO5;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D5 = CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  assign CLBLL_L_X2Y111_SLICE_X1Y111_D6 = CLBLM_R_X3Y111_SLICE_X3Y111_AO5;
  assign LIOI3_X0Y125_OLOGIC_X0Y126_T1 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_A1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_A2 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_A3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_A4 = CLBLM_R_X7Y105_SLICE_X8Y105_AO6;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_A5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_A6 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_D1 = CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_B1 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_B2 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_B3 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_B4 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_B5 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_B6 = 1'b1;
  assign LIOI3_X0Y125_OLOGIC_X0Y125_T1 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_C1 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_C2 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_C3 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_C4 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_C5 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_C6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_D1 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_D2 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_D3 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_D4 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_D5 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_A1 = CLBLM_R_X7Y104_SLICE_X9Y104_AO5;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_A2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_A3 = CLBLM_R_X7Y103_SLICE_X8Y103_CO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_A4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_A5 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = CLBLM_R_X3Y109_SLICE_X2Y109_BO5;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_B1 = CLBLM_R_X7Y104_SLICE_X9Y104_AO5;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_B2 = CLBLM_R_X7Y103_SLICE_X8Y103_DO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_B3 = CLBLM_R_X7Y103_SLICE_X8Y103_CO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_B4 = CLBLM_R_X7Y102_SLICE_X8Y102_BO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_B5 = CLBLM_R_X5Y103_SLICE_X6Y103_AO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_B6 = CLBLM_R_X7Y104_SLICE_X8Y104_AO5;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_C1 = CLBLM_R_X5Y104_SLICE_X6Y104_AO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_C2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_C3 = CLBLM_R_X5Y104_SLICE_X6Y104_DO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_C4 = CLBLM_R_X5Y105_SLICE_X6Y105_DO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_C5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_C6 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_D1 = CLBLM_R_X5Y104_SLICE_X6Y104_AO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_D2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_D3 = CLBLM_R_X5Y104_SLICE_X6Y104_DO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_D4 = CLBLM_R_X5Y105_SLICE_X6Y105_DO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_D5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_D6 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A1 = CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A4 = CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_A6 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B3 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B5 = CLBLL_L_X2Y112_SLICE_X0Y112_CO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_B6 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C2 = CLBLL_L_X2Y111_SLICE_X0Y111_CO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C5 = CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_C6 = CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  assign RIOI3_X105Y109_ILOGIC_X1Y110_D = RIOB33_X105Y109_IOB_X1Y110_I;
  assign RIOI3_X105Y109_ILOGIC_X1Y109_D = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D2 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y112_SLICE_X0Y112_D6 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A1 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A2 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_A6 = 1'b1;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B4 = CLBLL_L_X2Y111_SLICE_X1Y111_CO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_B6 = CLBLL_L_X2Y112_SLICE_X1Y112_CO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C2 = CLBLL_L_X2Y111_SLICE_X1Y111_BO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C5 = CLBLL_L_X2Y112_SLICE_X1Y112_DO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_C6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D1 = CLBLL_L_X2Y112_SLICE_X1Y112_AO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D2 = CLBLL_L_X2Y111_SLICE_X0Y111_CO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D3 = CLBLL_L_X2Y112_SLICE_X0Y112_DO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D4 = CLBLL_L_X2Y112_SLICE_X1Y112_AO5;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D5 = CLBLL_L_X2Y112_SLICE_X0Y112_BO6;
  assign CLBLL_L_X2Y112_SLICE_X1Y112_D6 = CLBLL_L_X2Y111_SLICE_X0Y111_BO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A2 = CLBLM_R_X7Y104_SLICE_X9Y104_BO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A3 = CLBLM_R_X7Y104_SLICE_X9Y104_AO5;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A4 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A5 = CLBLM_R_X7Y103_SLICE_X8Y103_CO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A6 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B1 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B2 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B3 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B4 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B5 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B6 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C1 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C2 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C3 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C4 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C5 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C6 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D1 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D2 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D3 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D4 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D5 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D6 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A1 = CLBLM_R_X5Y104_SLICE_X7Y104_AO5;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A2 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A3 = CLBLM_R_X5Y104_SLICE_X7Y104_AO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A4 = CLBLM_R_X7Y104_SLICE_X9Y104_BO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A6 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B2 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B3 = CLBLM_R_X5Y105_SLICE_X6Y105_DO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B5 = CLBLM_R_X5Y104_SLICE_X6Y104_AO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B6 = CLBLM_R_X5Y104_SLICE_X6Y104_CO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C2 = CLBLM_R_X5Y104_SLICE_X7Y104_AO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C4 = CLBLM_R_X7Y104_SLICE_X9Y104_BO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C6 = CLBLM_R_X5Y103_SLICE_X6Y103_BO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D1 = CLBLL_L_X4Y103_SLICE_X5Y103_AO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D2 = CLBLM_R_X5Y104_SLICE_X7Y104_AO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D3 = CLBLL_L_X4Y104_SLICE_X5Y104_AO5;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D4 = CLBLM_R_X7Y104_SLICE_X9Y104_BO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D5 = CLBLM_R_X5Y105_SLICE_X6Y105_AO5;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D6 = CLBLM_R_X5Y103_SLICE_X6Y103_BO6;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A2 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A4 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_A6 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_B6 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_C6 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X0Y113_D6 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_A6 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_B6 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_C6 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D1 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D2 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D3 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D4 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D5 = 1'b1;
  assign CLBLL_L_X2Y113_SLICE_X1Y113_D6 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A2 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A5 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A6 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B1 = CLBLM_R_X5Y105_SLICE_X7Y105_DO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B2 = CLBLM_R_X5Y101_SLICE_X7Y101_BO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B4 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B6 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C3 = CLBLM_R_X7Y102_SLICE_X8Y102_DO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C4 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C5 = CLBLM_R_X7Y103_SLICE_X8Y103_DO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D2 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D3 = CLBLM_R_X7Y102_SLICE_X8Y102_DO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D5 = CLBLM_R_X7Y103_SLICE_X8Y103_DO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A2 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A3 = CLBLM_R_X5Y104_SLICE_X7Y104_AO5;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A4 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A6 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B2 = CLBLM_R_X5Y105_SLICE_X6Y105_DO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B3 = CLBLM_R_X5Y104_SLICE_X7Y104_AO5;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B4 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B6 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C1 = CLBLM_R_X7Y104_SLICE_X9Y104_DO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C2 = CLBLM_R_X7Y106_SLICE_X9Y106_CO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C5 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D1 = CLBLM_R_X7Y104_SLICE_X9Y104_DO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D2 = CLBLM_R_X7Y106_SLICE_X9Y106_CO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D3 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_D1 = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign LIOI3_X0Y127_OLOGIC_X0Y128_T1 = 1'b1;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_D1 = CLBLM_R_X3Y111_SLICE_X3Y111_BO5;
  assign LIOI3_X0Y127_OLOGIC_X0Y127_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_D1 = CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y132_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_D1 = CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  assign LIOI3_TBYTESRC_X0Y131_OLOGIC_X0Y131_T1 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A1 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A5 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A6 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B4 = CLBLM_R_X7Y107_SLICE_X8Y107_CO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B6 = CLBLM_L_X8Y106_SLICE_X10Y106_CO6;
  assign RIOI3_X105Y111_ILOGIC_X1Y112_D = RIOB33_X105Y111_IOB_X1Y112_I;
  assign RIOI3_X105Y111_ILOGIC_X1Y111_D = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C3 = CLBLM_R_X7Y107_SLICE_X8Y107_CO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C4 = CLBLM_L_X8Y106_SLICE_X10Y106_CO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D1 = CLBLM_R_X5Y106_SLICE_X7Y106_AO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D2 = CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D3 = CLBLM_R_X5Y106_SLICE_X7Y106_AO5;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D4 = CLBLM_R_X5Y106_SLICE_X7Y106_CO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D5 = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D6 = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A2 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A5 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A6 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B3 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B4 = CLBLM_L_X8Y107_SLICE_X10Y107_CO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B6 = CLBLM_R_X7Y106_SLICE_X9Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C1 = CLBLM_R_X7Y106_SLICE_X9Y106_DO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C2 = CLBLM_R_X5Y105_SLICE_X7Y105_AO5;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C3 = CLBLM_L_X8Y107_SLICE_X10Y107_CO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C4 = CLBLM_R_X5Y106_SLICE_X6Y106_AO5;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C5 = CLBLM_R_X7Y107_SLICE_X9Y107_AO5;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C6 = CLBLM_R_X7Y106_SLICE_X9Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D2 = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D3 = CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D4 = CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D6 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A1 = CLBLM_R_X5Y105_SLICE_X7Y105_AO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A2 = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A3 = CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A4 = CLBLM_R_X7Y107_SLICE_X9Y107_DO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A5 = CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A6 = CLBLM_R_X5Y106_SLICE_X7Y106_AO5;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B2 = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B5 = CLBLM_R_X7Y107_SLICE_X8Y107_BO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C1 = CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C2 = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C3 = CLBLM_L_X8Y107_SLICE_X10Y107_DO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C4 = CLBLM_R_X7Y107_SLICE_X8Y107_CO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C5 = CLBLM_R_X5Y105_SLICE_X7Y105_AO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C6 = CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D1 = CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D2 = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D3 = CLBLM_R_X7Y107_SLICE_X9Y107_DO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D4 = CLBLM_R_X5Y106_SLICE_X7Y106_AO5;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D5 = CLBLM_R_X5Y105_SLICE_X7Y105_AO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D6 = CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A3 = CLBLM_R_X7Y107_SLICE_X8Y107_BO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A6 = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B2 = CLBLM_R_X7Y106_SLICE_X9Y106_BO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B6 = CLBLM_L_X8Y107_SLICE_X10Y107_CO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C3 = CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C4 = CLBLL_L_X4Y106_SLICE_X4Y106_AO5;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C6 = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D2 = CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D3 = CLBLM_R_X5Y107_SLICE_X7Y107_DO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D4 = CLBLM_R_X5Y106_SLICE_X7Y106_AO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D6 = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_D1 = CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y130_T1 = 1'b1;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_D1 = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign LIOI3_X0Y129_OLOGIC_X0Y129_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_D1 = CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y144_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_D1 = CLBLM_R_X3Y104_SLICE_X2Y104_DO6;
  assign LIOI3_TBYTESRC_X0Y143_OLOGIC_X0Y143_T1 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A1 = CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A2 = CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A3 = CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A4 = CLBLM_R_X7Y108_SLICE_X8Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A5 = CLBLM_R_X7Y107_SLICE_X8Y107_AO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_A6 = CLBLL_L_X4Y108_SLICE_X4Y108_AO5;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B1 = CLBLM_R_X5Y109_SLICE_X7Y109_BO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B2 = CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B3 = CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_B6 = CLBLM_R_X7Y106_SLICE_X9Y106_BO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C1 = CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C2 = CLBLM_R_X7Y108_SLICE_X8Y108_BO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C3 = CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C4 = CLBLL_L_X4Y108_SLICE_X4Y108_AO5;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C5 = CLBLM_R_X7Y108_SLICE_X9Y108_CO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_C6 = CLBLM_R_X3Y109_SLICE_X3Y109_AO5;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D1 = CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D2 = CLBLM_L_X10Y108_SLICE_X13Y108_BO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D3 = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D4 = CLBLM_R_X5Y109_SLICE_X7Y109_DO6;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D5 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X7Y108_D6 = CLBLM_L_X8Y109_SLICE_X10Y109_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A1 = CLBLM_R_X5Y109_SLICE_X6Y109_DO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A3 = CLBLM_R_X7Y108_SLICE_X8Y108_CO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_A6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B1 = CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B3 = CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B5 = CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_B6 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_B6 = 1'b1;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C1 = CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C2 = CLBLM_R_X5Y108_SLICE_X7Y108_CO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C5 = CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_C6 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D1 = CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D2 = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D3 = CLBLM_R_X5Y108_SLICE_X7Y108_DO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D4 = CLBLM_R_X7Y106_SLICE_X9Y106_BO6;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D5 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X5Y108_SLICE_X6Y108_D6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_C4 = 1'b1;
  assign CLBLM_R_X11Y103_SLICE_X15Y103_C6 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C4 = 1'b1;
  assign CLBLM_R_X7Y105_SLICE_X9Y105_C6 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A3 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A4 = CLBLM_R_X3Y109_SLICE_X2Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_A6 = 1'b1;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B1 = CLBLL_L_X2Y111_SLICE_X0Y111_DO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B2 = CLBLM_R_X3Y109_SLICE_X2Y109_AO5;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B3 = CLBLM_R_X11Y106_SLICE_X15Y106_DO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B4 = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B5 = CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_B6 = CLBLM_R_X5Y109_SLICE_X7Y109_CO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C4 = CLBLM_R_X7Y103_SLICE_X9Y103_AO5;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_C6 = CLBLM_R_X3Y109_SLICE_X2Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D1 = CLBLM_R_X5Y109_SLICE_X7Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D2 = CLBLM_R_X7Y103_SLICE_X9Y103_AO5;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D3 = CLBLL_L_X2Y111_SLICE_X0Y111_DO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D5 = CLBLM_R_X11Y106_SLICE_X15Y106_DO6;
  assign CLBLM_R_X5Y109_SLICE_X7Y109_D6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A1 = CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A2 = CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A4 = CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_A6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B1 = CLBLM_R_X5Y108_SLICE_X7Y108_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B3 = CLBLM_R_X5Y108_SLICE_X6Y108_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_B6 = CLBLM_R_X5Y109_SLICE_X6Y109_CO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C1 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C3 = CLBLM_R_X5Y110_SLICE_X7Y110_BO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C4 = CLBLM_R_X7Y109_SLICE_X8Y109_AO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_C6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D2 = CLBLM_R_X7Y110_SLICE_X8Y110_DO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D4 = CLBLM_R_X7Y109_SLICE_X8Y109_BO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D5 = CLBLM_R_X7Y109_SLICE_X9Y109_DO6;
  assign CLBLM_R_X5Y109_SLICE_X6Y109_D6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A1 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A2 = CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A5 = CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_A6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_D1 = 1'b0;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B1 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B4 = CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_B6 = CLBLM_R_X5Y110_SLICE_X7Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C1 = CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C2 = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C3 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C4 = CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C5 = CLBLL_L_X4Y103_SLICE_X5Y103_BO5;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_C6 = CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y134_T1 = 1'b1;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_D1 = CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D1 = CLBLM_R_X7Y110_SLICE_X8Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D2 = CLBLM_R_X7Y110_SLICE_X9Y110_BO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D3 = CLBLM_R_X5Y111_SLICE_X7Y111_DO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D4 = CLBLL_L_X4Y103_SLICE_X5Y103_BO5;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D5 = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X5Y110_SLICE_X7Y110_D6 = CLBLM_R_X7Y109_SLICE_X9Y109_AO6;
  assign LIOI3_X0Y133_OLOGIC_X0Y133_T1 = 1'b1;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A1 = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A2 = CLBLM_R_X5Y112_SLICE_X6Y112_AO5;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A3 = CLBLM_R_X7Y110_SLICE_X8Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A4 = CLBLM_L_X8Y109_SLICE_X11Y109_AO5;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A5 = CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_A6 = CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B1 = CLBLM_R_X5Y112_SLICE_X6Y112_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B2 = CLBLM_L_X8Y110_SLICE_X11Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B3 = CLBLM_R_X7Y110_SLICE_X9Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B4 = CLBLM_R_X3Y112_SLICE_X3Y112_AO5;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B5 = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_B6 = CLBLM_R_X5Y110_SLICE_X6Y110_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C1 = CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C2 = CLBLM_L_X8Y109_SLICE_X11Y109_AO5;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C3 = CLBLM_R_X5Y112_SLICE_X6Y112_AO5;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C4 = CLBLM_R_X7Y110_SLICE_X8Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C5 = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_C6 = CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D2 = CLBLM_R_X5Y110_SLICE_X7Y110_AO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D4 = CLBLM_R_X7Y111_SLICE_X8Y111_DO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D5 = CLBLM_R_X5Y111_SLICE_X6Y111_CO6;
  assign CLBLM_R_X5Y110_SLICE_X6Y110_D6 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A1 = CLBLM_R_X5Y111_SLICE_X7Y111_BO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A4 = CLBLM_R_X5Y112_SLICE_X7Y112_BO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_A6 = CLBLM_R_X7Y111_SLICE_X8Y111_AO5;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B1 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B4 = CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B5 = CLBLM_R_X7Y112_SLICE_X8Y112_AO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_B6 = CLBLM_L_X8Y111_SLICE_X11Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C1 = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C4 = CLBLM_R_X7Y111_SLICE_X8Y111_AO5;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_C6 = CLBLM_R_X5Y112_SLICE_X7Y112_BO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D1 = CLBLM_R_X5Y110_SLICE_X6Y110_AO6;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D4 = CLBLM_R_X7Y111_SLICE_X8Y111_AO5;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y111_SLICE_X7Y111_D6 = CLBLM_R_X5Y112_SLICE_X7Y112_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A1 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A2 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_A6 = 1'b1;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B1 = CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B2 = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B3 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B4 = CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_B6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C2 = CLBLM_R_X5Y111_SLICE_X7Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C3 = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C4 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_C6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D1 = CLBLM_R_X5Y111_SLICE_X6Y111_AO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D2 = CLBLL_L_X4Y113_SLICE_X5Y113_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D3 = CLBLM_R_X5Y110_SLICE_X6Y110_BO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D4 = CLBLM_R_X5Y111_SLICE_X6Y111_AO5;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D5 = CLBLM_R_X5Y111_SLICE_X7Y111_CO6;
  assign CLBLM_R_X5Y111_SLICE_X6Y111_D6 = CLBLM_R_X3Y111_SLICE_X3Y111_BO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A1 = CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A2 = CLBLM_R_X7Y107_SLICE_X9Y107_BO5;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_A6 = CLBLL_L_X4Y111_SLICE_X4Y111_AO5;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B2 = CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B5 = CLBLM_R_X5Y112_SLICE_X7Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_B6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_A1 = CLBLL_L_X4Y103_SLICE_X4Y103_AO5;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_A2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_A3 = CLBLM_R_X3Y103_SLICE_X3Y103_CO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C4 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C6 = 1'b1;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_A4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_A5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_A6 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_C2 = 1'b1;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_B2 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_B3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_B4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_B5 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_B6 = CLBLM_R_X5Y102_SLICE_X6Y102_CO6;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D6 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D1 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X7Y112_D2 = 1'b1;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_C1 = 1'b1;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_C2 = 1'b1;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_C3 = 1'b1;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_C4 = 1'b1;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_C5 = 1'b1;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_C6 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A2 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A5 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_A6 = 1'b1;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_D1 = 1'b1;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_D2 = 1'b1;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_D3 = 1'b1;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_D4 = 1'b1;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_D5 = 1'b1;
  assign CLBLM_R_X3Y102_SLICE_X3Y102_D6 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B1 = CLBLM_R_X7Y111_SLICE_X9Y111_BO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_B5 = CLBLL_L_X4Y111_SLICE_X5Y111_CO6;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_A1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C4 = CLBLM_R_X5Y112_SLICE_X6Y112_AO5;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C5 = CLBLM_L_X8Y112_SLICE_X10Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_C6 = CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_A2 = CLBLM_R_X3Y102_SLICE_X3Y102_BO6;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_A3 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_A5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_A6 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_B1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_B2 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_B4 = RIOB33_X105Y111_IOB_X1Y111_I;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_B5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_B6 = CLBLM_R_X3Y102_SLICE_X2Y102_AO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D1 = CLBLM_R_X5Y112_SLICE_X6Y112_AO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D2 = CLBLM_R_X7Y112_SLICE_X9Y112_CO6;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D3 = CLBLL_L_X4Y112_SLICE_X5Y112_CO6;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_C1 = 1'b1;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_C2 = 1'b1;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_C3 = 1'b1;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_C4 = 1'b1;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_C5 = 1'b1;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_C6 = 1'b1;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D5 = CLBLL_L_X4Y112_SLICE_X5Y112_AO5;
  assign CLBLM_R_X5Y112_SLICE_X6Y112_D6 = CLBLM_R_X5Y112_SLICE_X6Y112_BO6;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_D1 = 1'b1;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_D2 = 1'b1;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_D3 = 1'b1;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_D4 = 1'b1;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_D5 = 1'b1;
  assign CLBLM_R_X3Y102_SLICE_X2Y102_D6 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_D1 = CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y136_T1 = 1'b1;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_D1 = CLBLM_R_X3Y107_SLICE_X3Y107_AO6;
  assign LIOI3_X0Y135_OLOGIC_X0Y135_T1 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A1 = CLBLM_R_X3Y104_SLICE_X3Y104_DO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A2 = CLBLL_L_X4Y103_SLICE_X4Y103_AO5;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A5 = CLBLM_R_X3Y103_SLICE_X3Y103_CO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A6 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B1 = CLBLL_L_X4Y103_SLICE_X4Y103_DO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B2 = CLBLL_L_X4Y101_SLICE_X5Y101_AO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B5 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B6 = CLBLL_L_X4Y102_SLICE_X4Y102_AO5;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C2 = CLBLL_L_X4Y102_SLICE_X4Y102_AO5;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C3 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C4 = CLBLL_L_X4Y103_SLICE_X4Y103_DO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C6 = CLBLL_L_X4Y101_SLICE_X5Y101_AO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D2 = CLBLL_L_X2Y103_SLICE_X1Y103_BO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D3 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D5 = CLBLL_L_X4Y102_SLICE_X4Y102_DO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D6 = CLBLL_L_X2Y103_SLICE_X0Y103_AO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A1 = CLBLM_R_X3Y104_SLICE_X2Y104_CO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A2 = CLBLM_R_X3Y103_SLICE_X3Y103_DO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A3 = CLBLM_R_X3Y103_SLICE_X3Y103_AO5;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A4 = CLBLM_R_X3Y103_SLICE_X2Y103_BO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A5 = CLBLL_L_X2Y103_SLICE_X0Y103_CO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A6 = CLBLM_R_X3Y102_SLICE_X3Y102_AO5;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_B5 = CLBLM_R_X11Y105_SLICE_X15Y105_AO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_B6 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B1 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B2 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B3 = CLBLL_L_X2Y103_SLICE_X1Y103_BO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B4 = CLBLL_L_X2Y103_SLICE_X0Y103_AO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B6 = CLBLL_L_X4Y102_SLICE_X4Y102_DO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C1 = CLBLL_L_X2Y103_SLICE_X0Y103_CO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C2 = CLBLM_R_X3Y103_SLICE_X3Y103_AO5;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C3 = CLBLM_R_X3Y103_SLICE_X3Y103_DO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C4 = CLBLM_R_X3Y102_SLICE_X3Y102_AO5;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C5 = CLBLM_R_X3Y104_SLICE_X2Y104_CO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C6 = CLBLM_R_X3Y103_SLICE_X2Y103_BO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D1 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D2 = CLBLM_R_X3Y103_SLICE_X3Y103_AO5;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D3 = CLBLM_R_X3Y103_SLICE_X3Y103_DO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D4 = CLBLM_R_X3Y102_SLICE_X3Y102_AO5;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D5 = CLBLM_R_X3Y104_SLICE_X2Y104_CO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D6 = 1'b1;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_C3 = CLBLM_L_X10Y106_SLICE_X12Y106_CO6;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_C4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_C5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y104_SLICE_X15Y104_C6 = CLBLM_L_X12Y104_SLICE_X16Y104_AO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D4 = CLBLL_L_X4Y105_SLICE_X5Y105_AO5;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_B3 = CLBLM_L_X8Y105_SLICE_X10Y105_BO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C1 = CLBLM_L_X8Y106_SLICE_X10Y106_BO6;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_C2 = CLBLM_L_X8Y105_SLICE_X10Y105_CO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_C6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A1 = CLBLL_L_X4Y106_SLICE_X4Y106_DO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A2 = CLBLL_L_X4Y105_SLICE_X4Y105_BO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A3 = CLBLM_R_X3Y104_SLICE_X2Y104_AO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A4 = CLBLL_L_X4Y104_SLICE_X4Y104_BO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A5 = CLBLL_L_X4Y104_SLICE_X4Y104_BO5;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A6 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B1 = CLBLM_R_X3Y103_SLICE_X3Y103_BO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B2 = CLBLL_L_X4Y101_SLICE_X4Y101_CO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B6 = CLBLL_L_X4Y103_SLICE_X4Y103_BO5;
  assign CLBLM_R_X7Y106_SLICE_X9Y106_D1 = CLBLM_L_X8Y106_SLICE_X10Y106_AO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C1 = CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C2 = CLBLL_L_X4Y105_SLICE_X4Y105_BO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C3 = CLBLL_L_X4Y106_SLICE_X4Y106_DO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C4 = CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C5 = CLBLM_R_X3Y104_SLICE_X2Y104_AO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C6 = CLBLL_L_X4Y106_SLICE_X5Y106_AO5;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D2 = CLBLL_L_X4Y101_SLICE_X4Y101_CO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D4 = CLBLL_L_X4Y103_SLICE_X4Y103_BO5;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D6 = CLBLM_R_X3Y103_SLICE_X3Y103_BO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A2 = CLBLL_L_X4Y104_SLICE_X4Y104_DO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A3 = CLBLM_R_X3Y105_SLICE_X3Y105_BO5;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A4 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A6 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B1 = CLBLL_L_X4Y105_SLICE_X4Y105_DO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B2 = CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B3 = CLBLM_R_X3Y105_SLICE_X3Y105_BO5;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B4 = CLBLL_L_X4Y104_SLICE_X4Y104_BO5;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B5 = CLBLL_L_X4Y104_SLICE_X4Y104_DO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B6 = CLBLM_R_X3Y105_SLICE_X3Y105_CO5;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C1 = CLBLM_R_X3Y103_SLICE_X3Y103_AO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C2 = CLBLM_R_X3Y104_SLICE_X2Y104_AO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C3 = CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C4 = CLBLM_R_X3Y104_SLICE_X2Y104_AO5;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C5 = CLBLL_L_X4Y105_SLICE_X4Y105_DO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C6 = CLBLL_L_X4Y104_SLICE_X4Y104_BO5;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D1 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D2 = CLBLM_R_X3Y104_SLICE_X3Y104_CO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D3 = CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D4 = CLBLM_R_X3Y104_SLICE_X2Y104_AO5;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D5 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D6 = 1'b1;
  assign LIOB33_SING_X0Y149_IOB_X0Y149_O = CLBLL_L_X2Y106_SLICE_X0Y106_AO5;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_D1 = CLBLL_L_X4Y106_SLICE_X4Y106_BO5;
  assign LIOI3_X0Y139_OLOGIC_X0Y140_T1 = 1'b1;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_D1 = CLBLL_L_X4Y106_SLICE_X4Y106_BO6;
  assign LIOI3_X0Y139_OLOGIC_X0Y139_T1 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A1 = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A2 = CLBLL_L_X4Y104_SLICE_X4Y104_AO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A6 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B2 = CLBLL_L_X4Y103_SLICE_X4Y103_BO5;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B5 = CLBLL_L_X4Y101_SLICE_X4Y101_CO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B6 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C2 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C4 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C5 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C6 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D1 = RIOB33_X105Y101_IOB_X1Y102_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D2 = RIOB33_X105Y103_IOB_X1Y103_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D4 = CLBLM_R_X3Y105_SLICE_X3Y105_AO5;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D5 = CLBLL_L_X4Y103_SLICE_X5Y103_CO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D6 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign LIOB33_X0Y117_IOB_X0Y118_O = CLBLL_L_X2Y113_SLICE_X0Y113_AO5;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A1 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A2 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A3 = CLBLM_R_X3Y103_SLICE_X3Y103_AO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A4 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A5 = CLBLM_R_X3Y104_SLICE_X2Y104_BO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A6 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B1 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B2 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B3 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B4 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B5 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B6 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C1 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C2 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C3 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C4 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C5 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C6 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D1 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D2 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D3 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D4 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D5 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D6 = 1'b1;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y108_D = RIOB33_X105Y107_IOB_X1Y108_I;
  assign RIOI3_TBYTESRC_X105Y107_ILOGIC_X1Y107_D = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A1 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A2 = CLBLL_L_X4Y106_SLICE_X4Y106_AO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A4 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A5 = CLBLM_R_X5Y105_SLICE_X6Y105_BO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A6 = 1'b1;
  assign LIOB33_X0Y119_IOB_X0Y119_O = CLBLM_R_X3Y109_SLICE_X2Y109_BO5;
  assign LIOB33_X0Y119_IOB_X0Y120_O = CLBLL_L_X2Y112_SLICE_X0Y112_AO5;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B1 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B2 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B3 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B4 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B5 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B6 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C1 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C2 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C3 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C4 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C5 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C6 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D1 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D2 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D3 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D4 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D5 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D6 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A1 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A2 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A3 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A4 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A5 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A6 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B1 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B2 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B3 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B4 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B5 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B6 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C1 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C2 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C3 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C4 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C5 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C6 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D1 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D2 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D3 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D4 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D5 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D6 = 1'b1;
  assign LIOB33_X0Y121_IOB_X0Y122_O = CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  assign LIOB33_X0Y121_IOB_X0Y121_O = CLBLL_L_X2Y112_SLICE_X0Y112_BO5;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A1 = CLBLM_R_X3Y107_SLICE_X3Y107_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A2 = CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A3 = CLBLM_R_X3Y106_SLICE_X3Y106_AO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A4 = CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A5 = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A6 = CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B1 = CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B2 = CLBLM_R_X3Y107_SLICE_X2Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B3 = CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B4 = CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B5 = CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B6 = CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_D1 = CLBLM_R_X3Y104_SLICE_X3Y104_AO5;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_D = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C1 = CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C2 = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C3 = CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C4 = CLBLM_R_X5Y108_SLICE_X7Y108_BO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C5 = CLBLL_L_X4Y106_SLICE_X4Y106_AO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C6 = CLBLM_R_X5Y105_SLICE_X6Y105_BO6;
  assign LIOI3_X0Y141_OLOGIC_X0Y142_T1 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D1 = CLBLM_R_X5Y105_SLICE_X6Y105_BO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D2 = CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D3 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D4 = CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D5 = CLBLL_L_X4Y106_SLICE_X4Y106_AO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D6 = 1'b1;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_D = LIOB33_X0Y103_IOB_X0Y103_I;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_D1 = CLBLM_R_X3Y104_SLICE_X3Y104_AO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A2 = CLBLM_R_X3Y107_SLICE_X3Y107_DO5;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A4 = CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A6 = 1'b1;
  assign LIOI3_X0Y141_OLOGIC_X0Y141_T1 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B2 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B4 = CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B5 = CLBLM_R_X5Y106_SLICE_X7Y106_DO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C1 = CLBLM_R_X5Y106_SLICE_X7Y106_DO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C6 = CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D1 = CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D2 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D3 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D4 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D5 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D6 = CLBLM_R_X3Y107_SLICE_X2Y107_BO6;
  assign LIOB33_X0Y123_IOB_X0Y124_O = CLBLM_R_X3Y113_SLICE_X2Y113_AO6;
  assign LIOB33_X0Y123_IOB_X0Y123_O = CLBLL_L_X2Y112_SLICE_X1Y112_BO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A1 = CLBLM_R_X3Y107_SLICE_X2Y107_DO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A2 = CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A3 = CLBLM_R_X3Y106_SLICE_X3Y106_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A4 = CLBLM_R_X5Y108_SLICE_X6Y108_DO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A5 = CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A6 = CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B1 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B2 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B3 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B4 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B6 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C1 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C2 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C3 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C4 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C6 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D1 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D2 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D3 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D4 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D6 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A1 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A2 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A3 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A4 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A6 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B1 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B2 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B3 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B4 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B6 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_B5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C1 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C2 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C3 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C4 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C6 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D1 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D2 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D3 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D4 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D6 = 1'b1;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C1 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_R_X11Y105_SLICE_X15Y105_C2 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign LIOB33_X0Y125_IOB_X0Y126_O = CLBLM_R_X3Y113_SLICE_X3Y113_AO6;
  assign LIOB33_X0Y125_IOB_X0Y125_O = CLBLM_R_X3Y112_SLICE_X3Y112_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B4 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_B6 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C3 = CLBLM_L_X10Y108_SLICE_X12Y108_AO6;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_C4 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A1 = CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A2 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A4 = CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D6 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D5 = CLBLM_R_X7Y108_SLICE_X9Y108_BO5;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A1 = CLBLL_L_X2Y111_SLICE_X0Y111_DO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A6 = 1'b1;
  assign CLBLM_R_X7Y107_SLICE_X9Y107_D6 = CLBLM_L_X8Y106_SLICE_X11Y106_AO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D3 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D4 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D6 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_A1 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_A2 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_A3 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_A4 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_A5 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_A6 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_B1 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_B2 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_B3 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_B4 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_B5 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_B6 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_C1 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_C2 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_C3 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_C4 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_C5 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_C6 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_D1 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_D2 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_D3 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_D4 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_D5 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X17Y104_D6 = 1'b1;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_D1 = CLBLM_R_X3Y103_SLICE_X2Y103_AO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_A1 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_A2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_A3 = CLBLM_R_X11Y105_SLICE_X15Y105_AO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_A4 = CLBLM_L_X12Y104_SLICE_X16Y104_BO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_A5 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_A6 = CLBLM_L_X12Y104_SLICE_X16Y104_CO6;
  assign LIOI3_X0Y145_OLOGIC_X0Y146_T1 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_B1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_B2 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_B3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_B4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_B5 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_B6 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_D1 = CLBLM_R_X3Y103_SLICE_X2Y103_DO6;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_C1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_C2 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_C3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_C4 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_C5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_C6 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOI3_X0Y145_OLOGIC_X0Y145_T1 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_D1 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_D2 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_D3 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_D4 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_D5 = 1'b1;
  assign CLBLM_L_X12Y104_SLICE_X16Y104_D6 = 1'b1;
  assign LIOB33_X0Y127_IOB_X0Y128_O = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign LIOB33_X0Y127_IOB_X0Y127_O = CLBLM_R_X3Y111_SLICE_X3Y111_BO5;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A2 = CLBLM_R_X3Y111_SLICE_X3Y111_CO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A4 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A6 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B1 = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B2 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B3 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B4 = CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B6 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C1 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C2 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C3 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C4 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C6 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D1 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D2 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D3 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D4 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D6 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A4 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_B4 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B4 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_L_X8Y101_SLICE_X10Y101_B5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C1 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C2 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C5 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C6 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D2 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D3 = CLBLM_R_X3Y111_SLICE_X3Y111_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D5 = CLBLM_R_X5Y110_SLICE_X6Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign LIOB33_X0Y129_IOB_X0Y130_O = CLBLL_L_X2Y113_SLICE_X0Y113_AO6;
  assign LIOB33_X0Y129_IOB_X0Y129_O = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A1 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A3 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_A6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B1 = CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B2 = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_B6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C2 = CLBLM_R_X5Y111_SLICE_X6Y111_BO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C3 = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C4 = CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_C6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D1 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D2 = CLBLL_L_X4Y111_SLICE_X4Y111_DO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D3 = CLBLM_R_X5Y111_SLICE_X6Y111_DO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D4 = CLBLM_R_X3Y113_SLICE_X3Y113_CO6;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y111_SLICE_X3Y111_D6 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A2 = CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A3 = CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A5 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_A6 = 1'b1;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B3 = CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B5 = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_B6 = CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C1 = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C2 = CLBLM_R_X3Y111_SLICE_X3Y111_AO5;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C3 = CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C4 = CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C5 = CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_C6 = CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D1 = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D2 = CLBLM_R_X3Y111_SLICE_X3Y111_AO5;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D3 = CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D4 = CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D5 = CLBLM_R_X3Y111_SLICE_X3Y111_AO6;
  assign CLBLM_R_X3Y111_SLICE_X2Y111_D6 = CLBLL_L_X2Y111_SLICE_X1Y111_AO6;
  assign LIOB33_X0Y131_IOB_X0Y132_O = CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  assign LIOB33_X0Y131_IOB_X0Y131_O = CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_D1 = CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y148_T1 = 1'b1;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_D1 = CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  assign LIOI3_X0Y147_OLOGIC_X0Y147_T1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A4 = CLBLM_R_X3Y112_SLICE_X3Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_A6 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B2 = CLBLM_R_X3Y112_SLICE_X2Y112_BO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B4 = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B5 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_B6 = CLBLM_R_X3Y112_SLICE_X3Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C2 = CLBLL_L_X4Y111_SLICE_X4Y111_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C5 = CLBLM_R_X3Y112_SLICE_X2Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_C6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D3 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D4 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D5 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y112_SLICE_X3Y112_D6 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A3 = CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A5 = CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_A6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B1 = CLBLL_L_X2Y112_SLICE_X1Y112_CO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B3 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B5 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_B6 = CLBLL_L_X2Y111_SLICE_X1Y111_CO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C1 = CLBLM_R_X3Y111_SLICE_X2Y111_BO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C2 = CLBLL_L_X2Y111_SLICE_X1Y111_DO6;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_C6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D1 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D2 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D3 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D4 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D5 = 1'b1;
  assign CLBLM_R_X3Y112_SLICE_X2Y112_D6 = 1'b1;
  assign LIOB33_X0Y133_IOB_X0Y134_O = 1'b0;
  assign LIOB33_X0Y133_IOB_X0Y133_O = CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A1 = CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A4 = CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_A6 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B4 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B5 = CLBLL_L_X4Y112_SLICE_X4Y112_CO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_B6 = CLBLM_R_X3Y113_SLICE_X2Y113_DO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A4 = CLBLM_R_X11Y106_SLICE_X15Y106_BO6;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A5 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C1 = CLBLL_L_X4Y113_SLICE_X4Y113_AO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C2 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C3 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_A6 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C5 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_C6 = CLBLM_R_X3Y113_SLICE_X3Y113_BO6;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D1 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D2 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D3 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D4 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D5 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X3Y113_D6 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A1 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A2 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A3 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A5 = CLBLM_R_X3Y113_SLICE_X2Y113_CO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_A6 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B1 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B2 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B3 = 1'b1;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_B6 = 1'b1;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B3 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B4 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C1 = CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C3 = CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C4 = RIOB33_SING_X105Y100_IOB_X1Y100_I;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C5 = CLBLL_L_X2Y112_SLICE_X1Y112_CO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_C6 = RIOB33_X105Y105_IOB_X1Y106_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_R_X11Y106_SLICE_X15Y106_B6 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign LIOB33_X0Y135_IOB_X0Y135_O = CLBLM_R_X3Y107_SLICE_X3Y107_AO6;
  assign LIOB33_X0Y135_IOB_X0Y136_O = CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D1 = CLBLM_R_X3Y112_SLICE_X2Y112_AO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D2 = CLBLL_L_X4Y112_SLICE_X4Y112_BO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D3 = CLBLL_L_X2Y112_SLICE_X1Y112_CO6;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D4 = CLBLM_R_X3Y113_SLICE_X2Y113_AO5;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D5 = CLBLM_R_X3Y113_SLICE_X2Y113_BO5;
  assign CLBLM_R_X3Y113_SLICE_X2Y113_D6 = CLBLM_R_X3Y113_SLICE_X2Y113_BO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D4 = CLBLM_L_X10Y110_SLICE_X13Y110_DO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D5 = CLBLM_L_X10Y109_SLICE_X12Y109_AO6;
  assign CLBLM_L_X10Y110_SLICE_X12Y110_D6 = CLBLM_L_X10Y111_SLICE_X12Y111_AO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A1 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_A3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_B1 = 1'b1;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C1 = CLBLM_L_X8Y108_SLICE_X10Y108_AO6;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_C2 = CLBLM_R_X7Y109_SLICE_X9Y109_CO6;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D2 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D3 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D4 = 1'b1;
  assign CLBLM_L_X8Y112_SLICE_X10Y112_D5 = 1'b1;
  assign LIOB33_X0Y137_IOB_X0Y138_O = CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  assign LIOB33_X0Y137_IOB_X0Y137_O = CLBLL_L_X4Y107_SLICE_X4Y107_AO5;
  assign CLBLM_R_X7Y108_SLICE_X9Y108_D6 = 1'b1;
  assign LIOB33_X0Y139_IOB_X0Y140_O = CLBLL_L_X4Y106_SLICE_X4Y106_BO5;
  assign LIOB33_X0Y139_IOB_X0Y139_O = CLBLL_L_X4Y106_SLICE_X4Y106_BO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_B4 = CLBLM_L_X10Y101_SLICE_X12Y101_CO6;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_C1 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_C2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_C3 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X8Y102_SLICE_X10Y102_D5 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign LIOB33_X0Y141_IOB_X0Y142_O = CLBLM_R_X3Y104_SLICE_X3Y104_AO5;
  assign LIOB33_X0Y141_IOB_X0Y141_O = CLBLM_R_X3Y104_SLICE_X3Y104_AO6;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_A1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_A2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_A3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_A4 = RIOB33_X105Y109_IOB_X1Y110_I;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_A5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_A6 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_B1 = RIOB33_X105Y113_IOB_X1Y113_I;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_B2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_B3 = RIOB33_X105Y109_IOB_X1Y109_I;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_B4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_B5 = RIOB33_X105Y111_IOB_X1Y112_I;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_B6 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_D = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_C1 = 1'b1;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_C2 = 1'b1;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_C3 = 1'b1;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_C4 = 1'b1;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_C5 = 1'b1;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_C6 = 1'b1;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_D1 = 1'b1;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_D2 = 1'b1;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_D3 = 1'b1;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_D4 = 1'b1;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_D5 = 1'b1;
  assign CLBLM_L_X10Y101_SLICE_X13Y101_D6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y137_OLOGIC_X0Y138_T1 = 1'b1;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_A1 = CLBLM_L_X8Y102_SLICE_X11Y102_CO6;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_A2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_A3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_A4 = CLBLM_L_X10Y103_SLICE_X13Y103_BO6;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_A5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_A6 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_B1 = CLBLM_L_X8Y102_SLICE_X11Y102_CO6;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_B2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_B3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_B4 = CLBLM_L_X10Y103_SLICE_X13Y103_BO6;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_B5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_B6 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_C1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_C2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_C3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_C4 = CLBLM_R_X11Y103_SLICE_X14Y103_AO6;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_C5 = CLBLM_L_X10Y101_SLICE_X12Y101_DO6;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_C6 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_D1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_D2 = CLBLM_L_X10Y103_SLICE_X13Y103_AO5;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_D3 = CLBLM_L_X8Y102_SLICE_X11Y102_CO6;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_D4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_D5 = CLBLM_L_X8Y102_SLICE_X11Y102_AO5;
  assign CLBLM_L_X10Y101_SLICE_X12Y101_D6 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign LIOB33_X0Y143_IOB_X0Y143_O = CLBLM_R_X3Y104_SLICE_X2Y104_DO6;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_D1 = CLBLL_L_X2Y106_SLICE_X0Y106_AO5;
  assign LIOI3_SING_X0Y149_OLOGIC_X0Y149_T1 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_A2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_A4 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_A5 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_A6 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C3 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C4 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_B1 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_B2 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_B4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_B5 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_B6 = 1'b1;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_C5 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_C1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_C2 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_C3 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_C4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_C5 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_C6 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_D1 = CLBLM_L_X10Y102_SLICE_X13Y102_CO6;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_D2 = CLBLM_R_X7Y102_SLICE_X9Y102_BO6;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_D3 = CLBLM_R_X11Y104_SLICE_X14Y104_DO6;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_D4 = CLBLM_L_X10Y103_SLICE_X13Y103_DO6;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_D5 = CLBLM_L_X10Y102_SLICE_X13Y102_BO5;
  assign CLBLM_L_X10Y102_SLICE_X13Y102_D6 = CLBLM_L_X10Y103_SLICE_X13Y103_BO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_A1 = CLBLM_R_X11Y103_SLICE_X14Y103_AO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_A2 = CLBLM_L_X10Y102_SLICE_X13Y102_BO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_A3 = CLBLM_L_X10Y102_SLICE_X13Y102_AO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_A4 = CLBLM_L_X10Y102_SLICE_X12Y102_BO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_A5 = CLBLM_L_X8Y102_SLICE_X10Y102_AO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_A6 = CLBLM_L_X10Y101_SLICE_X12Y101_AO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_B1 = CLBLM_L_X8Y103_SLICE_X10Y103_CO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_B2 = CLBLM_L_X10Y103_SLICE_X13Y103_BO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_B3 = CLBLM_L_X10Y102_SLICE_X13Y102_CO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_B4 = CLBLM_R_X7Y102_SLICE_X9Y102_AO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_B5 = CLBLM_R_X7Y102_SLICE_X9Y102_BO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_B6 = CLBLL_L_X4Y103_SLICE_X4Y103_AO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D1 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_C1 = CLBLM_L_X8Y102_SLICE_X10Y102_AO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_C2 = CLBLM_L_X10Y101_SLICE_X12Y101_AO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_C3 = CLBLM_L_X10Y102_SLICE_X13Y102_AO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_C4 = CLBLM_L_X10Y102_SLICE_X13Y102_BO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_C5 = CLBLM_R_X11Y103_SLICE_X14Y103_AO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_C6 = CLBLM_L_X10Y102_SLICE_X12Y102_BO6;
  assign CLBLM_L_X10Y111_SLICE_X13Y111_D4 = 1'b1;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_D1 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_D2 = CLBLM_L_X10Y101_SLICE_X12Y101_AO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_D3 = CLBLM_R_X11Y103_SLICE_X14Y103_AO6;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_D4 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_D5 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y102_SLICE_X12Y102_D6 = CLBLM_L_X10Y102_SLICE_X12Y102_BO6;
  assign LIOB33_X0Y145_IOB_X0Y146_O = CLBLM_R_X3Y103_SLICE_X2Y103_AO6;
  assign LIOB33_X0Y145_IOB_X0Y145_O = CLBLM_R_X3Y103_SLICE_X2Y103_DO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_B6 = CLBLM_L_X10Y110_SLICE_X13Y110_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B1 = CLBLM_L_X10Y106_SLICE_X13Y106_AO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C5 = CLBLM_L_X10Y111_SLICE_X12Y111_DO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_B2 = CLBLM_R_X11Y108_SLICE_X15Y108_BO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_C6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A1 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A2 = CLBLM_L_X12Y104_SLICE_X16Y104_BO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A4 = CLBLM_L_X10Y101_SLICE_X13Y101_BO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A5 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_A6 = 1'b1;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B1 = CLBLM_L_X10Y101_SLICE_X13Y101_AO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B2 = CLBLM_L_X12Y104_SLICE_X16Y104_BO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B3 = CLBLM_L_X10Y102_SLICE_X13Y102_CO5;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B4 = CLBLM_R_X5Y101_SLICE_X7Y101_AO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B5 = CLBLM_L_X10Y101_SLICE_X13Y101_BO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_B6 = CLBLL_L_X4Y103_SLICE_X4Y103_BO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D2 = CLBLM_L_X10Y110_SLICE_X13Y110_CO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C5 = CLBLM_R_X11Y108_SLICE_X15Y108_BO6;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C4 = CLBLM_R_X11Y105_SLICE_X15Y105_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D3 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C2 = CLBLM_L_X12Y104_SLICE_X16Y104_BO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C4 = RIOB33_X105Y107_IOB_X1Y108_I;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C5 = CLBLM_L_X10Y101_SLICE_X13Y101_AO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D4 = RIOB33_X105Y101_IOB_X1Y101_I;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C6 = CLBLM_L_X10Y101_SLICE_X13Y101_BO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_C3 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X11Y107_SLICE_X15Y107_C6 = CLBLM_R_X11Y106_SLICE_X15Y106_CO6;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_L_X10Y111_SLICE_X12Y111_D6 = CLBLM_L_X8Y111_SLICE_X11Y111_BO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D1 = CLBLM_L_X10Y101_SLICE_X13Y101_BO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D2 = CLBLM_R_X5Y101_SLICE_X7Y101_AO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D3 = CLBLL_L_X4Y103_SLICE_X4Y103_BO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D4 = CLBLM_L_X10Y102_SLICE_X13Y102_CO5;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D6 = CLBLM_L_X12Y104_SLICE_X16Y104_BO6;
  assign CLBLM_L_X10Y103_SLICE_X13Y103_D5 = CLBLM_L_X10Y101_SLICE_X13Y101_AO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A1 = CLBLM_L_X10Y102_SLICE_X12Y102_DO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A4 = CLBLM_L_X10Y104_SLICE_X13Y104_AO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_A6 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B1 = CLBLM_L_X10Y102_SLICE_X12Y102_DO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B3 = RIOB33_X105Y105_IOB_X1Y105_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B4 = CLBLM_R_X11Y103_SLICE_X14Y103_BO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B5 = RIOB33_X105Y103_IOB_X1Y104_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_B6 = CLBLM_L_X10Y103_SLICE_X12Y103_CO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C1 = RIOB33_X105Y107_IOB_X1Y107_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C2 = CLBLM_L_X10Y101_SLICE_X12Y101_DO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C3 = CLBLM_R_X11Y103_SLICE_X14Y103_AO6;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C4 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_L_X10Y103_SLICE_X12Y103_C5 = RIOB33_X105Y105_IOB_X1Y105_I;
endmodule
