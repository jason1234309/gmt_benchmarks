module top(
  input LIOB33_SING_X0Y100_IOB_X0Y100_IPAD,
  input LIOB33_X0Y101_IOB_X0Y101_IPAD,
  input LIOB33_X0Y101_IOB_X0Y102_IPAD,
  input LIOB33_X0Y103_IOB_X0Y103_IPAD,
  input LIOB33_X0Y103_IOB_X0Y104_IPAD,
  input LIOB33_X0Y105_IOB_X0Y105_IPAD,
  input LIOB33_X0Y105_IOB_X0Y106_IPAD,
  input LIOB33_X0Y107_IOB_X0Y107_IPAD,
  input LIOB33_X0Y107_IOB_X0Y108_IPAD,
  input LIOB33_X0Y109_IOB_X0Y109_IPAD,
  input LIOB33_X0Y109_IOB_X0Y110_IPAD,
  input LIOB33_X0Y111_IOB_X0Y111_IPAD,
  input LIOB33_X0Y111_IOB_X0Y112_IPAD,
  input LIOB33_X0Y113_IOB_X0Y113_IPAD,
  input LIOB33_X0Y113_IOB_X0Y114_IPAD,
  input LIOB33_X0Y115_IOB_X0Y115_IPAD,
  input LIOB33_X0Y115_IOB_X0Y116_IPAD,
  input LIOB33_X0Y117_IOB_X0Y117_IPAD,
  input LIOB33_X0Y117_IOB_X0Y118_IPAD,
  input LIOB33_X0Y127_IOB_X0Y128_IPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD
  );
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A1;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A2;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A3;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A4;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_AO5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_AO6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_AQ;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A_CY;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_A_XOR;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B1;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B2;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B3;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B4;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_BO5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_BO6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_BQ;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B_CY;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_B_XOR;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C1;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C2;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C3;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C4;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_CLK;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_CO5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_CO6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C_CY;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_C_XOR;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D1;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D2;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D3;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D4;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_DO5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_DO6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D_CY;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X0Y103_D_XOR;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A1;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A2;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A3;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A4;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_AO5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_AO6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_AQ;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A_CY;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_A_XOR;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B1;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B2;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B3;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B4;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_BO5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_BO6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_BQ;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B_CY;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_B_XOR;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C1;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C2;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C3;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C4;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_CLK;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_CMUX;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_CO5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_CO6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C_CY;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_C_XOR;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D1;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D2;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D3;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D4;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_DO5;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_DO6;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D_CY;
  wire [0:0] CLBLL_L_X2Y103_SLICE_X1Y103_D_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_AO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_AO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_AQ;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_A_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_BO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_BO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_BQ;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_B_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_CLK;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_CMUX;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_CO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_CO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_C_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_DO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_DO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X0Y104_D_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_AMUX;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_AO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_AO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_A_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_BO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_BO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_B_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_CO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_CO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_C_XOR;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D1;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D2;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D3;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D4;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_DO5;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_DO6;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D_CY;
  wire [0:0] CLBLL_L_X2Y104_SLICE_X1Y104_D_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_AO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_AO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_AQ;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_BO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_BO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_BQ;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_CLK;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_CO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_CO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_CQ;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_DO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_DO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_DQ;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_AMUX;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_AO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_AO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_BO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_BO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_BQ;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_CLK;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_CO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_CO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_DO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_DO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_AMUX;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_AO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_BO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_BQ;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_CLK;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_CMUX;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_CO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_DO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_DO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A5Q;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_AMUX;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_AO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_AQ;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_AX;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_BO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_BQ;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_CLK;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_CMUX;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_CO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_CO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_DO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_DO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_AMUX;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_AO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_BO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_BO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_BQ;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_CLK;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_CO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_CO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_CQ;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_DMUX;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_DO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_DO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_AO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_AQ;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_BO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_BO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_BQ;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_CLK;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_CO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_CO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_CQ;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_DMUX;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_DO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_DO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A5Q;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_AMUX;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_AO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_AQ;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_AX;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_BMUX;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_BO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_BO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_BQ;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_BX;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_CLK;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_CO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_DO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_DO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_AO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_BO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_CO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_CO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_DO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_AO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_AO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_AQ;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_A_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_BO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_BO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_B_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_CLK;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_CO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_CO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_C_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_DO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_DO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X4Y103_D_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_AO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_AO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_AQ;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_A_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_BO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_BO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_BQ;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_B_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_CLK;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_CO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_CO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_CQ;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_C_XOR;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D1;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D2;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D3;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D4;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_DO5;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_DO6;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D_CY;
  wire [0:0] CLBLL_L_X4Y103_SLICE_X5Y103_D_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_AO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_AO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_AQ;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_BO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_BO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_BQ;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_CLK;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_CMUX;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_CO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_DO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_DO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_AMUX;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_AO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_AO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_AQ;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_BMUX;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_BO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_BO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_CLK;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_CO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_CO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_DO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_DO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_AO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_AO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_AQ;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_BO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_BO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_CLK;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_CO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_DO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_DO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_AO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_AO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_AQ;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_BO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_BQ;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_CLK;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_CO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_CO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_CQ;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_DO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_DO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_AMUX;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_AO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_AO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_AQ;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_AX;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_BMUX;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_BO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_BO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_CLK;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_CMUX;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_CO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_DO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_DO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_AO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_AO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_AQ;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_BO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_BO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_CLK;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_CO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_CO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_DO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_DO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_AO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_AQ;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_BO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_BQ;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_CLK;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_CO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_CQ;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_DO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_DO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_AO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_AO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_AQ;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_BO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_BQ;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_CLK;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_CO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_DO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_AO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_AO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_AQ;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_A_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_BO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_BO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_BQ;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_B_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_CLK;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_CO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_CO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_CQ;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_C_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_DO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_DO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X2Y103_D_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_AO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_AO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_AQ;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_A_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_BO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_BO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_BQ;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_B_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_CLK;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_CO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_CO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_C_XOR;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D1;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D2;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D3;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D4;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_DO5;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_DO6;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D_CY;
  wire [0:0] CLBLM_R_X3Y103_SLICE_X3Y103_D_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_AO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_AO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_AQ;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_BO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_BO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_BQ;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_CLK;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_CO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_CO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_DO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_DO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_AO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_AO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_AQ;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_BO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_BQ;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_CLK;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_CO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_CO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_DO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_DO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A5Q;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_AMUX;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_AO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_AQ;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_AX;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B5Q;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_BMUX;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_BO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_BO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_BQ;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_BX;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_CLK;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_CMUX;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_CO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_CO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_DMUX;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_DO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_DO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_AO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_AO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_AQ;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_BO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_CLK;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_CO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_DO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_DO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_AMUX;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_AO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_AO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_AQ;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_BO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_BO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_BQ;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_CLK;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_CMUX;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_CO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_DO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_DO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_AMUX;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_AO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_AO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_BO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_CO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_CO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_DO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_DO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_AO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_AQ;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_BO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_BO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_BQ;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_CLK;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_CO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_DO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_DO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_AMUX;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_AO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_AO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_BMUX;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_BO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_BO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_CO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_DMUX;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_DO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_DO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D_XOR;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A1;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A2;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A3;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A4;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_AO5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_AO6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_AQ;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A_CY;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_A_XOR;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B1;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B2;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B3;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B4;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_BO5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_BO6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_BQ;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B_CY;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_B_XOR;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C1;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C2;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C3;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C4;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_CLK;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_CO5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_CO6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_CQ;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C_CY;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_C_XOR;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D1;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D2;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D3;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D4;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_DO5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_DO6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D_CY;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X6Y103_D_XOR;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A1;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A2;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A3;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A4;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_AO5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_AO6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A_CY;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_A_XOR;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B1;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B2;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B3;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B4;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_BO5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_BO6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B_CY;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_B_XOR;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C1;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C2;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C3;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C4;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_CO5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_CO6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C_CY;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_C_XOR;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D1;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D2;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D3;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D4;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_DO5;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_DO6;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D_CY;
  wire [0:0] CLBLM_R_X5Y103_SLICE_X7Y103_D_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_AO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_AO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_AQ;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_A_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_BO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_BO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_BQ;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_B_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_CLK;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_CO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_CO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_C_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_DO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_DO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X6Y104_D_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_AO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_AO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_AQ;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_A_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_BO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_BO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_BQ;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_B_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_CLK;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_CO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_CO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_C_XOR;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D1;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D2;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D3;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D4;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_DO5;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_DO6;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D_CY;
  wire [0:0] CLBLM_R_X5Y104_SLICE_X7Y104_D_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_AO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_AQ;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_BO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_BO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_BQ;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_CLK;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_CMUX;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_CO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_CO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_DO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_DO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_AO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_AO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_AQ;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_BO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_BO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_CLK;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_CO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_DO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_DO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_AMUX;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_AO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_BO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_CO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_DO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_AO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_AO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_AQ;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_BO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_CLK;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_CO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_CO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_DO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_DO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_AO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_AQ;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_A_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_BO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_BQ;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_B_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_CLK;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_CO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_CO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_CQ;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_C_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_DO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_DQ;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X6Y107_D_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_AO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_AO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_A_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_BO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_B_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_CO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_CO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_C_XOR;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D1;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D2;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D3;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D4;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_DO5;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_DO6;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D_CY;
  wire [0:0] CLBLM_R_X5Y107_SLICE_X7Y107_D_XOR;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_I;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_I;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_D;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_O;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y118_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y118_O;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_D;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_O;


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y103_SLICE_X0Y103_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y103_SLICE_X0Y103_AO6),
.Q(CLBLL_L_X2Y103_SLICE_X0Y103_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y103_SLICE_X0Y103_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y103_SLICE_X0Y103_BO6),
.Q(CLBLL_L_X2Y103_SLICE_X0Y103_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0455040004550400)
  ) CLBLL_L_X2Y103_SLICE_X0Y103_DLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(CLBLL_L_X2Y106_SLICE_X1Y106_BQ),
.I3(CLBLL_L_X2Y104_SLICE_X0Y104_CO5),
.I4(CLBLL_L_X2Y103_SLICE_X0Y103_BQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y103_SLICE_X0Y103_DO5),
.O6(CLBLL_L_X2Y103_SLICE_X0Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0455045504000400)
  ) CLBLL_L_X2Y103_SLICE_X0Y103_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(CLBLL_L_X2Y106_SLICE_X1Y106_BQ),
.I3(CLBLL_L_X2Y104_SLICE_X0Y104_CO5),
.I4(1'b1),
.I5(CLBLL_L_X2Y103_SLICE_X0Y103_AQ),
.O5(CLBLL_L_X2Y103_SLICE_X0Y103_CO5),
.O6(CLBLL_L_X2Y103_SLICE_X0Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefaeeaafafaaaaa)
  ) CLBLL_L_X2Y103_SLICE_X0Y103_BLUT (
.I0(CLBLL_L_X2Y103_SLICE_X0Y103_DO6),
.I1(CLBLL_L_X2Y104_SLICE_X0Y104_CO6),
.I2(CLBLL_L_X2Y103_SLICE_X0Y103_AQ),
.I3(CLBLL_L_X2Y106_SLICE_X1Y106_BQ),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(LIOB33_X0Y111_IOB_X0Y111_I),
.O5(CLBLL_L_X2Y103_SLICE_X0Y103_BO5),
.O6(CLBLL_L_X2Y103_SLICE_X0Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffeca0a0a0)
  ) CLBLL_L_X2Y103_SLICE_X0Y103_ALUT (
.I0(CLBLL_L_X2Y104_SLICE_X0Y104_AQ),
.I1(CLBLL_L_X2Y104_SLICE_X0Y104_CO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLL_L_X2Y106_SLICE_X1Y106_BQ),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(CLBLL_L_X2Y103_SLICE_X0Y103_CO6),
.O5(CLBLL_L_X2Y103_SLICE_X0Y103_AO5),
.O6(CLBLL_L_X2Y103_SLICE_X0Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y103_SLICE_X1Y103_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y103_SLICE_X1Y103_AO6),
.Q(CLBLL_L_X2Y103_SLICE_X1Y103_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y103_SLICE_X1Y103_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y103_SLICE_X1Y103_BO6),
.Q(CLBLL_L_X2Y103_SLICE_X1Y103_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5faf5faf5faf5af)
  ) CLBLL_L_X2Y103_SLICE_X1Y103_DLUT (
.I0(CLBLL_L_X2Y103_SLICE_X0Y103_AQ),
.I1(1'b1),
.I2(CLBLL_L_X2Y104_SLICE_X0Y104_AQ),
.I3(CLBLM_R_X3Y103_SLICE_X2Y103_CQ),
.I4(CLBLL_L_X2Y104_SLICE_X0Y104_BQ),
.I5(CLBLL_L_X2Y103_SLICE_X0Y103_BQ),
.O5(CLBLL_L_X2Y103_SLICE_X1Y103_DO5),
.O6(CLBLL_L_X2Y103_SLICE_X1Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hddffeeffffddffee)
  ) CLBLL_L_X2Y103_SLICE_X1Y103_CLUT (
.I0(CLBLL_L_X2Y103_SLICE_X1Y103_BQ),
.I1(CLBLL_L_X2Y103_SLICE_X1Y103_DO6),
.I2(1'b1),
.I3(CLBLL_L_X2Y103_SLICE_X1Y103_AQ),
.I4(CLBLL_L_X2Y104_SLICE_X0Y104_BQ),
.I5(CLBLL_L_X2Y103_SLICE_X0Y103_BQ),
.O5(CLBLL_L_X2Y103_SLICE_X1Y103_CO5),
.O6(CLBLL_L_X2Y103_SLICE_X1Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f08822f0f00000)
  ) CLBLL_L_X2Y103_SLICE_X1Y103_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLL_L_X2Y103_SLICE_X1Y103_BQ),
.I2(CLBLL_L_X2Y103_SLICE_X1Y103_AQ),
.I3(CLBLL_L_X2Y104_SLICE_X1Y104_AO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLL_L_X2Y103_SLICE_X1Y103_CO6),
.O5(CLBLL_L_X2Y103_SLICE_X1Y103_BO5),
.O6(CLBLL_L_X2Y103_SLICE_X1Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa78aa00aa00aa00)
  ) CLBLL_L_X2Y103_SLICE_X1Y103_ALUT (
.I0(CLBLM_R_X3Y103_SLICE_X2Y103_CQ),
.I1(CLBLM_R_X3Y103_SLICE_X3Y103_CO6),
.I2(CLBLL_L_X2Y103_SLICE_X1Y103_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLL_L_X2Y103_SLICE_X1Y103_CO6),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLL_L_X2Y103_SLICE_X1Y103_AO5),
.O6(CLBLL_L_X2Y103_SLICE_X1Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y104_SLICE_X0Y104_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y104_SLICE_X0Y104_AO6),
.Q(CLBLL_L_X2Y104_SLICE_X0Y104_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y104_SLICE_X0Y104_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y104_SLICE_X0Y104_BO6),
.Q(CLBLL_L_X2Y104_SLICE_X0Y104_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0055000000f500a0)
  ) CLBLL_L_X2Y104_SLICE_X0Y104_DLUT (
.I0(CLBLL_L_X2Y104_SLICE_X0Y104_CO5),
.I1(1'b1),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLL_L_X2Y104_SLICE_X0Y104_BQ),
.I5(CLBLL_L_X2Y106_SLICE_X1Y106_BQ),
.O5(CLBLL_L_X2Y104_SLICE_X0Y104_DO5),
.O6(CLBLL_L_X2Y104_SLICE_X0Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0155015503ff03ff)
  ) CLBLL_L_X2Y104_SLICE_X0Y104_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLL_L_X2Y103_SLICE_X1Y103_CO6),
.I2(CLBLL_L_X2Y105_SLICE_X0Y105_BQ),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y104_SLICE_X0Y104_CO5),
.O6(CLBLL_L_X2Y104_SLICE_X0Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeeefaaaeeeeaaaa)
  ) CLBLL_L_X2Y104_SLICE_X0Y104_BLUT (
.I0(CLBLL_L_X2Y104_SLICE_X0Y104_DO6),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y111_IOB_X0Y112_I),
.I3(CLBLL_L_X2Y106_SLICE_X1Y106_BQ),
.I4(CLBLL_L_X2Y103_SLICE_X0Y103_BQ),
.I5(CLBLL_L_X2Y104_SLICE_X0Y104_CO6),
.O5(CLBLL_L_X2Y104_SLICE_X0Y104_BO5),
.O6(CLBLL_L_X2Y104_SLICE_X0Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff0084c0ff000000)
  ) CLBLL_L_X2Y104_SLICE_X0Y104_ALUT (
.I0(CLBLL_L_X2Y104_SLICE_X1Y104_AO6),
.I1(CLBLL_L_X2Y103_SLICE_X1Y103_CO6),
.I2(CLBLL_L_X2Y104_SLICE_X0Y104_AQ),
.I3(CLBLL_L_X2Y103_SLICE_X1Y103_BQ),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLL_L_X2Y104_SLICE_X0Y104_AO5),
.O6(CLBLL_L_X2Y104_SLICE_X0Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffbfffffaaeaaaaa)
  ) CLBLL_L_X2Y104_SLICE_X1Y104_DLUT (
.I0(CLBLL_L_X2Y105_SLICE_X1Y105_AO6),
.I1(CLBLM_R_X3Y103_SLICE_X3Y103_CO6),
.I2(CLBLL_L_X2Y103_SLICE_X1Y103_BQ),
.I3(CLBLL_L_X2Y104_SLICE_X1Y104_AO5),
.I4(CLBLM_R_X5Y104_SLICE_X6Y104_DO6),
.I5(CLBLM_R_X3Y103_SLICE_X3Y103_DO6),
.O5(CLBLL_L_X2Y104_SLICE_X1Y104_DO5),
.O6(CLBLL_L_X2Y104_SLICE_X1Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff7fffff0f8f0f0)
  ) CLBLL_L_X2Y104_SLICE_X1Y104_CLUT (
.I0(CLBLL_L_X2Y103_SLICE_X1Y103_BQ),
.I1(CLBLM_R_X3Y103_SLICE_X3Y103_CO6),
.I2(CLBLL_L_X2Y105_SLICE_X1Y105_AO5),
.I3(CLBLL_L_X2Y104_SLICE_X1Y104_AO5),
.I4(CLBLM_R_X5Y104_SLICE_X6Y104_DO6),
.I5(CLBLM_R_X3Y103_SLICE_X3Y103_DO6),
.O5(CLBLL_L_X2Y104_SLICE_X1Y104_CO5),
.O6(CLBLL_L_X2Y104_SLICE_X1Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h78f0f0f0f0f0f0f0)
  ) CLBLL_L_X2Y104_SLICE_X1Y104_BLUT (
.I0(CLBLM_R_X3Y103_SLICE_X2Y103_CQ),
.I1(CLBLM_R_X3Y103_SLICE_X3Y103_CO6),
.I2(CLBLM_R_X3Y103_SLICE_X3Y103_DO6),
.I3(CLBLL_L_X2Y103_SLICE_X1Y103_BQ),
.I4(CLBLL_L_X2Y103_SLICE_X1Y103_AQ),
.I5(CLBLM_R_X5Y104_SLICE_X6Y104_DO6),
.O5(CLBLL_L_X2Y104_SLICE_X1Y104_BO5),
.O6(CLBLL_L_X2Y104_SLICE_X1Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f7f7f7f5f5f5f5f)
  ) CLBLL_L_X2Y104_SLICE_X1Y104_ALUT (
.I0(CLBLM_R_X3Y103_SLICE_X2Y103_CQ),
.I1(CLBLM_R_X3Y103_SLICE_X3Y103_CO6),
.I2(CLBLL_L_X2Y103_SLICE_X1Y103_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y104_SLICE_X1Y104_AO5),
.O6(CLBLL_L_X2Y104_SLICE_X1Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y105_SLICE_X0Y105_AO6),
.Q(CLBLL_L_X2Y105_SLICE_X0Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y105_SLICE_X0Y105_BO6),
.Q(CLBLL_L_X2Y105_SLICE_X0Y105_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y105_SLICE_X0Y105_CO6),
.Q(CLBLL_L_X2Y105_SLICE_X0Y105_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y105_SLICE_X0Y105_DO6),
.Q(CLBLL_L_X2Y105_SLICE_X0Y105_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff109800001098)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_DLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(CLBLL_L_X2Y105_SLICE_X0Y105_DQ),
.I3(CLBLM_R_X3Y104_SLICE_X2Y104_BQ),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLL_L_X2Y105_SLICE_X1Y105_BQ),
.O5(CLBLL_L_X2Y105_SLICE_X0Y105_DO5),
.O6(CLBLL_L_X2Y105_SLICE_X0Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff0f0f4f0fef0)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_CLUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(CLBLL_L_X2Y105_SLICE_X0Y105_CQ),
.I2(CLBLM_R_X3Y105_SLICE_X2Y105_CO6),
.I3(CLBLM_R_X3Y105_SLICE_X2Y105_B5Q),
.I4(CLBLL_L_X2Y105_SLICE_X0Y105_BQ),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLL_L_X2Y105_SLICE_X0Y105_CO5),
.O6(CLBLL_L_X2Y105_SLICE_X0Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffbaaaaaafbaa)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_BLUT (
.I0(CLBLM_R_X3Y105_SLICE_X2Y105_CO6),
.I1(CLBLL_L_X2Y105_SLICE_X0Y105_BQ),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(CLBLM_R_X3Y105_SLICE_X2Y105_B5Q),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_R_X3Y104_SLICE_X2Y104_BQ),
.O5(CLBLL_L_X2Y105_SLICE_X0Y105_BO5),
.O6(CLBLL_L_X2Y105_SLICE_X0Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb888b88888aa88aa)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_ALUT (
.I0(CLBLL_L_X2Y106_SLICE_X1Y106_A5Q),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLL_L_X2Y105_SLICE_X0Y105_AQ),
.I3(CLBLL_L_X2Y103_SLICE_X1Y103_CO6),
.I4(1'b1),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLL_L_X2Y105_SLICE_X0Y105_AO5),
.O6(CLBLL_L_X2Y105_SLICE_X0Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y105_SLICE_X1Y105_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y105_SLICE_X1Y105_BO6),
.Q(CLBLL_L_X2Y105_SLICE_X1Y105_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000055555555)
  ) CLBLL_L_X2Y105_SLICE_X1Y105_DLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(CLBLL_L_X2Y105_SLICE_X0Y105_BQ),
.O5(CLBLL_L_X2Y105_SLICE_X1Y105_DO5),
.O6(CLBLL_L_X2Y105_SLICE_X1Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ff00ff0a)
  ) CLBLL_L_X2Y105_SLICE_X1Y105_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y108_I),
.I1(1'b1),
.I2(CLBLL_L_X4Y107_SLICE_X5Y107_DO6),
.I3(CLBLL_L_X2Y105_SLICE_X0Y105_BQ),
.I4(CLBLL_L_X2Y105_SLICE_X0Y105_AQ),
.I5(CLBLM_R_X3Y105_SLICE_X2Y105_AQ),
.O5(CLBLL_L_X2Y105_SLICE_X1Y105_CO5),
.O6(CLBLL_L_X2Y105_SLICE_X1Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa0ff00ffe0ffc0)
  ) CLBLL_L_X2Y105_SLICE_X1Y105_BLUT (
.I0(CLBLL_L_X2Y105_SLICE_X1Y105_DO6),
.I1(CLBLL_L_X2Y104_SLICE_X1Y104_DO6),
.I2(CLBLL_L_X2Y106_SLICE_X0Y106_CO5),
.I3(CLBLM_R_X3Y105_SLICE_X3Y105_CO6),
.I4(CLBLL_L_X2Y104_SLICE_X1Y104_CO6),
.I5(CLBLL_L_X2Y105_SLICE_X1Y105_CO6),
.O5(CLBLL_L_X2Y105_SLICE_X1Y105_BO5),
.O6(CLBLL_L_X2Y105_SLICE_X1Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000aa22222222)
  ) CLBLL_L_X2Y105_SLICE_X1Y105_ALUT (
.I0(CLBLM_R_X3Y106_SLICE_X3Y106_CO6),
.I1(LIOB33_X0Y111_IOB_X0Y112_I),
.I2(1'b1),
.I3(CLBLM_R_X3Y105_SLICE_X2Y105_AQ),
.I4(CLBLL_L_X4Y107_SLICE_X5Y107_DO6),
.I5(1'b1),
.O5(CLBLL_L_X2Y105_SLICE_X1Y105_AO5),
.O6(CLBLL_L_X2Y105_SLICE_X1Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y106_SLICE_X0Y106_BO6),
.Q(CLBLL_L_X2Y106_SLICE_X0Y106_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8888888800808880)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_DLUT (
.I0(CLBLM_R_X3Y105_SLICE_X2Y105_AQ),
.I1(CLBLL_L_X2Y106_SLICE_X1Y106_CO6),
.I2(CLBLL_L_X2Y106_SLICE_X1Y106_AQ),
.I3(CLBLL_L_X2Y105_SLICE_X0Y105_BQ),
.I4(LIOB33_X0Y115_IOB_X0Y115_I),
.I5(CLBLL_L_X2Y107_SLICE_X0Y107_BQ),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_DO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00be1450500000)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLL_L_X2Y108_SLICE_X0Y108_BQ),
.I2(CLBLM_R_X3Y106_SLICE_X3Y106_DO6),
.I3(CLBLL_L_X2Y108_SLICE_X0Y108_A5Q),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_CO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf222f222f000f000)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_BLUT (
.I0(CLBLL_L_X2Y106_SLICE_X0Y106_DO6),
.I1(CLBLL_L_X2Y104_SLICE_X1Y104_BO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLL_L_X2Y105_SLICE_X0Y105_DQ),
.I4(1'b1),
.I5(CLBLL_L_X2Y106_SLICE_X0Y106_AO5),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_BO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00fa00ccaafaaaff)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_ALUT (
.I0(CLBLL_L_X2Y107_SLICE_X0Y107_CQ),
.I1(CLBLL_L_X2Y107_SLICE_X0Y107_BQ),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(CLBLL_L_X2Y105_SLICE_X0Y105_BQ),
.I4(CLBLL_L_X2Y106_SLICE_X1Y106_AQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_AO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y106_SLICE_X1Y106_CO5),
.Q(CLBLL_L_X2Y106_SLICE_X1Y106_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y106_SLICE_X1Y106_AO6),
.Q(CLBLL_L_X2Y106_SLICE_X1Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y106_SLICE_X1Y106_BO6),
.Q(CLBLL_L_X2Y106_SLICE_X1Y106_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcd01cc00cd01ff33)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_DLUT (
.I0(LIOB33_X0Y115_IOB_X0Y115_I),
.I1(CLBLL_L_X2Y105_SLICE_X0Y105_BQ),
.I2(CLBLL_L_X2Y107_SLICE_X0Y107_CQ),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(CLBLL_L_X2Y106_SLICE_X1Y106_AQ),
.I5(CLBLL_L_X2Y107_SLICE_X0Y107_BQ),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_DO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h05050505fbab5101)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLL_L_X2Y103_SLICE_X1Y103_CO6),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLL_L_X2Y106_SLICE_X1Y106_A5Q),
.I4(CLBLL_L_X2Y106_SLICE_X1Y106_AQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_CO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f00000ccff)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y106_SLICE_X1Y106_BQ),
.I2(CLBLL_L_X4Y104_SLICE_X5Y104_AQ),
.I3(CLBLL_L_X2Y104_SLICE_X1Y104_BO6),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_BO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcacac0c0c0c0cccc)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_ALUT (
.I0(CLBLL_L_X2Y106_SLICE_X1Y106_AQ),
.I1(CLBLL_L_X2Y106_SLICE_X1Y106_BQ),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(1'b1),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLL_L_X2Y103_SLICE_X1Y103_CO6),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_AO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y107_SLICE_X0Y107_BO6),
.Q(CLBLL_L_X2Y107_SLICE_X0Y107_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y107_SLICE_X0Y107_CO6),
.Q(CLBLL_L_X2Y107_SLICE_X0Y107_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h07050705080a080a)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLL_L_X2Y103_SLICE_X1Y103_CO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLL_L_X2Y105_SLICE_X0Y105_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_DO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeeefcccfaaaf000)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_CLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(CLBLL_L_X2Y107_SLICE_X0Y107_CQ),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLL_L_X2Y107_SLICE_X0Y107_BQ),
.I4(CLBLL_L_X2Y107_SLICE_X0Y107_DO6),
.I5(CLBLL_L_X2Y107_SLICE_X0Y107_DO5),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_CO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeca0eca0eca0)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_BLUT (
.I0(CLBLL_L_X2Y107_SLICE_X0Y107_DO6),
.I1(CLBLL_L_X2Y107_SLICE_X0Y107_BQ),
.I2(LIOB33_X0Y101_IOB_X0Y102_I),
.I3(CLBLL_L_X2Y107_SLICE_X0Y107_DO5),
.I4(CLBLM_R_X3Y105_SLICE_X2Y105_AQ),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_BO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff005f005f00)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_ALUT (
.I0(CLBLL_L_X2Y103_SLICE_X1Y103_CO6),
.I1(1'b1),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLL_L_X2Y105_SLICE_X0Y105_BQ),
.I4(LIOB33_X0Y109_IOB_X0Y110_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_AO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y107_SLICE_X1Y107_AO6),
.Q(CLBLL_L_X2Y107_SLICE_X1Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y107_SLICE_X1Y107_BO6),
.Q(CLBLL_L_X2Y107_SLICE_X1Y107_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y107_SLICE_X1Y107_CO6),
.Q(CLBLL_L_X2Y107_SLICE_X1Y107_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000aeaa51555155)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_DLUT (
.I0(CLBLL_L_X2Y105_SLICE_X0Y105_BQ),
.I1(CLBLL_L_X2Y103_SLICE_X1Y103_CO6),
.I2(LIOB33_X0Y115_IOB_X0Y116_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_DO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hefffaa00ba00aa00)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_R_X3Y106_SLICE_X2Y106_AO5),
.I2(CLBLL_L_X2Y107_SLICE_X1Y107_BQ),
.I3(CLBLL_L_X2Y107_SLICE_X1Y107_AQ),
.I4(CLBLL_L_X2Y107_SLICE_X1Y107_DO6),
.I5(CLBLL_L_X2Y107_SLICE_X1Y107_CQ),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_CO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf888f888f222f222)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_BLUT (
.I0(CLBLL_L_X2Y107_SLICE_X1Y107_DO6),
.I1(CLBLM_R_X3Y106_SLICE_X2Y106_AO5),
.I2(CLBLM_R_X3Y106_SLICE_X2Y106_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(1'b1),
.I5(CLBLL_L_X2Y107_SLICE_X1Y107_BQ),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_BO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaebaaeb00500050)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_R_X3Y106_SLICE_X2Y106_AO5),
.I2(CLBLL_L_X2Y107_SLICE_X1Y107_AQ),
.I3(CLBLL_L_X2Y107_SLICE_X1Y107_DO5),
.I4(1'b1),
.I5(CLBLL_L_X2Y107_SLICE_X1Y107_BQ),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_AO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y108_SLICE_X0Y108_BO6),
.Q(CLBLL_L_X2Y108_SLICE_X0Y108_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y108_SLICE_X0Y108_AO6),
.Q(CLBLL_L_X2Y108_SLICE_X0Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y106_SLICE_X0Y106_CO6),
.Q(CLBLL_L_X2Y108_SLICE_X0Y108_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_DO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555555555555555)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_CLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_CO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0ccf0aa33335555)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_BLUT (
.I0(CLBLL_L_X2Y108_SLICE_X0Y108_A5Q),
.I1(CLBLM_R_X3Y104_SLICE_X2Y104_CO6),
.I2(CLBLL_L_X2Y108_SLICE_X0Y108_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y107_IOB_X0Y107_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_BO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc0cfc0cfc0cfc0c)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y104_SLICE_X2Y104_CO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(LIOB33_X0Y117_IOB_X0Y118_I),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_AO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_DO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_CO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_BO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_AO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y103_SLICE_X4Y103_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y103_SLICE_X4Y103_AO6),
.Q(CLBLL_L_X4Y103_SLICE_X4Y103_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8b038b03cf03cf03)
  ) CLBLL_L_X4Y103_SLICE_X4Y103_DLUT (
.I0(CLBLM_R_X5Y105_SLICE_X7Y105_AQ),
.I1(CLBLL_L_X2Y105_SLICE_X1Y105_CO6),
.I2(CLBLL_L_X4Y103_SLICE_X4Y103_AQ),
.I3(CLBLM_R_X3Y105_SLICE_X3Y105_AQ),
.I4(1'b1),
.I5(CLBLM_R_X5Y105_SLICE_X7Y105_BO6),
.O5(CLBLL_L_X4Y103_SLICE_X4Y103_DO5),
.O6(CLBLL_L_X4Y103_SLICE_X4Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff2f3fffff3f3f)
  ) CLBLL_L_X4Y103_SLICE_X4Y103_CLUT (
.I0(CLBLM_R_X3Y103_SLICE_X3Y103_BQ),
.I1(CLBLL_L_X2Y105_SLICE_X1Y105_CO6),
.I2(CLBLM_R_X5Y104_SLICE_X7Y104_BQ),
.I3(CLBLL_L_X4Y103_SLICE_X5Y103_CQ),
.I4(CLBLL_L_X4Y103_SLICE_X4Y103_DO6),
.I5(CLBLL_L_X4Y105_SLICE_X5Y105_DO6),
.O5(CLBLL_L_X4Y103_SLICE_X4Y103_CO5),
.O6(CLBLL_L_X4Y103_SLICE_X4Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff33df13ff33ff33)
  ) CLBLL_L_X4Y103_SLICE_X4Y103_BLUT (
.I0(CLBLL_L_X4Y105_SLICE_X5Y105_DO6),
.I1(CLBLL_L_X2Y105_SLICE_X1Y105_CO6),
.I2(CLBLL_L_X4Y103_SLICE_X4Y103_AQ),
.I3(CLBLM_R_X5Y104_SLICE_X6Y104_CO6),
.I4(CLBLM_R_X3Y103_SLICE_X3Y103_BQ),
.I5(CLBLL_L_X4Y103_SLICE_X5Y103_CQ),
.O5(CLBLL_L_X4Y103_SLICE_X4Y103_BO5),
.O6(CLBLL_L_X4Y103_SLICE_X4Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaebaaeb00410041)
  ) CLBLL_L_X4Y103_SLICE_X4Y103_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLL_L_X4Y103_SLICE_X5Y103_DO6),
.I2(CLBLL_L_X4Y103_SLICE_X4Y103_AQ),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y103_SLICE_X5Y103_CQ),
.O5(CLBLL_L_X4Y103_SLICE_X4Y103_AO5),
.O6(CLBLL_L_X4Y103_SLICE_X4Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y103_SLICE_X5Y103_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y103_SLICE_X5Y103_AO6),
.Q(CLBLL_L_X4Y103_SLICE_X5Y103_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y103_SLICE_X5Y103_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y103_SLICE_X5Y103_BO6),
.Q(CLBLL_L_X4Y103_SLICE_X5Y103_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y103_SLICE_X5Y103_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y103_SLICE_X5Y103_CO6),
.Q(CLBLL_L_X4Y103_SLICE_X5Y103_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff73fff3ff73fff3)
  ) CLBLL_L_X4Y103_SLICE_X5Y103_DLUT (
.I0(CLBLL_L_X4Y104_SLICE_X5Y104_DO6),
.I1(CLBLL_L_X4Y103_SLICE_X5Y103_CQ),
.I2(CLBLL_L_X2Y105_SLICE_X0Y105_CQ),
.I3(CLBLM_R_X3Y103_SLICE_X3Y103_BQ),
.I4(CLBLL_L_X4Y105_SLICE_X5Y105_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y103_SLICE_X5Y103_DO5),
.O6(CLBLL_L_X4Y103_SLICE_X5Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hee44bb11aa00aa00)
  ) CLBLL_L_X4Y103_SLICE_X5Y103_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLL_L_X4Y104_SLICE_X5Y104_CO6),
.I2(1'b1),
.I3(CLBLM_R_X3Y103_SLICE_X3Y103_BQ),
.I4(CLBLL_L_X4Y103_SLICE_X5Y103_CQ),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLL_L_X4Y103_SLICE_X5Y103_CO5),
.O6(CLBLL_L_X4Y103_SLICE_X5Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f03000f0f0cc00)
  ) CLBLL_L_X4Y103_SLICE_X5Y103_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y103_SLICE_X5Y103_BQ),
.I2(CLBLL_L_X4Y103_SLICE_X5Y103_AQ),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLL_L_X4Y104_SLICE_X4Y104_CO5),
.O5(CLBLL_L_X4Y103_SLICE_X5Y103_BO5),
.O6(CLBLL_L_X4Y103_SLICE_X5Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff02ffa0000200a0)
  ) CLBLL_L_X4Y103_SLICE_X5Y103_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLL_L_X4Y103_SLICE_X5Y103_BQ),
.I2(CLBLL_L_X4Y103_SLICE_X5Y103_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLL_L_X4Y104_SLICE_X4Y104_CO5),
.I5(CLBLL_L_X4Y105_SLICE_X5Y105_BQ),
.O5(CLBLL_L_X4Y103_SLICE_X5Y103_AO5),
.O6(CLBLL_L_X4Y103_SLICE_X5Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y104_SLICE_X4Y104_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y104_SLICE_X4Y104_AO6),
.Q(CLBLL_L_X4Y104_SLICE_X4Y104_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y104_SLICE_X4Y104_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y104_SLICE_X4Y104_BO6),
.Q(CLBLL_L_X4Y104_SLICE_X4Y104_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000070f0f0f)
  ) CLBLL_L_X4Y104_SLICE_X4Y104_DLUT (
.I0(CLBLL_L_X4Y104_SLICE_X5Y104_AQ),
.I1(CLBLL_L_X4Y104_SLICE_X4Y104_CO5),
.I2(CLBLL_L_X4Y104_SLICE_X5Y104_BO6),
.I3(CLBLM_R_X3Y104_SLICE_X2Y104_BQ),
.I4(CLBLL_L_X4Y103_SLICE_X5Y103_BQ),
.I5(CLBLL_L_X4Y105_SLICE_X4Y105_BO6),
.O5(CLBLL_L_X4Y104_SLICE_X4Y104_DO5),
.O6(CLBLL_L_X4Y104_SLICE_X4Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbff00004000f0f0)
  ) CLBLL_L_X4Y104_SLICE_X4Y104_CLUT (
.I0(CLBLL_L_X4Y103_SLICE_X4Y103_BO6),
.I1(CLBLL_L_X4Y105_SLICE_X5Y105_BQ),
.I2(CLBLL_L_X4Y104_SLICE_X4Y104_BQ),
.I3(CLBLM_R_X5Y104_SLICE_X7Y104_BQ),
.I4(CLBLL_L_X2Y105_SLICE_X0Y105_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y104_SLICE_X4Y104_CO5),
.O6(CLBLL_L_X4Y104_SLICE_X4Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf044f044f010f000)
  ) CLBLL_L_X4Y104_SLICE_X4Y104_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLL_L_X4Y104_SLICE_X4Y104_BQ),
.I2(CLBLL_L_X4Y104_SLICE_X4Y104_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_R_X3Y104_SLICE_X3Y104_BQ),
.I5(CLBLL_L_X4Y104_SLICE_X4Y104_CO6),
.O5(CLBLL_L_X4Y104_SLICE_X4Y104_BO5),
.O6(CLBLL_L_X4Y104_SLICE_X4Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff500050ff010010)
  ) CLBLL_L_X4Y104_SLICE_X4Y104_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLL_L_X4Y104_SLICE_X4Y104_BQ),
.I2(CLBLL_L_X4Y104_SLICE_X4Y104_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_R_X3Y104_SLICE_X3Y104_BQ),
.I5(CLBLL_L_X4Y104_SLICE_X4Y104_CO6),
.O5(CLBLL_L_X4Y104_SLICE_X4Y104_AO5),
.O6(CLBLL_L_X4Y104_SLICE_X4Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y104_SLICE_X5Y104_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y104_SLICE_X5Y104_AO6),
.Q(CLBLL_L_X4Y104_SLICE_X5Y104_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000055500000055)
  ) CLBLL_L_X4Y104_SLICE_X5Y104_DLUT (
.I0(CLBLL_L_X4Y105_SLICE_X4Y105_AQ),
.I1(1'b1),
.I2(CLBLM_R_X5Y105_SLICE_X7Y105_AQ),
.I3(CLBLM_R_X3Y105_SLICE_X3Y105_AQ),
.I4(CLBLL_L_X4Y105_SLICE_X5Y105_AQ),
.I5(CLBLM_R_X5Y105_SLICE_X7Y105_BO6),
.O5(CLBLL_L_X4Y104_SLICE_X5Y104_DO5),
.O6(CLBLL_L_X4Y104_SLICE_X5Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff00ef00)
  ) CLBLL_L_X4Y104_SLICE_X5Y104_CLUT (
.I0(CLBLL_L_X4Y105_SLICE_X4Y105_AQ),
.I1(CLBLM_R_X5Y104_SLICE_X6Y104_CO6),
.I2(CLBLL_L_X4Y105_SLICE_X5Y105_CQ),
.I3(CLBLL_L_X2Y105_SLICE_X0Y105_CQ),
.I4(CLBLL_L_X4Y105_SLICE_X5Y105_AQ),
.I5(CLBLM_R_X3Y103_SLICE_X3Y103_BQ),
.O5(CLBLL_L_X4Y104_SLICE_X5Y104_CO5),
.O6(CLBLL_L_X4Y104_SLICE_X5Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h01000000ffffffff)
  ) CLBLL_L_X4Y104_SLICE_X5Y104_BLUT (
.I0(CLBLL_L_X4Y105_SLICE_X5Y105_AQ),
.I1(CLBLM_R_X5Y104_SLICE_X6Y104_CO6),
.I2(CLBLL_L_X4Y105_SLICE_X4Y105_AQ),
.I3(CLBLM_R_X3Y104_SLICE_X2Y104_AQ),
.I4(CLBLL_L_X4Y105_SLICE_X5Y105_CQ),
.I5(CLBLL_L_X2Y105_SLICE_X0Y105_BQ),
.O5(CLBLL_L_X4Y104_SLICE_X5Y104_BO5),
.O6(CLBLL_L_X4Y104_SLICE_X5Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hde30cc00f000f000)
  ) CLBLL_L_X4Y104_SLICE_X5Y104_ALUT (
.I0(CLBLL_L_X4Y104_SLICE_X4Y104_CO5),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLL_L_X4Y104_SLICE_X5Y104_AQ),
.I3(CLBLL_L_X4Y103_SLICE_X5Y103_BQ),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y104_SLICE_X5Y104_AO5),
.O6(CLBLL_L_X4Y104_SLICE_X5Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y105_SLICE_X4Y105_AO6),
.Q(CLBLL_L_X4Y105_SLICE_X4Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000100)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_DLUT (
.I0(CLBLL_L_X4Y105_SLICE_X5Y105_AQ),
.I1(CLBLL_L_X4Y105_SLICE_X4Y105_AQ),
.I2(CLBLM_R_X3Y107_SLICE_X3Y107_AO5),
.I3(CLBLM_R_X3Y104_SLICE_X3Y104_CO6),
.I4(CLBLL_L_X4Y106_SLICE_X4Y106_CO6),
.I5(CLBLM_R_X5Y104_SLICE_X6Y104_CO6),
.O5(CLBLL_L_X4Y105_SLICE_X4Y105_DO5),
.O6(CLBLL_L_X4Y105_SLICE_X4Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0eeffff00eeffff)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_CLUT (
.I0(CLBLL_L_X4Y103_SLICE_X4Y103_AQ),
.I1(CLBLL_L_X4Y103_SLICE_X5Y103_DO6),
.I2(CLBLM_R_X5Y105_SLICE_X6Y105_CO6),
.I3(CLBLL_L_X2Y105_SLICE_X1Y105_CO6),
.I4(CLBLL_L_X4Y107_SLICE_X5Y107_DO6),
.I5(CLBLM_R_X3Y105_SLICE_X3Y105_AQ),
.O5(CLBLL_L_X4Y105_SLICE_X4Y105_CO5),
.O6(CLBLL_L_X4Y105_SLICE_X4Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000accce000a000a)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_BLUT (
.I0(CLBLM_R_X5Y107_SLICE_X6Y107_DQ),
.I1(CLBLM_R_X5Y105_SLICE_X7Y105_BO6),
.I2(CLBLM_R_X5Y106_SLICE_X6Y106_AO6),
.I3(CLBLL_L_X2Y105_SLICE_X0Y105_DQ),
.I4(CLBLM_R_X5Y105_SLICE_X7Y105_AQ),
.I5(CLBLM_R_X3Y105_SLICE_X2Y105_BQ),
.O5(CLBLL_L_X4Y105_SLICE_X4Y105_BO5),
.O6(CLBLL_L_X4Y105_SLICE_X4Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000030033003)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(CLBLL_L_X4Y105_SLICE_X4Y105_AQ),
.I3(CLBLM_R_X5Y104_SLICE_X6Y104_CO6),
.I4(CLBLL_L_X4Y103_SLICE_X4Y103_AQ),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLL_L_X4Y105_SLICE_X4Y105_AO5),
.O6(CLBLL_L_X4Y105_SLICE_X4Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y105_SLICE_X5Y105_AO6),
.Q(CLBLL_L_X4Y105_SLICE_X5Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y105_SLICE_X5Y105_BO6),
.Q(CLBLL_L_X4Y105_SLICE_X5Y105_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y105_SLICE_X5Y105_CO6),
.Q(CLBLL_L_X4Y105_SLICE_X5Y105_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff04ff00ff44ff)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_DLUT (
.I0(CLBLL_L_X4Y105_SLICE_X4Y105_AQ),
.I1(CLBLL_L_X4Y105_SLICE_X5Y105_CQ),
.I2(CLBLM_R_X3Y105_SLICE_X3Y105_AQ),
.I3(CLBLL_L_X2Y105_SLICE_X0Y105_CQ),
.I4(CLBLL_L_X4Y105_SLICE_X5Y105_AQ),
.I5(CLBLM_R_X5Y105_SLICE_X7Y105_CO6),
.O5(CLBLL_L_X4Y105_SLICE_X5Y105_DO5),
.O6(CLBLL_L_X4Y105_SLICE_X5Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000044444441)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLL_L_X4Y105_SLICE_X5Y105_CQ),
.I2(CLBLM_R_X5Y104_SLICE_X6Y104_CO6),
.I3(CLBLL_L_X4Y105_SLICE_X4Y105_AQ),
.I4(CLBLL_L_X4Y105_SLICE_X5Y105_AQ),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLL_L_X4Y105_SLICE_X5Y105_CO5),
.O6(CLBLL_L_X4Y105_SLICE_X5Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00c3cc0000)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y105_SLICE_X5Y105_BQ),
.I2(CLBLL_L_X4Y103_SLICE_X4Y103_BO6),
.I3(CLBLM_R_X5Y104_SLICE_X7Y104_BQ),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLL_L_X4Y105_SLICE_X5Y105_BO5),
.O6(CLBLL_L_X4Y105_SLICE_X5Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0fa0009f0fa0009)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_ALUT (
.I0(CLBLL_L_X4Y105_SLICE_X5Y105_AQ),
.I1(CLBLM_R_X5Y104_SLICE_X6Y104_CO6),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(CLBLL_L_X4Y105_SLICE_X4Y105_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y105_SLICE_X5Y105_AO5),
.O6(CLBLL_L_X4Y105_SLICE_X5Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y106_SLICE_X4Y106_BO5),
.Q(CLBLL_L_X4Y106_SLICE_X4Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc8c8c8c8c8fec8c8)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_DLUT (
.I0(CLBLL_L_X4Y106_SLICE_X4Y106_CO5),
.I1(CLBLL_L_X4Y106_SLICE_X4Y106_AQ),
.I2(CLBLL_L_X2Y106_SLICE_X1Y106_DO6),
.I3(CLBLL_L_X4Y106_SLICE_X4Y106_AO5),
.I4(CLBLL_L_X4Y106_SLICE_X5Y106_AQ),
.I5(CLBLM_R_X3Y106_SLICE_X2Y106_DO6),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_DO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdfdfccdf0f0f000f)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_CLUT (
.I0(CLBLL_L_X2Y106_SLICE_X0Y106_AO6),
.I1(CLBLL_L_X4Y106_SLICE_X4Y106_AQ),
.I2(CLBLM_R_X3Y106_SLICE_X2Y106_AQ),
.I3(CLBLL_L_X2Y105_SLICE_X0Y105_BQ),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_CO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0fffffffcddc1010)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_BLUT (
.I0(CLBLM_R_X3Y106_SLICE_X2Y106_CO5),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLL_L_X4Y106_SLICE_X4Y106_AQ),
.I3(CLBLM_R_X3Y104_SLICE_X2Y104_DO6),
.I4(CLBLL_L_X4Y106_SLICE_X5Y106_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_BO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0bbbf44444444444)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_ALUT (
.I0(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I1(CLBLL_L_X2Y105_SLICE_X0Y105_BQ),
.I2(CLBLM_R_X3Y106_SLICE_X2Y106_BQ),
.I3(CLBLL_L_X2Y106_SLICE_X0Y106_AO6),
.I4(CLBLL_L_X4Y106_SLICE_X5Y106_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_AO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y106_SLICE_X5Y106_AO6),
.Q(CLBLL_L_X4Y106_SLICE_X5Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_DO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_CO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_BO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3c003c003c00)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y104_SLICE_X2Y104_DO6),
.I2(CLBLL_L_X4Y106_SLICE_X5Y106_AQ),
.I3(CLBLM_R_X3Y106_SLICE_X2Y106_CO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLL_L_X4Y105_SLICE_X5Y105_CQ),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_AO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y107_SLICE_X4Y107_AO6),
.Q(CLBLL_L_X4Y107_SLICE_X4Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y107_SLICE_X4Y107_BO6),
.Q(CLBLL_L_X4Y107_SLICE_X4Y107_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y107_SLICE_X4Y107_CO6),
.Q(CLBLL_L_X4Y107_SLICE_X4Y107_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6fffff6ff6fffff6)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_DLUT (
.I0(CLBLL_L_X4Y107_SLICE_X5Y107_AQ),
.I1(CLBLM_R_X3Y106_SLICE_X2Y106_BQ),
.I2(CLBLL_L_X2Y107_SLICE_X1Y107_AQ),
.I3(CLBLM_R_X3Y106_SLICE_X2Y106_AQ),
.I4(CLBLL_L_X4Y107_SLICE_X5Y107_BQ),
.I5(CLBLM_R_X3Y107_SLICE_X2Y107_AQ),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_DO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc9cfcccf000f000)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_CLUT (
.I0(CLBLL_L_X4Y106_SLICE_X4Y106_BO6),
.I1(CLBLL_L_X4Y107_SLICE_X4Y107_CQ),
.I2(CLBLL_L_X4Y107_SLICE_X4Y107_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLL_L_X4Y107_SLICE_X4Y107_BQ),
.I5(CLBLM_R_X3Y106_SLICE_X2Y106_CO6),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_CO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heca0b3a0eca0b3a0)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_BLUT (
.I0(CLBLL_L_X4Y106_SLICE_X4Y106_AQ),
.I1(CLBLL_L_X4Y107_SLICE_X4Y107_BQ),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_R_X3Y106_SLICE_X2Y106_CO6),
.I4(CLBLL_L_X4Y106_SLICE_X4Y106_BO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_BO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc0acc06cc0acc06)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_ALUT (
.I0(CLBLL_L_X4Y107_SLICE_X4Y107_AQ),
.I1(CLBLL_L_X4Y107_SLICE_X4Y107_BQ),
.I2(CLBLM_R_X3Y106_SLICE_X2Y106_CO5),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLL_L_X4Y106_SLICE_X4Y106_BO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_AO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y107_SLICE_X5Y107_AO6),
.Q(CLBLL_L_X4Y107_SLICE_X5Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y107_SLICE_X5Y107_BO6),
.Q(CLBLL_L_X4Y107_SLICE_X5Y107_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff0fff0fff0fff0)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X4Y107_SLICE_X4Y107_DO6),
.I3(CLBLL_L_X4Y107_SLICE_X5Y107_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_DO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaffffaaaaffffa9)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_CLUT (
.I0(CLBLL_L_X2Y107_SLICE_X1Y107_CQ),
.I1(CLBLM_R_X3Y107_SLICE_X2Y107_AQ),
.I2(CLBLL_L_X4Y107_SLICE_X5Y107_BQ),
.I3(CLBLM_R_X3Y107_SLICE_X2Y107_BQ),
.I4(CLBLL_L_X2Y107_SLICE_X1Y107_BQ),
.I5(CLBLL_L_X4Y107_SLICE_X5Y107_AQ),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_CO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeeefcccfaaaf000)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_BLUT (
.I0(CLBLL_L_X2Y107_SLICE_X0Y107_DO6),
.I1(CLBLL_L_X2Y107_SLICE_X0Y107_DO5),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLL_L_X4Y107_SLICE_X5Y107_AQ),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(CLBLL_L_X4Y107_SLICE_X5Y107_BQ),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_BO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefafcf0eeaacc00)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_ALUT (
.I0(CLBLL_L_X2Y107_SLICE_X0Y107_DO6),
.I1(CLBLL_L_X2Y107_SLICE_X0Y107_DO5),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLL_L_X4Y107_SLICE_X5Y107_AQ),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(CLBLL_L_X2Y107_SLICE_X1Y107_CQ),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_AO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y103_SLICE_X2Y103_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y103_SLICE_X2Y103_AO6),
.Q(CLBLM_R_X3Y103_SLICE_X2Y103_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y103_SLICE_X2Y103_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y103_SLICE_X2Y103_BO6),
.Q(CLBLM_R_X3Y103_SLICE_X2Y103_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y103_SLICE_X2Y103_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y103_SLICE_X2Y103_CO6),
.Q(CLBLM_R_X3Y103_SLICE_X2Y103_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y103_SLICE_X2Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y103_SLICE_X2Y103_DO5),
.O6(CLBLM_R_X3Y103_SLICE_X2Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa3000c000)
  ) CLBLM_R_X3Y103_SLICE_X2Y103_CLUT (
.I0(CLBLL_L_X2Y105_SLICE_X0Y105_AQ),
.I1(CLBLM_R_X3Y103_SLICE_X3Y103_CO6),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLL_L_X2Y103_SLICE_X1Y103_CO6),
.I4(CLBLM_R_X3Y103_SLICE_X2Y103_CQ),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X3Y103_SLICE_X2Y103_CO5),
.O6(CLBLM_R_X3Y103_SLICE_X2Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf030f088f0f0f000)
  ) CLBLM_R_X3Y103_SLICE_X2Y103_BLUT (
.I0(CLBLM_R_X3Y103_SLICE_X2Y103_BQ),
.I1(CLBLM_R_X5Y103_SLICE_X7Y103_AO6),
.I2(CLBLM_R_X3Y103_SLICE_X2Y103_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLL_L_X2Y105_SLICE_X0Y105_CQ),
.O5(CLBLM_R_X3Y103_SLICE_X2Y103_BO5),
.O6(CLBLM_R_X3Y103_SLICE_X2Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff620040ffaa0000)
  ) CLBLM_R_X3Y103_SLICE_X2Y103_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X5Y103_SLICE_X7Y103_AO6),
.I2(CLBLM_R_X3Y103_SLICE_X2Y103_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_R_X3Y103_SLICE_X3Y103_AQ),
.I5(CLBLL_L_X2Y105_SLICE_X0Y105_CQ),
.O5(CLBLM_R_X3Y103_SLICE_X2Y103_AO5),
.O6(CLBLM_R_X3Y103_SLICE_X2Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y103_SLICE_X3Y103_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y103_SLICE_X3Y103_AO6),
.Q(CLBLM_R_X3Y103_SLICE_X3Y103_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y103_SLICE_X3Y103_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y103_SLICE_X3Y103_BO6),
.Q(CLBLM_R_X3Y103_SLICE_X3Y103_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0cfc0cf55555555)
  ) CLBLM_R_X3Y103_SLICE_X3Y103_DLUT (
.I0(CLBLL_L_X4Y103_SLICE_X4Y103_AQ),
.I1(CLBLM_R_X5Y105_SLICE_X7Y105_AQ),
.I2(CLBLM_R_X3Y105_SLICE_X3Y105_AQ),
.I3(CLBLM_R_X3Y105_SLICE_X2Y105_A5Q),
.I4(1'b1),
.I5(CLBLL_L_X2Y105_SLICE_X1Y105_CO6),
.O5(CLBLM_R_X3Y103_SLICE_X3Y103_DO5),
.O6(CLBLM_R_X3Y103_SLICE_X3Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcecccececccccece)
  ) CLBLM_R_X3Y103_SLICE_X3Y103_CLUT (
.I0(CLBLL_L_X4Y105_SLICE_X5Y105_BQ),
.I1(CLBLL_L_X2Y105_SLICE_X0Y105_BQ),
.I2(CLBLL_L_X4Y103_SLICE_X4Y103_CO6),
.I3(CLBLL_L_X4Y104_SLICE_X5Y104_AO5),
.I4(CLBLL_L_X2Y105_SLICE_X0Y105_CQ),
.I5(CLBLL_L_X4Y104_SLICE_X4Y104_BQ),
.O5(CLBLM_R_X3Y103_SLICE_X3Y103_CO5),
.O6(CLBLM_R_X3Y103_SLICE_X3Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff6600000066)
  ) CLBLM_R_X3Y103_SLICE_X3Y103_BLUT (
.I0(CLBLL_L_X4Y105_SLICE_X5Y105_DO6),
.I1(CLBLM_R_X3Y103_SLICE_X3Y103_BQ),
.I2(1'b1),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLM_R_X3Y105_SLICE_X2Y105_A5Q),
.O5(CLBLM_R_X3Y103_SLICE_X3Y103_BO5),
.O6(CLBLM_R_X3Y103_SLICE_X3Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc50888888)
  ) CLBLM_R_X3Y103_SLICE_X3Y103_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X3Y104_SLICE_X3Y104_AQ),
.I2(CLBLM_R_X3Y103_SLICE_X3Y103_AQ),
.I3(CLBLL_L_X2Y105_SLICE_X0Y105_CQ),
.I4(CLBLM_R_X5Y103_SLICE_X7Y103_AO6),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X3Y103_SLICE_X3Y103_AO5),
.O6(CLBLM_R_X3Y103_SLICE_X3Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y104_SLICE_X2Y104_AO6),
.Q(CLBLM_R_X3Y104_SLICE_X2Y104_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y104_SLICE_X2Y104_BO6),
.Q(CLBLM_R_X3Y104_SLICE_X2Y104_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8800000000000000)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_DLUT (
.I0(CLBLM_R_X3Y104_SLICE_X3Y104_AQ),
.I1(CLBLM_R_X3Y103_SLICE_X2Y103_AQ),
.I2(1'b1),
.I3(CLBLL_L_X2Y108_SLICE_X0Y108_BO5),
.I4(CLBLM_R_X3Y103_SLICE_X3Y103_AQ),
.I5(CLBLM_R_X3Y103_SLICE_X2Y103_BQ),
.O5(CLBLM_R_X3Y104_SLICE_X2Y104_DO5),
.O6(CLBLM_R_X3Y104_SLICE_X2Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0f8f0f0e0)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_CLUT (
.I0(CLBLM_R_X3Y104_SLICE_X3Y104_AQ),
.I1(CLBLM_R_X3Y103_SLICE_X2Y103_AQ),
.I2(CLBLL_L_X2Y108_SLICE_X0Y108_AQ),
.I3(CLBLM_R_X3Y103_SLICE_X2Y103_BQ),
.I4(CLBLM_R_X3Y103_SLICE_X3Y103_AQ),
.I5(LIOB33_X0Y107_IOB_X0Y107_I),
.O5(CLBLM_R_X3Y104_SLICE_X2Y104_CO5),
.O6(CLBLM_R_X3Y104_SLICE_X2Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0a0a04444)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X3Y104_SLICE_X2Y104_BQ),
.I2(CLBLM_R_X3Y104_SLICE_X2Y104_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X3Y104_SLICE_X2Y104_BO5),
.O6(CLBLM_R_X3Y104_SLICE_X2Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee00dc10ee00dc10)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_R_X3Y104_SLICE_X2Y104_AQ),
.I3(CLBLM_R_X3Y105_SLICE_X2Y105_BQ),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y104_SLICE_X2Y104_AO5),
.O6(CLBLM_R_X3Y104_SLICE_X2Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y104_SLICE_X3Y104_AO6),
.Q(CLBLM_R_X3Y104_SLICE_X3Y104_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y104_SLICE_X3Y104_BO6),
.Q(CLBLM_R_X3Y104_SLICE_X3Y104_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y104_SLICE_X3Y104_DO5),
.O6(CLBLM_R_X3Y104_SLICE_X3Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000800000000000)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_CLUT (
.I0(CLBLM_R_X3Y104_SLICE_X2Y104_AQ),
.I1(CLBLL_L_X2Y105_SLICE_X0Y105_BQ),
.I2(CLBLL_L_X2Y104_SLICE_X0Y104_AQ),
.I3(CLBLL_L_X4Y105_SLICE_X5Y105_CQ),
.I4(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I5(LIOB33_X0Y103_IOB_X0Y104_I),
.O5(CLBLM_R_X3Y104_SLICE_X3Y104_CO5),
.O6(CLBLM_R_X3Y104_SLICE_X3Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f04400f0f04411)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X3Y104_SLICE_X3Y104_BQ),
.I2(CLBLM_R_X3Y103_SLICE_X2Y103_BQ),
.I3(CLBLL_L_X4Y104_SLICE_X4Y104_CO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLL_L_X4Y104_SLICE_X4Y104_BQ),
.O5(CLBLM_R_X3Y104_SLICE_X3Y104_BO5),
.O6(CLBLM_R_X3Y104_SLICE_X3Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaacc00aaaa3030)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_ALUT (
.I0(CLBLL_L_X4Y107_SLICE_X4Y107_CQ),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(CLBLM_R_X3Y104_SLICE_X3Y104_AQ),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_R_X5Y104_SLICE_X7Y104_CO6),
.O5(CLBLM_R_X3Y104_SLICE_X3Y104_AO5),
.O6(CLBLM_R_X3Y104_SLICE_X3Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y105_SLICE_X2Y105_CO5),
.Q(CLBLM_R_X3Y105_SLICE_X2Y105_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y105_SLICE_X2Y105_DO5),
.Q(CLBLM_R_X3Y105_SLICE_X2Y105_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y105_SLICE_X2Y105_AO6),
.Q(CLBLM_R_X3Y105_SLICE_X2Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y105_SLICE_X2Y105_BO6),
.Q(CLBLM_R_X3Y105_SLICE_X2Y105_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a0fc0cf000)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_DLUT (
.I0(CLBLM_R_X3Y107_SLICE_X2Y107_AQ),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLL_L_X2Y107_SLICE_X0Y107_CQ),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y105_SLICE_X2Y105_DO5),
.O6(CLBLM_R_X3Y105_SLICE_X2Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h11113333c0c0c0f3)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y105_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_R_X5Y105_SLICE_X7Y105_AQ),
.I3(CLBLM_R_X3Y105_SLICE_X2Y105_A5Q),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y105_SLICE_X2Y105_CO5),
.O6(CLBLM_R_X3Y105_SLICE_X2Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000004a404a4)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_BLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X3Y105_SLICE_X2Y105_BQ),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(CLBLL_L_X2Y105_SLICE_X0Y105_DQ),
.I4(CLBLM_R_X3Y105_SLICE_X2Y105_B5Q),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X3Y105_SLICE_X2Y105_BO5),
.O6(CLBLM_R_X3Y105_SLICE_X2Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfabaaaaaffffaaaa)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_ALUT (
.I0(CLBLM_R_X3Y105_SLICE_X2Y105_DO6),
.I1(CLBLL_L_X2Y104_SLICE_X1Y104_BO6),
.I2(CLBLM_R_X3Y105_SLICE_X2Y105_AQ),
.I3(CLBLL_L_X4Y107_SLICE_X5Y107_DO6),
.I4(CLBLL_L_X2Y107_SLICE_X1Y107_DO6),
.I5(CLBLL_L_X4Y105_SLICE_X4Y105_CO6),
.O5(CLBLM_R_X3Y105_SLICE_X2Y105_AO5),
.O6(CLBLM_R_X3Y105_SLICE_X2Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y105_SLICE_X3Y105_AO6),
.Q(CLBLM_R_X3Y105_SLICE_X3Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y105_SLICE_X3Y105_DO5),
.O6(CLBLM_R_X3Y105_SLICE_X3Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccfc0030cccc0000)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_CLUT (
.I0(1'b1),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLL_L_X2Y105_SLICE_X0Y105_BQ),
.I4(CLBLM_R_X3Y105_SLICE_X3Y105_AQ),
.I5(CLBLM_R_X3Y105_SLICE_X3Y105_BO6),
.O5(CLBLM_R_X3Y105_SLICE_X3Y105_CO5),
.O6(CLBLM_R_X3Y105_SLICE_X3Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcf4cc44f8f08800)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_BLUT (
.I0(CLBLL_L_X2Y105_SLICE_X0Y105_CQ),
.I1(CLBLL_L_X2Y105_SLICE_X1Y105_CO6),
.I2(CLBLM_R_X3Y105_SLICE_X2Y105_A5Q),
.I3(CLBLL_L_X4Y104_SLICE_X5Y104_AQ),
.I4(LIOB33_X0Y113_IOB_X0Y113_I),
.I5(CLBLL_L_X4Y105_SLICE_X5Y105_BQ),
.O5(CLBLM_R_X3Y105_SLICE_X3Y105_BO5),
.O6(CLBLM_R_X3Y105_SLICE_X3Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaf8fbf8faf8f8f8)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_ALUT (
.I0(CLBLL_L_X2Y105_SLICE_X0Y105_CQ),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_R_X3Y105_SLICE_X2Y105_CO6),
.I3(CLBLM_R_X3Y105_SLICE_X2Y105_B5Q),
.I4(LIOB33_X0Y101_IOB_X0Y102_I),
.I5(CLBLM_R_X3Y105_SLICE_X3Y105_AQ),
.O5(CLBLM_R_X3Y105_SLICE_X3Y105_AO5),
.O6(CLBLM_R_X3Y105_SLICE_X3Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y106_SLICE_X2Y106_AO6),
.Q(CLBLM_R_X3Y106_SLICE_X2Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y106_SLICE_X2Y106_BO6),
.Q(CLBLM_R_X3Y106_SLICE_X2Y106_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000a8a80000aa00)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_DLUT (
.I0(CLBLM_R_X3Y106_SLICE_X2Y106_BQ),
.I1(CLBLL_L_X2Y107_SLICE_X0Y107_CQ),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(CLBLL_L_X2Y107_SLICE_X0Y107_BQ),
.I4(CLBLL_L_X2Y105_SLICE_X0Y105_BQ),
.I5(CLBLL_L_X2Y106_SLICE_X1Y106_AQ),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_DO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4444544433330333)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_CLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLL_L_X2Y105_SLICE_X0Y105_BQ),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLL_L_X2Y103_SLICE_X1Y103_CO6),
.I4(LIOB33_X0Y113_IOB_X0Y114_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_CO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8f28822f8f28822)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_BLUT (
.I0(CLBLL_L_X2Y107_SLICE_X1Y107_DO6),
.I1(CLBLM_R_X3Y106_SLICE_X2Y106_BQ),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLL_L_X4Y105_SLICE_X4Y105_CO6),
.I4(CLBLL_L_X2Y104_SLICE_X0Y104_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_BO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdccd1010ff0fffff)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_ALUT (
.I0(CLBLL_L_X2Y107_SLICE_X1Y107_DO5),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_R_X3Y106_SLICE_X2Y106_AQ),
.I3(CLBLL_L_X4Y105_SLICE_X4Y105_CO6),
.I4(CLBLM_R_X3Y106_SLICE_X2Y106_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_AO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff00000a2a)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_DLUT (
.I0(CLBLM_R_X3Y106_SLICE_X3Y106_AO6),
.I1(CLBLM_R_X3Y107_SLICE_X3Y107_AO6),
.I2(CLBLM_R_X3Y107_SLICE_X3Y107_AO5),
.I3(CLBLL_L_X4Y106_SLICE_X4Y106_DO6),
.I4(CLBLM_R_X3Y107_SLICE_X3Y107_BO6),
.I5(CLBLM_R_X3Y107_SLICE_X3Y107_DO6),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_DO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffff7f3f)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_CLUT (
.I0(CLBLL_L_X4Y107_SLICE_X4Y107_AQ),
.I1(CLBLL_L_X4Y106_SLICE_X4Y106_CO6),
.I2(CLBLM_R_X3Y107_SLICE_X3Y107_AO5),
.I3(CLBLM_R_X3Y106_SLICE_X3Y106_AO5),
.I4(CLBLM_R_X3Y107_SLICE_X3Y107_BO6),
.I5(CLBLL_L_X4Y106_SLICE_X4Y106_AO6),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_CO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff00e0ffff00ff)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_BLUT (
.I0(CLBLL_L_X4Y106_SLICE_X4Y106_DO6),
.I1(CLBLM_R_X3Y107_SLICE_X3Y107_AO6),
.I2(CLBLM_R_X3Y107_SLICE_X3Y107_AO5),
.I3(CLBLM_R_X3Y107_SLICE_X3Y107_DO6),
.I4(CLBLL_L_X2Y108_SLICE_X0Y108_BQ),
.I5(CLBLM_R_X3Y107_SLICE_X3Y107_CO6),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_BO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf4ff44fff4f44444)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_ALUT (
.I0(LIOB33_X0Y109_IOB_X0Y110_I),
.I1(CLBLL_L_X2Y105_SLICE_X0Y105_BQ),
.I2(CLBLL_L_X2Y107_SLICE_X1Y107_AQ),
.I3(CLBLL_L_X4Y107_SLICE_X4Y107_AQ),
.I4(CLBLL_L_X2Y106_SLICE_X0Y106_AO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_AO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y107_SLICE_X2Y107_AO6),
.Q(CLBLM_R_X3Y107_SLICE_X2Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y107_SLICE_X2Y107_BO6),
.Q(CLBLM_R_X3Y107_SLICE_X2Y107_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000fcaa0000)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_DLUT (
.I0(CLBLL_L_X2Y107_SLICE_X0Y107_BQ),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(CLBLL_L_X2Y107_SLICE_X0Y107_CQ),
.I3(CLBLL_L_X2Y106_SLICE_X1Y106_AQ),
.I4(CLBLL_L_X2Y107_SLICE_X1Y107_AQ),
.I5(CLBLL_L_X2Y105_SLICE_X0Y105_BQ),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_DO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff0355ffff)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_CLUT (
.I0(CLBLL_L_X2Y107_SLICE_X0Y107_BQ),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(CLBLL_L_X2Y107_SLICE_X0Y107_CQ),
.I3(CLBLL_L_X2Y106_SLICE_X1Y106_AQ),
.I4(CLBLL_L_X2Y107_SLICE_X1Y107_CQ),
.I5(CLBLL_L_X2Y105_SLICE_X0Y105_BQ),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_CO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff8f8f8ff888888)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_BLUT (
.I0(CLBLL_L_X2Y107_SLICE_X0Y107_DO5),
.I1(CLBLM_R_X3Y107_SLICE_X2Y107_BQ),
.I2(LIOB33_X0Y115_IOB_X0Y115_I),
.I3(CLBLL_L_X4Y107_SLICE_X5Y107_BQ),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLL_L_X2Y107_SLICE_X0Y107_DO6),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_BO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeca0eca0eca0)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_ALUT (
.I0(CLBLL_L_X2Y107_SLICE_X0Y107_DO5),
.I1(CLBLM_R_X3Y107_SLICE_X2Y107_BQ),
.I2(CLBLM_R_X3Y107_SLICE_X2Y107_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLL_L_X2Y107_SLICE_X0Y107_DO6),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_AO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h117755ff107350ff)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_DLUT (
.I0(CLBLL_L_X4Y107_SLICE_X4Y107_AQ),
.I1(CLBLM_R_X3Y107_SLICE_X2Y107_CO6),
.I2(CLBLM_R_X3Y107_SLICE_X2Y107_DO6),
.I3(CLBLL_L_X4Y107_SLICE_X4Y107_CQ),
.I4(CLBLM_R_X3Y107_SLICE_X3Y107_BO5),
.I5(CLBLL_L_X2Y107_SLICE_X0Y107_AO6),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_DO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3c3cf0f03c14f050)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_CLUT (
.I0(CLBLL_L_X4Y107_SLICE_X4Y107_AQ),
.I1(CLBLM_R_X3Y107_SLICE_X2Y107_CO6),
.I2(CLBLL_L_X4Y107_SLICE_X4Y107_CQ),
.I3(CLBLM_R_X3Y107_SLICE_X2Y107_DO6),
.I4(CLBLM_R_X3Y107_SLICE_X3Y107_BO5),
.I5(CLBLL_L_X2Y107_SLICE_X0Y107_AO6),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_CO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5aaa5666ffff3333)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_BLUT (
.I0(CLBLL_L_X4Y107_SLICE_X4Y107_CQ),
.I1(CLBLL_L_X2Y105_SLICE_X0Y105_BQ),
.I2(CLBLL_L_X2Y106_SLICE_X0Y106_AO6),
.I3(CLBLL_L_X2Y107_SLICE_X1Y107_CQ),
.I4(LIOB33_X0Y111_IOB_X0Y111_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_BO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5f001300ff5fff13)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_ALUT (
.I0(CLBLL_L_X2Y107_SLICE_X1Y107_BQ),
.I1(CLBLL_L_X2Y105_SLICE_X0Y105_BQ),
.I2(CLBLL_L_X2Y106_SLICE_X0Y106_AO6),
.I3(CLBLL_L_X4Y107_SLICE_X4Y107_BQ),
.I4(LIOB33_X0Y109_IOB_X0Y109_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_AO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y103_SLICE_X6Y103_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y103_SLICE_X6Y103_AO6),
.Q(CLBLM_R_X5Y103_SLICE_X6Y103_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y103_SLICE_X6Y103_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y103_SLICE_X6Y103_BO6),
.Q(CLBLM_R_X5Y103_SLICE_X6Y103_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y103_SLICE_X6Y103_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y103_SLICE_X6Y103_CO6),
.Q(CLBLM_R_X5Y103_SLICE_X6Y103_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4040c0c00000c0c0)
  ) CLBLM_R_X5Y103_SLICE_X6Y103_DLUT (
.I0(CLBLM_R_X5Y105_SLICE_X7Y105_AQ),
.I1(CLBLM_R_X5Y103_SLICE_X6Y103_CQ),
.I2(CLBLM_R_X5Y103_SLICE_X6Y103_AQ),
.I3(1'b1),
.I4(CLBLM_R_X3Y105_SLICE_X3Y105_AQ),
.I5(CLBLM_R_X5Y105_SLICE_X7Y105_BO6),
.O5(CLBLM_R_X5Y103_SLICE_X6Y103_DO5),
.O6(CLBLM_R_X5Y103_SLICE_X6Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf8f8f2f208080202)
  ) CLBLM_R_X5Y103_SLICE_X6Y103_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X5Y103_SLICE_X6Y103_CQ),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(1'b1),
.I4(CLBLM_R_X5Y104_SLICE_X6Y104_CO6),
.I5(CLBLL_L_X4Y104_SLICE_X4Y104_BQ),
.O5(CLBLM_R_X5Y103_SLICE_X6Y103_CO5),
.O6(CLBLM_R_X5Y103_SLICE_X6Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cc640000)
  ) CLBLM_R_X5Y103_SLICE_X6Y103_BLUT (
.I0(CLBLM_R_X5Y103_SLICE_X6Y103_CQ),
.I1(CLBLM_R_X5Y103_SLICE_X6Y103_BQ),
.I2(CLBLM_R_X5Y103_SLICE_X6Y103_AQ),
.I3(CLBLM_R_X5Y104_SLICE_X6Y104_CO6),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X5Y103_SLICE_X6Y103_BO5),
.O6(CLBLM_R_X5Y103_SLICE_X6Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaf0520000)
  ) CLBLM_R_X5Y103_SLICE_X6Y103_ALUT (
.I0(CLBLM_R_X5Y103_SLICE_X6Y103_CQ),
.I1(CLBLM_R_X5Y103_SLICE_X6Y103_BQ),
.I2(CLBLM_R_X5Y103_SLICE_X6Y103_AQ),
.I3(CLBLM_R_X5Y104_SLICE_X6Y104_CO6),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X5Y103_SLICE_X6Y103_AO5),
.O6(CLBLM_R_X5Y103_SLICE_X6Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y103_SLICE_X7Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y103_SLICE_X7Y103_DO5),
.O6(CLBLM_R_X5Y103_SLICE_X7Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y103_SLICE_X7Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y103_SLICE_X7Y103_CO5),
.O6(CLBLM_R_X5Y103_SLICE_X7Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y103_SLICE_X7Y103_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y103_SLICE_X7Y103_BO5),
.O6(CLBLM_R_X5Y103_SLICE_X7Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaff22ffffffffff)
  ) CLBLM_R_X5Y103_SLICE_X7Y103_ALUT (
.I0(CLBLM_R_X3Y105_SLICE_X3Y105_AQ),
.I1(CLBLM_R_X5Y105_SLICE_X7Y105_BO6),
.I2(1'b1),
.I3(CLBLM_R_X5Y103_SLICE_X6Y103_BQ),
.I4(CLBLM_R_X5Y105_SLICE_X7Y105_AQ),
.I5(CLBLM_R_X5Y103_SLICE_X6Y103_CQ),
.O5(CLBLM_R_X5Y103_SLICE_X7Y103_AO5),
.O6(CLBLM_R_X5Y103_SLICE_X7Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y104_SLICE_X6Y104_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y104_SLICE_X6Y104_AO6),
.Q(CLBLM_R_X5Y104_SLICE_X6Y104_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y104_SLICE_X6Y104_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y104_SLICE_X6Y104_BO6),
.Q(CLBLM_R_X5Y104_SLICE_X6Y104_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h1000000000000000)
  ) CLBLM_R_X5Y104_SLICE_X6Y104_DLUT (
.I0(CLBLL_L_X4Y103_SLICE_X5Y103_DO6),
.I1(CLBLL_L_X4Y103_SLICE_X4Y103_BO6),
.I2(CLBLM_R_X5Y104_SLICE_X7Y104_DO6),
.I3(CLBLM_R_X5Y103_SLICE_X6Y103_DO6),
.I4(CLBLL_L_X4Y105_SLICE_X4Y105_DO6),
.I5(CLBLM_R_X5Y104_SLICE_X7Y104_BQ),
.O5(CLBLM_R_X5Y104_SLICE_X6Y104_DO5),
.O6(CLBLM_R_X5Y104_SLICE_X6Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffdf0000ffff0000)
  ) CLBLM_R_X5Y104_SLICE_X6Y104_CLUT (
.I0(CLBLM_R_X5Y104_SLICE_X6Y104_BQ),
.I1(CLBLM_R_X5Y106_SLICE_X6Y106_CO6),
.I2(CLBLM_R_X5Y104_SLICE_X6Y104_AQ),
.I3(CLBLM_R_X5Y105_SLICE_X7Y105_AQ),
.I4(CLBLM_R_X3Y105_SLICE_X3Y105_AQ),
.I5(CLBLM_R_X5Y105_SLICE_X6Y105_BQ),
.O5(CLBLM_R_X5Y104_SLICE_X6Y104_CO5),
.O6(CLBLM_R_X5Y104_SLICE_X6Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f09ccc0000)
  ) CLBLM_R_X5Y104_SLICE_X6Y104_BLUT (
.I0(CLBLM_R_X5Y106_SLICE_X6Y106_CO6),
.I1(CLBLM_R_X5Y104_SLICE_X6Y104_BQ),
.I2(CLBLM_R_X5Y104_SLICE_X6Y104_AQ),
.I3(CLBLM_R_X5Y105_SLICE_X6Y105_BQ),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X5Y104_SLICE_X6Y104_BO5),
.O6(CLBLM_R_X5Y104_SLICE_X6Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccf0cc00cc3ccc00)
  ) CLBLM_R_X5Y104_SLICE_X6Y104_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y105_SLICE_X6Y105_BQ),
.I2(CLBLM_R_X5Y104_SLICE_X6Y104_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLM_R_X5Y106_SLICE_X6Y106_CO6),
.O5(CLBLM_R_X5Y104_SLICE_X6Y104_AO5),
.O6(CLBLM_R_X5Y104_SLICE_X6Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y104_SLICE_X7Y104_AO6),
.Q(CLBLM_R_X5Y104_SLICE_X7Y104_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y104_SLICE_X7Y104_BO6),
.Q(CLBLM_R_X5Y104_SLICE_X7Y104_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c8c8c8c0c0c0c0c)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_DLUT (
.I0(CLBLM_R_X5Y103_SLICE_X6Y103_CQ),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(CLBLL_L_X2Y105_SLICE_X0Y105_CQ),
.I3(CLBLM_R_X5Y105_SLICE_X7Y105_CO6),
.I4(CLBLM_R_X3Y105_SLICE_X3Y105_AQ),
.I5(CLBLM_R_X5Y103_SLICE_X6Y103_BQ),
.O5(CLBLM_R_X5Y104_SLICE_X7Y104_DO5),
.O6(CLBLM_R_X5Y104_SLICE_X7Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h2f0fafaf0f0f0f0f)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_CLUT (
.I0(CLBLM_R_X5Y103_SLICE_X6Y103_CQ),
.I1(CLBLM_R_X5Y105_SLICE_X7Y105_AQ),
.I2(CLBLL_L_X2Y105_SLICE_X0Y105_CQ),
.I3(CLBLM_R_X5Y105_SLICE_X7Y105_BO6),
.I4(CLBLM_R_X3Y105_SLICE_X3Y105_AQ),
.I5(CLBLM_R_X5Y103_SLICE_X6Y103_BQ),
.O5(CLBLM_R_X5Y104_SLICE_X7Y104_CO5),
.O6(CLBLM_R_X5Y104_SLICE_X7Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf098f000f098f000)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_BLUT (
.I0(CLBLL_L_X4Y103_SLICE_X4Y103_BO6),
.I1(CLBLM_R_X5Y104_SLICE_X7Y104_BQ),
.I2(CLBLM_R_X5Y104_SLICE_X7Y104_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y104_SLICE_X7Y104_BO5),
.O6(CLBLM_R_X5Y104_SLICE_X7Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00a1a10000)
  ) CLBLM_R_X5Y104_SLICE_X7Y104_ALUT (
.I0(CLBLL_L_X4Y103_SLICE_X4Y103_BO6),
.I1(CLBLM_R_X5Y104_SLICE_X7Y104_BQ),
.I2(CLBLM_R_X5Y104_SLICE_X7Y104_AQ),
.I3(CLBLM_R_X5Y103_SLICE_X6Y103_BQ),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X5Y104_SLICE_X7Y104_AO5),
.O6(CLBLM_R_X5Y104_SLICE_X7Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y105_SLICE_X6Y105_AO6),
.Q(CLBLM_R_X5Y105_SLICE_X6Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y105_SLICE_X6Y105_BO6),
.Q(CLBLM_R_X5Y105_SLICE_X6Y105_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hefffccffffffffff)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_DLUT (
.I0(CLBLM_R_X5Y106_SLICE_X6Y106_AO6),
.I1(CLBLM_R_X5Y105_SLICE_X6Y105_AQ),
.I2(CLBLM_R_X5Y107_SLICE_X6Y107_DQ),
.I3(CLBLM_R_X5Y105_SLICE_X6Y105_BQ),
.I4(CLBLM_R_X3Y105_SLICE_X3Y105_AQ),
.I5(CLBLM_R_X5Y106_SLICE_X7Y106_AQ),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_DO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff7fffffaaaa0000)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_CLUT (
.I0(CLBLM_R_X5Y104_SLICE_X6Y104_AQ),
.I1(CLBLM_R_X5Y105_SLICE_X7Y105_AQ),
.I2(CLBLM_R_X5Y105_SLICE_X6Y105_BQ),
.I3(CLBLM_R_X5Y106_SLICE_X6Y106_CO6),
.I4(CLBLM_R_X5Y104_SLICE_X6Y104_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_CO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff09ff0900090009)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_BLUT (
.I0(CLBLM_R_X5Y106_SLICE_X6Y106_CO6),
.I1(CLBLM_R_X5Y105_SLICE_X6Y105_BQ),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(1'b1),
.I5(CLBLM_R_X5Y106_SLICE_X7Y106_AQ),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_BO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888b88b9a8b)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_ALUT (
.I0(CLBLM_R_X5Y107_SLICE_X6Y107_DQ),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_R_X5Y105_SLICE_X6Y105_AQ),
.I3(CLBLM_R_X3Y105_SLICE_X3Y105_AQ),
.I4(CLBLM_R_X5Y106_SLICE_X6Y106_AO6),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_AO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y105_SLICE_X7Y105_AO6),
.Q(CLBLM_R_X5Y105_SLICE_X7Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_DO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffbfffffffff)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_CLUT (
.I0(CLBLM_R_X5Y105_SLICE_X6Y105_AQ),
.I1(CLBLM_R_X5Y106_SLICE_X7Y106_AQ),
.I2(CLBLM_R_X5Y105_SLICE_X6Y105_CO5),
.I3(CLBLM_R_X5Y106_SLICE_X6Y106_BO6),
.I4(CLBLM_R_X5Y105_SLICE_X7Y105_AQ),
.I5(CLBLM_R_X5Y105_SLICE_X6Y105_BQ),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_CO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000008000)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_BLUT (
.I0(CLBLM_R_X5Y104_SLICE_X6Y104_BQ),
.I1(CLBLM_R_X5Y106_SLICE_X7Y106_AQ),
.I2(CLBLM_R_X5Y104_SLICE_X6Y104_AQ),
.I3(CLBLM_R_X5Y105_SLICE_X6Y105_BQ),
.I4(CLBLM_R_X5Y105_SLICE_X6Y105_AQ),
.I5(CLBLM_R_X5Y106_SLICE_X6Y106_BO6),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_BO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff22ff1200220022)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_ALUT (
.I0(CLBLM_R_X5Y105_SLICE_X7Y105_AQ),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(CLBLM_R_X5Y104_SLICE_X6Y104_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLM_R_X5Y105_SLICE_X6Y105_DO6),
.I5(CLBLM_R_X5Y104_SLICE_X6Y104_BQ),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_AO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffeeffffaaaaaaaa)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_DLUT (
.I0(CLBLM_R_X5Y105_SLICE_X6Y105_AQ),
.I1(CLBLM_R_X5Y107_SLICE_X6Y107_CQ),
.I2(1'b1),
.I3(CLBLM_R_X5Y106_SLICE_X6Y106_AO5),
.I4(CLBLM_R_X5Y107_SLICE_X6Y107_DQ),
.I5(CLBLM_R_X3Y105_SLICE_X3Y105_AQ),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_DO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffdfffff5f5f5f5)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_CLUT (
.I0(CLBLM_R_X5Y106_SLICE_X7Y106_AQ),
.I1(CLBLM_R_X5Y107_SLICE_X6Y107_CQ),
.I2(CLBLM_R_X5Y105_SLICE_X6Y105_AQ),
.I3(CLBLM_R_X5Y106_SLICE_X6Y106_AO5),
.I4(CLBLM_R_X5Y107_SLICE_X6Y107_DQ),
.I5(CLBLM_R_X3Y105_SLICE_X3Y105_AQ),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_CO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0d0f0f0f0f0f0)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_BLUT (
.I0(CLBLM_R_X5Y107_SLICE_X6Y107_DQ),
.I1(CLBLM_R_X3Y106_SLICE_X3Y106_BO6),
.I2(CLBLM_R_X3Y105_SLICE_X3Y105_AQ),
.I3(CLBLM_R_X5Y107_SLICE_X6Y107_BQ),
.I4(CLBLM_R_X5Y107_SLICE_X6Y107_CQ),
.I5(CLBLM_R_X5Y107_SLICE_X6Y107_AQ),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_BO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff7fff7fff7ff)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_ALUT (
.I0(CLBLM_R_X3Y106_SLICE_X3Y106_DO6),
.I1(CLBLM_R_X5Y107_SLICE_X6Y107_BQ),
.I2(CLBLL_L_X2Y108_SLICE_X0Y108_BQ),
.I3(CLBLM_R_X5Y107_SLICE_X6Y107_AQ),
.I4(CLBLM_R_X5Y107_SLICE_X6Y107_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_AO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y106_SLICE_X7Y106_AO6),
.Q(CLBLM_R_X5Y106_SLICE_X7Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_DO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_CO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_BO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hb88b8888b88b8888)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_ALUT (
.I0(CLBLM_R_X5Y105_SLICE_X6Y105_AQ),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_R_X5Y106_SLICE_X7Y106_AQ),
.I3(CLBLM_R_X5Y106_SLICE_X6Y106_DO6),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_AO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y107_SLICE_X6Y107_AO6),
.Q(CLBLM_R_X5Y107_SLICE_X6Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y107_SLICE_X6Y107_BO6),
.Q(CLBLM_R_X5Y107_SLICE_X6Y107_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y107_SLICE_X6Y107_CO6),
.Q(CLBLM_R_X5Y107_SLICE_X6Y107_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y107_SLICE_X6Y107_DO6),
.Q(CLBLM_R_X5Y107_SLICE_X6Y107_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc50415041)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X5Y107_SLICE_X6Y107_CQ),
.I2(CLBLM_R_X5Y107_SLICE_X6Y107_DQ),
.I3(CLBLM_R_X5Y106_SLICE_X6Y106_AO5),
.I4(1'b1),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_DO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f044114411)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLM_R_X5Y107_SLICE_X6Y107_CQ),
.I2(CLBLM_R_X5Y107_SLICE_X6Y107_BQ),
.I3(CLBLM_R_X5Y106_SLICE_X6Y106_AO5),
.I4(1'b1),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_CO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0dff000f020f000)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_BLUT (
.I0(CLBLM_R_X3Y106_SLICE_X3Y106_DO6),
.I1(CLBLL_L_X2Y108_SLICE_X0Y108_BQ),
.I2(CLBLM_R_X5Y107_SLICE_X6Y107_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLM_R_X5Y107_SLICE_X6Y107_BQ),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_BO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccd2d20000)
  ) CLBLM_R_X5Y107_SLICE_X6Y107_ALUT (
.I0(CLBLM_R_X3Y106_SLICE_X3Y106_DO6),
.I1(CLBLL_L_X2Y108_SLICE_X0Y108_BQ),
.I2(CLBLM_R_X5Y107_SLICE_X6Y107_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X5Y107_SLICE_X6Y107_AO5),
.O6(CLBLM_R_X5Y107_SLICE_X6Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_DO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_CO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_BO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y107_SLICE_X7Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y107_SLICE_X7Y107_AO5),
.O6(CLBLM_R_X5Y107_SLICE_X7Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(LIOB33_X0Y127_IOB_X0Y128_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y101_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y101_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y102_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y102_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y103_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y103_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y104_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y104_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y105_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y105_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y106_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y106_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y107_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y107_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y108_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y108_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y109_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y109_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y110_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y110_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y111_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y111_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y112_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y112_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y113_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y113_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y114_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y114_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y115_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y115_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y116_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y116_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y117_IOB_X0Y117_IBUF (
.I(LIOB33_X0Y117_IOB_X0Y117_IPAD),
.O(LIOB33_X0Y117_IOB_X0Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y117_IOB_X0Y118_IBUF (
.I(LIOB33_X0Y117_IOB_X0Y118_IPAD),
.O(LIOB33_X0Y117_IOB_X0Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUF (
.I(CLBLL_L_X2Y108_SLICE_X0Y108_CO6),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUF (
.I(CLBLL_L_X4Y104_SLICE_X4Y104_DO6),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUF (
.I(CLBLL_L_X2Y105_SLICE_X1Y105_BQ),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUF (
.I(CLBLL_L_X2Y107_SLICE_X0Y107_AO5),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUF (
.I(CLBLL_L_X2Y106_SLICE_X0Y106_BQ),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(CLBLL_L_X2Y106_SLICE_X0Y106_BQ),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y127_IOB_X0Y128_IBUF (
.I(LIOB33_X0Y127_IOB_X0Y128_IPAD),
.O(LIOB33_X0Y127_IOB_X0Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y100_IOB_X0Y100_IBUF (
.I(LIOB33_SING_X0Y100_IOB_X0Y100_IPAD),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_I)
  );
  assign CLBLL_L_X2Y103_SLICE_X0Y103_A = CLBLL_L_X2Y103_SLICE_X0Y103_AO6;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_B = CLBLL_L_X2Y103_SLICE_X0Y103_BO6;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_C = CLBLL_L_X2Y103_SLICE_X0Y103_CO6;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_D = CLBLL_L_X2Y103_SLICE_X0Y103_DO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_A = CLBLL_L_X2Y103_SLICE_X1Y103_AO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_B = CLBLL_L_X2Y103_SLICE_X1Y103_BO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_C = CLBLL_L_X2Y103_SLICE_X1Y103_CO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_D = CLBLL_L_X2Y103_SLICE_X1Y103_DO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_CMUX = CLBLL_L_X2Y103_SLICE_X1Y103_CO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A = CLBLL_L_X2Y104_SLICE_X0Y104_AO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B = CLBLL_L_X2Y104_SLICE_X0Y104_BO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C = CLBLL_L_X2Y104_SLICE_X0Y104_CO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D = CLBLL_L_X2Y104_SLICE_X0Y104_DO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_CMUX = CLBLL_L_X2Y104_SLICE_X0Y104_CO5;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A = CLBLL_L_X2Y104_SLICE_X1Y104_AO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B = CLBLL_L_X2Y104_SLICE_X1Y104_BO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C = CLBLL_L_X2Y104_SLICE_X1Y104_CO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D = CLBLL_L_X2Y104_SLICE_X1Y104_DO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_AMUX = CLBLL_L_X2Y104_SLICE_X1Y104_AO5;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A = CLBLL_L_X2Y105_SLICE_X0Y105_AO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B = CLBLL_L_X2Y105_SLICE_X0Y105_BO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C = CLBLL_L_X2Y105_SLICE_X0Y105_CO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D = CLBLL_L_X2Y105_SLICE_X0Y105_DO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A = CLBLL_L_X2Y105_SLICE_X1Y105_AO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B = CLBLL_L_X2Y105_SLICE_X1Y105_BO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C = CLBLL_L_X2Y105_SLICE_X1Y105_CO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D = CLBLL_L_X2Y105_SLICE_X1Y105_DO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_AMUX = CLBLL_L_X2Y105_SLICE_X1Y105_AO5;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A = CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B = CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C = CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D = CLBLL_L_X2Y106_SLICE_X0Y106_DO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_AMUX = CLBLL_L_X2Y106_SLICE_X0Y106_AO5;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_CMUX = CLBLL_L_X2Y106_SLICE_X0Y106_CO5;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A = CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B = CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C = CLBLL_L_X2Y106_SLICE_X1Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D = CLBLL_L_X2Y106_SLICE_X1Y106_DO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_AMUX = CLBLL_L_X2Y106_SLICE_X1Y106_A5Q;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_CMUX = CLBLL_L_X2Y106_SLICE_X1Y106_CO5;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B = CLBLL_L_X2Y107_SLICE_X0Y107_BO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C = CLBLL_L_X2Y107_SLICE_X0Y107_CO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D = CLBLL_L_X2Y107_SLICE_X0Y107_DO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_AMUX = CLBLL_L_X2Y107_SLICE_X0Y107_AO5;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_DMUX = CLBLL_L_X2Y107_SLICE_X0Y107_DO5;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A = CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B = CLBLL_L_X2Y107_SLICE_X1Y107_BO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C = CLBLL_L_X2Y107_SLICE_X1Y107_CO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D = CLBLL_L_X2Y107_SLICE_X1Y107_DO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_DMUX = CLBLL_L_X2Y107_SLICE_X1Y107_DO5;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A = CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B = CLBLL_L_X2Y108_SLICE_X0Y108_BO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C = CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D = CLBLL_L_X2Y108_SLICE_X0Y108_DO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_AMUX = CLBLL_L_X2Y108_SLICE_X0Y108_A5Q;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_BMUX = CLBLL_L_X2Y108_SLICE_X0Y108_BO5;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A = CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B = CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C = CLBLL_L_X2Y108_SLICE_X1Y108_CO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D = CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A = CLBLL_L_X4Y103_SLICE_X4Y103_AO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B = CLBLL_L_X4Y103_SLICE_X4Y103_BO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C = CLBLL_L_X4Y103_SLICE_X4Y103_CO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D = CLBLL_L_X4Y103_SLICE_X4Y103_DO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A = CLBLL_L_X4Y103_SLICE_X5Y103_AO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B = CLBLL_L_X4Y103_SLICE_X5Y103_BO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C = CLBLL_L_X4Y103_SLICE_X5Y103_CO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D = CLBLL_L_X4Y103_SLICE_X5Y103_DO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A = CLBLL_L_X4Y104_SLICE_X4Y104_AO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B = CLBLL_L_X4Y104_SLICE_X4Y104_BO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C = CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D = CLBLL_L_X4Y104_SLICE_X4Y104_DO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_CMUX = CLBLL_L_X4Y104_SLICE_X4Y104_CO5;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A = CLBLL_L_X4Y104_SLICE_X5Y104_AO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B = CLBLL_L_X4Y104_SLICE_X5Y104_BO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C = CLBLL_L_X4Y104_SLICE_X5Y104_CO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D = CLBLL_L_X4Y104_SLICE_X5Y104_DO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_AMUX = CLBLL_L_X4Y104_SLICE_X5Y104_AO5;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_BMUX = CLBLL_L_X4Y104_SLICE_X5Y104_BO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A = CLBLL_L_X4Y105_SLICE_X4Y105_AO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B = CLBLL_L_X4Y105_SLICE_X4Y105_BO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C = CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D = CLBLL_L_X4Y105_SLICE_X4Y105_DO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A = CLBLL_L_X4Y105_SLICE_X5Y105_AO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C = CLBLL_L_X4Y105_SLICE_X5Y105_CO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D = CLBLL_L_X4Y105_SLICE_X5Y105_DO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A = CLBLL_L_X4Y106_SLICE_X4Y106_AO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B = CLBLL_L_X4Y106_SLICE_X4Y106_BO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C = CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D = CLBLL_L_X4Y106_SLICE_X4Y106_DO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_AMUX = CLBLL_L_X4Y106_SLICE_X4Y106_AO5;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_BMUX = CLBLL_L_X4Y106_SLICE_X4Y106_BO5;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_CMUX = CLBLL_L_X4Y106_SLICE_X4Y106_CO5;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A = CLBLL_L_X4Y106_SLICE_X5Y106_AO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B = CLBLL_L_X4Y106_SLICE_X5Y106_BO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C = CLBLL_L_X4Y106_SLICE_X5Y106_CO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D = CLBLL_L_X4Y106_SLICE_X5Y106_DO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A = CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B = CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C = CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D = CLBLL_L_X4Y107_SLICE_X4Y107_DO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A = CLBLL_L_X4Y107_SLICE_X5Y107_AO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B = CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C = CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D = CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A = CLBLM_R_X3Y103_SLICE_X2Y103_AO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B = CLBLM_R_X3Y103_SLICE_X2Y103_BO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C = CLBLM_R_X3Y103_SLICE_X2Y103_CO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D = CLBLM_R_X3Y103_SLICE_X2Y103_DO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A = CLBLM_R_X3Y103_SLICE_X3Y103_AO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B = CLBLM_R_X3Y103_SLICE_X3Y103_BO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C = CLBLM_R_X3Y103_SLICE_X3Y103_CO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D = CLBLM_R_X3Y103_SLICE_X3Y103_DO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A = CLBLM_R_X3Y104_SLICE_X2Y104_AO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B = CLBLM_R_X3Y104_SLICE_X2Y104_BO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C = CLBLM_R_X3Y104_SLICE_X2Y104_CO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D = CLBLM_R_X3Y104_SLICE_X2Y104_DO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A = CLBLM_R_X3Y104_SLICE_X3Y104_AO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B = CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C = CLBLM_R_X3Y104_SLICE_X3Y104_CO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D = CLBLM_R_X3Y104_SLICE_X3Y104_DO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A = CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B = CLBLM_R_X3Y105_SLICE_X2Y105_BO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C = CLBLM_R_X3Y105_SLICE_X2Y105_CO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D = CLBLM_R_X3Y105_SLICE_X2Y105_DO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_AMUX = CLBLM_R_X3Y105_SLICE_X2Y105_A5Q;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_BMUX = CLBLM_R_X3Y105_SLICE_X2Y105_B5Q;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_CMUX = CLBLM_R_X3Y105_SLICE_X2Y105_CO5;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_DMUX = CLBLM_R_X3Y105_SLICE_X2Y105_DO5;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A = CLBLM_R_X3Y105_SLICE_X3Y105_AO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B = CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C = CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D = CLBLM_R_X3Y105_SLICE_X3Y105_DO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A = CLBLM_R_X3Y106_SLICE_X2Y106_AO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B = CLBLM_R_X3Y106_SLICE_X2Y106_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C = CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D = CLBLM_R_X3Y106_SLICE_X2Y106_DO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_AMUX = CLBLM_R_X3Y106_SLICE_X2Y106_AO5;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_CMUX = CLBLM_R_X3Y106_SLICE_X2Y106_CO5;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A = CLBLM_R_X3Y106_SLICE_X3Y106_AO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B = CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C = CLBLM_R_X3Y106_SLICE_X3Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D = CLBLM_R_X3Y106_SLICE_X3Y106_DO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_AMUX = CLBLM_R_X3Y106_SLICE_X3Y106_AO5;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A = CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B = CLBLM_R_X3Y107_SLICE_X2Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C = CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D = CLBLM_R_X3Y107_SLICE_X2Y107_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A = CLBLM_R_X3Y107_SLICE_X3Y107_AO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B = CLBLM_R_X3Y107_SLICE_X3Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C = CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D = CLBLM_R_X3Y107_SLICE_X3Y107_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_AMUX = CLBLM_R_X3Y107_SLICE_X3Y107_AO5;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_BMUX = CLBLM_R_X3Y107_SLICE_X3Y107_BO5;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_DMUX = CLBLM_R_X3Y107_SLICE_X3Y107_DO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_A = CLBLM_R_X5Y103_SLICE_X6Y103_AO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_B = CLBLM_R_X5Y103_SLICE_X6Y103_BO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_C = CLBLM_R_X5Y103_SLICE_X6Y103_CO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_D = CLBLM_R_X5Y103_SLICE_X6Y103_DO6;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_A = CLBLM_R_X5Y103_SLICE_X7Y103_AO6;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_B = CLBLM_R_X5Y103_SLICE_X7Y103_BO6;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_C = CLBLM_R_X5Y103_SLICE_X7Y103_CO6;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_D = CLBLM_R_X5Y103_SLICE_X7Y103_DO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A = CLBLM_R_X5Y104_SLICE_X6Y104_AO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B = CLBLM_R_X5Y104_SLICE_X6Y104_BO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C = CLBLM_R_X5Y104_SLICE_X6Y104_CO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D = CLBLM_R_X5Y104_SLICE_X6Y104_DO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A = CLBLM_R_X5Y104_SLICE_X7Y104_AO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B = CLBLM_R_X5Y104_SLICE_X7Y104_BO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C = CLBLM_R_X5Y104_SLICE_X7Y104_CO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D = CLBLM_R_X5Y104_SLICE_X7Y104_DO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A = CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B = CLBLM_R_X5Y105_SLICE_X6Y105_BO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C = CLBLM_R_X5Y105_SLICE_X6Y105_CO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D = CLBLM_R_X5Y105_SLICE_X6Y105_DO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_CMUX = CLBLM_R_X5Y105_SLICE_X6Y105_CO5;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A = CLBLM_R_X5Y105_SLICE_X7Y105_AO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B = CLBLM_R_X5Y105_SLICE_X7Y105_BO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C = CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D = CLBLM_R_X5Y105_SLICE_X7Y105_DO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A = CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B = CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C = CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D = CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_AMUX = CLBLM_R_X5Y106_SLICE_X6Y106_AO5;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A = CLBLM_R_X5Y106_SLICE_X7Y106_AO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B = CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C = CLBLM_R_X5Y106_SLICE_X7Y106_CO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D = CLBLM_R_X5Y106_SLICE_X7Y106_DO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A = CLBLM_R_X5Y107_SLICE_X6Y107_AO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B = CLBLM_R_X5Y107_SLICE_X6Y107_BO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C = CLBLM_R_X5Y107_SLICE_X6Y107_CO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D = CLBLM_R_X5Y107_SLICE_X6Y107_DO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A = CLBLM_R_X5Y107_SLICE_X7Y107_AO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B = CLBLM_R_X5Y107_SLICE_X7Y107_BO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C = CLBLM_R_X5Y107_SLICE_X7Y107_CO6;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D = CLBLM_R_X5Y107_SLICE_X7Y107_DO6;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_O = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_O = LIOB33_X0Y101_IOB_X0Y101_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_O = LIOB33_X0Y103_IOB_X0Y104_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_O = LIOB33_X0Y103_IOB_X0Y103_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_O = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_O = LIOB33_X0Y105_IOB_X0Y105_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_O = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_O = LIOB33_X0Y109_IOB_X0Y109_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_O = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_O = LIOB33_X0Y111_IOB_X0Y111_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_O = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_O = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y118_O = LIOB33_X0Y117_IOB_X0Y118_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_O = LIOB33_X0Y117_IOB_X0Y117_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = CLBLL_L_X2Y107_SLICE_X0Y107_AO5;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = CLBLL_L_X2Y105_SLICE_X1Y105_BQ;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = CLBLL_L_X2Y106_SLICE_X0Y106_BQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = CLBLL_L_X2Y106_SLICE_X0Y106_BQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_O = LIOB33_X0Y127_IOB_X0Y128_I;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_O = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O = LIOB33_X0Y107_IOB_X0Y107_I;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = CLBLL_L_X4Y104_SLICE_X4Y104_DO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_A1 = CLBLM_R_X3Y105_SLICE_X3Y105_AQ;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_A2 = CLBLM_R_X5Y105_SLICE_X7Y105_BO6;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_A3 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_A4 = CLBLM_R_X5Y103_SLICE_X6Y103_BQ;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_A5 = CLBLM_R_X5Y105_SLICE_X7Y105_AQ;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_A6 = CLBLM_R_X5Y103_SLICE_X6Y103_CQ;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_B1 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_B2 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_B3 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_B4 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_B5 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_B6 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A1 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A2 = CLBLL_L_X2Y105_SLICE_X0Y105_BQ;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A3 = CLBLL_L_X2Y107_SLICE_X1Y107_AQ;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A4 = CLBLL_L_X4Y107_SLICE_X4Y107_AQ;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A5 = CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A6 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_C1 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_C2 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_C3 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B1 = CLBLL_L_X4Y106_SLICE_X4Y106_DO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B2 = CLBLM_R_X3Y107_SLICE_X3Y107_AO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B3 = CLBLM_R_X3Y107_SLICE_X3Y107_AO5;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B4 = CLBLM_R_X3Y107_SLICE_X3Y107_DO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B5 = CLBLL_L_X2Y108_SLICE_X0Y108_BQ;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B6 = CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_D4 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C1 = CLBLL_L_X4Y107_SLICE_X4Y107_AQ;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C2 = CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C3 = CLBLM_R_X3Y107_SLICE_X3Y107_AO5;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C4 = CLBLM_R_X3Y106_SLICE_X3Y106_AO5;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C5 = CLBLM_R_X3Y107_SLICE_X3Y107_BO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C6 = CLBLL_L_X4Y106_SLICE_X4Y106_AO6;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_D2 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_D3 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_D5 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_A1 = CLBLM_R_X5Y103_SLICE_X6Y103_CQ;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_A2 = CLBLM_R_X5Y103_SLICE_X6Y103_BQ;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_A3 = CLBLM_R_X5Y103_SLICE_X6Y103_AQ;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_A4 = CLBLM_R_X5Y104_SLICE_X6Y104_CO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_A6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_A5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D1 = CLBLM_R_X3Y106_SLICE_X3Y106_AO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D2 = CLBLM_R_X3Y107_SLICE_X3Y107_AO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D3 = CLBLM_R_X3Y107_SLICE_X3Y107_AO5;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_B1 = CLBLM_R_X5Y103_SLICE_X6Y103_CQ;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_B2 = CLBLM_R_X5Y103_SLICE_X6Y103_BQ;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_B3 = CLBLM_R_X5Y103_SLICE_X6Y103_AQ;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_B4 = CLBLM_R_X5Y104_SLICE_X6Y104_CO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_B5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D4 = CLBLL_L_X4Y106_SLICE_X4Y106_DO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D5 = CLBLM_R_X3Y107_SLICE_X3Y107_BO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D6 = CLBLM_R_X3Y107_SLICE_X3Y107_DO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_C1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_C2 = CLBLM_R_X5Y103_SLICE_X6Y103_CQ;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A1 = CLBLL_L_X2Y107_SLICE_X1Y107_DO5;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_C4 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_C5 = CLBLM_R_X5Y104_SLICE_X6Y104_CO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_C3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_C6 = CLBLL_L_X4Y104_SLICE_X4Y104_BQ;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A3 = CLBLM_R_X3Y106_SLICE_X2Y106_AQ;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A5 = CLBLM_R_X3Y106_SLICE_X2Y106_BQ;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A6 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B1 = CLBLL_L_X2Y107_SLICE_X1Y107_DO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B2 = CLBLM_R_X3Y106_SLICE_X2Y106_BQ;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_D1 = CLBLM_R_X5Y105_SLICE_X7Y105_AQ;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B4 = CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_D3 = CLBLM_R_X5Y103_SLICE_X6Y103_AQ;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_D4 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_D5 = CLBLM_R_X3Y105_SLICE_X3Y105_AQ;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_D6 = CLBLM_R_X5Y105_SLICE_X7Y105_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C4 = CLBLL_L_X2Y103_SLICE_X1Y103_CO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C6 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D1 = CLBLM_R_X3Y106_SLICE_X2Y106_BQ;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D2 = CLBLL_L_X2Y107_SLICE_X0Y107_CQ;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D4 = CLBLL_L_X2Y107_SLICE_X0Y107_BQ;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D5 = CLBLL_L_X2Y105_SLICE_X0Y105_BQ;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D6 = CLBLL_L_X2Y106_SLICE_X1Y106_AQ;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0 = LIOB33_X0Y127_IOB_X0Y128_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X6Y103_D2 = CLBLM_R_X5Y103_SLICE_X6Y103_CQ;
  assign LIOB33_X0Y121_IOB_X0Y122_O = CLBLL_L_X2Y107_SLICE_X0Y107_AO5;
  assign LIOB33_X0Y121_IOB_X0Y121_O = CLBLL_L_X2Y105_SLICE_X1Y105_BQ;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A1 = CLBLL_L_X4Y103_SLICE_X4Y103_BO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A2 = CLBLM_R_X5Y104_SLICE_X7Y104_BQ;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A3 = CLBLM_R_X5Y104_SLICE_X7Y104_AQ;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A4 = CLBLM_R_X5Y103_SLICE_X6Y103_BQ;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_A6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B1 = CLBLL_L_X4Y103_SLICE_X4Y103_BO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B2 = CLBLM_R_X5Y104_SLICE_X7Y104_BQ;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B3 = CLBLM_R_X5Y104_SLICE_X7Y104_AQ;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_B6 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A1 = CLBLL_L_X2Y107_SLICE_X1Y107_BQ;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A2 = CLBLL_L_X2Y105_SLICE_X0Y105_BQ;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A3 = CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A4 = CLBLL_L_X4Y107_SLICE_X4Y107_BQ;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A5 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A6 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C1 = CLBLM_R_X5Y103_SLICE_X6Y103_CQ;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C2 = CLBLM_R_X5Y105_SLICE_X7Y105_AQ;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C3 = CLBLL_L_X2Y105_SLICE_X0Y105_CQ;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B1 = CLBLL_L_X4Y107_SLICE_X4Y107_CQ;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B2 = CLBLL_L_X2Y105_SLICE_X0Y105_BQ;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B3 = CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B4 = CLBLL_L_X2Y107_SLICE_X1Y107_CQ;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B5 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B6 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D1 = CLBLM_R_X5Y103_SLICE_X6Y103_CQ;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C1 = CLBLL_L_X4Y107_SLICE_X4Y107_AQ;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C2 = CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C3 = CLBLL_L_X4Y107_SLICE_X4Y107_CQ;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C4 = CLBLM_R_X3Y107_SLICE_X2Y107_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C5 = CLBLM_R_X3Y107_SLICE_X3Y107_BO5;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C6 = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D3 = CLBLL_L_X2Y105_SLICE_X0Y105_CQ;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D4 = CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A1 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A2 = CLBLM_R_X5Y105_SLICE_X6Y105_BQ;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A3 = CLBLM_R_X5Y104_SLICE_X6Y104_AQ;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D1 = CLBLL_L_X4Y107_SLICE_X4Y107_AQ;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D2 = CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_A6 = CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D3 = CLBLM_R_X3Y107_SLICE_X2Y107_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D4 = CLBLL_L_X4Y107_SLICE_X4Y107_CQ;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D5 = CLBLM_R_X3Y107_SLICE_X3Y107_BO5;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D6 = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B4 = CLBLM_R_X5Y105_SLICE_X6Y105_BQ;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B1 = CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A1 = CLBLL_L_X2Y107_SLICE_X0Y107_DO5;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A2 = CLBLM_R_X3Y107_SLICE_X2Y107_BQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A3 = CLBLM_R_X3Y107_SLICE_X2Y107_AQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A6 = CLBLL_L_X2Y107_SLICE_X0Y107_DO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C1 = CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C1 = CLBLM_R_X5Y104_SLICE_X6Y104_BQ;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C2 = CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B1 = CLBLL_L_X2Y107_SLICE_X0Y107_DO5;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C2 = CLBLL_L_X4Y106_SLICE_X4Y106_AQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B2 = CLBLM_R_X3Y107_SLICE_X2Y107_BQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B4 = CLBLL_L_X4Y107_SLICE_X5Y107_BQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B6 = CLBLL_L_X2Y107_SLICE_X0Y107_DO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D1 = CLBLL_L_X4Y103_SLICE_X5Y103_DO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C1 = CLBLL_L_X2Y107_SLICE_X0Y107_BQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C3 = CLBLL_L_X2Y107_SLICE_X0Y107_CQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C4 = CLBLL_L_X2Y106_SLICE_X1Y106_AQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C5 = CLBLL_L_X2Y107_SLICE_X1Y107_CQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C6 = CLBLL_L_X2Y105_SLICE_X0Y105_BQ;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D2 = CLBLL_L_X4Y103_SLICE_X4Y103_BO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D3 = CLBLM_R_X5Y104_SLICE_X7Y104_DO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D5 = CLBLL_L_X4Y105_SLICE_X4Y105_DO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C6 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D1 = CLBLL_L_X2Y107_SLICE_X0Y107_BQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D3 = CLBLL_L_X2Y107_SLICE_X0Y107_CQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D4 = CLBLL_L_X2Y106_SLICE_X1Y106_AQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D5 = CLBLL_L_X2Y107_SLICE_X1Y107_AQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D6 = CLBLL_L_X2Y105_SLICE_X0Y105_BQ;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_D = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_D = LIOB33_X0Y111_IOB_X0Y111_I;
  assign LIOB33_X0Y123_IOB_X0Y124_O = CLBLL_L_X2Y106_SLICE_X0Y106_BQ;
  assign LIOB33_X0Y123_IOB_X0Y123_O = CLBLL_L_X2Y106_SLICE_X0Y106_BQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A1 = CLBLM_R_X5Y105_SLICE_X7Y105_AQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A3 = CLBLM_R_X5Y104_SLICE_X6Y104_AQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A5 = CLBLM_R_X5Y105_SLICE_X6Y105_DO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A6 = CLBLM_R_X5Y104_SLICE_X6Y104_BQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B1 = CLBLM_R_X5Y104_SLICE_X6Y104_BQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B2 = CLBLM_R_X5Y106_SLICE_X7Y106_AQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B3 = CLBLM_R_X5Y104_SLICE_X6Y104_AQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B4 = CLBLM_R_X5Y105_SLICE_X6Y105_BQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B5 = CLBLM_R_X5Y105_SLICE_X6Y105_AQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B6 = CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C1 = CLBLM_R_X5Y105_SLICE_X6Y105_AQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C2 = CLBLM_R_X5Y106_SLICE_X7Y106_AQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C3 = CLBLM_R_X5Y105_SLICE_X6Y105_CO5;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C4 = CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C5 = CLBLM_R_X5Y105_SLICE_X7Y105_AQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C6 = CLBLM_R_X5Y105_SLICE_X6Y105_BQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D1 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D2 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D3 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D4 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D5 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D6 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A1 = CLBLM_R_X5Y107_SLICE_X6Y107_DQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A3 = CLBLM_R_X5Y105_SLICE_X6Y105_AQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A4 = CLBLM_R_X3Y105_SLICE_X3Y105_AQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A5 = CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B1 = CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B2 = CLBLM_R_X5Y105_SLICE_X6Y105_BQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B5 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B6 = CLBLM_R_X5Y106_SLICE_X7Y106_AQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C1 = CLBLM_R_X5Y104_SLICE_X6Y104_AQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C2 = CLBLM_R_X5Y105_SLICE_X7Y105_AQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C3 = CLBLM_R_X5Y105_SLICE_X6Y105_BQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C4 = CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C5 = CLBLM_R_X5Y104_SLICE_X6Y104_BQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C6 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B5 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B6 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D1 = CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D2 = CLBLM_R_X5Y105_SLICE_X6Y105_AQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D3 = CLBLM_R_X5Y107_SLICE_X6Y107_DQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D4 = CLBLM_R_X5Y105_SLICE_X6Y105_BQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D5 = CLBLM_R_X3Y105_SLICE_X3Y105_AQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D6 = CLBLM_R_X5Y106_SLICE_X7Y106_AQ;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C4 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C5 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C6 = 1'b1;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_D = LIOB33_X0Y127_IOB_X0Y128_I;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C6 = CLBLM_R_X3Y103_SLICE_X3Y103_DO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A1 = CLBLM_R_X5Y105_SLICE_X6Y105_AQ;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A3 = CLBLM_R_X5Y106_SLICE_X7Y106_AQ;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A4 = CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A6 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B1 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B2 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B3 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B4 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B5 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B6 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C1 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C2 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C3 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C4 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C5 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C6 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D1 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D2 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D3 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D4 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D5 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D6 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A1 = CLBLM_R_X3Y106_SLICE_X3Y106_DO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A2 = CLBLM_R_X5Y107_SLICE_X6Y107_BQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A3 = CLBLL_L_X2Y108_SLICE_X0Y108_BQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A4 = CLBLM_R_X5Y107_SLICE_X6Y107_AQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A5 = CLBLM_R_X5Y107_SLICE_X6Y107_CQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A6 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B1 = CLBLM_R_X5Y107_SLICE_X6Y107_DQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B2 = CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B3 = CLBLM_R_X3Y105_SLICE_X3Y105_AQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B4 = CLBLM_R_X5Y107_SLICE_X6Y107_BQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B5 = CLBLM_R_X5Y107_SLICE_X6Y107_CQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B6 = CLBLM_R_X5Y107_SLICE_X6Y107_AQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C1 = CLBLM_R_X5Y106_SLICE_X7Y106_AQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C2 = CLBLM_R_X5Y107_SLICE_X6Y107_CQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C3 = CLBLM_R_X5Y105_SLICE_X6Y105_AQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C4 = CLBLM_R_X5Y106_SLICE_X6Y106_AO5;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C5 = CLBLM_R_X5Y107_SLICE_X6Y107_DQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C6 = CLBLM_R_X3Y105_SLICE_X3Y105_AQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D1 = CLBLM_R_X5Y105_SLICE_X6Y105_AQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D2 = CLBLM_R_X5Y107_SLICE_X6Y107_CQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D3 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D4 = CLBLM_R_X5Y106_SLICE_X6Y106_AO5;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D5 = CLBLM_R_X5Y107_SLICE_X6Y107_DQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D6 = CLBLM_R_X3Y105_SLICE_X3Y105_AQ;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A2 = CLBLL_L_X4Y103_SLICE_X5Y103_DO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A3 = CLBLL_L_X4Y103_SLICE_X4Y103_AQ;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A5 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_A6 = CLBLL_L_X4Y103_SLICE_X5Y103_CQ;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B1 = CLBLL_L_X4Y105_SLICE_X5Y105_DO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B2 = CLBLL_L_X2Y105_SLICE_X1Y105_CO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B3 = CLBLL_L_X4Y103_SLICE_X4Y103_AQ;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B4 = CLBLM_R_X5Y104_SLICE_X6Y104_CO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B5 = CLBLM_R_X3Y103_SLICE_X3Y103_BQ;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_B6 = CLBLL_L_X4Y103_SLICE_X5Y103_CQ;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C1 = CLBLM_R_X3Y103_SLICE_X3Y103_BQ;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C2 = CLBLL_L_X2Y105_SLICE_X1Y105_CO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C3 = CLBLM_R_X5Y104_SLICE_X7Y104_BQ;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C4 = CLBLL_L_X4Y103_SLICE_X5Y103_CQ;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C5 = CLBLL_L_X4Y103_SLICE_X4Y103_DO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_C6 = CLBLL_L_X4Y105_SLICE_X5Y105_DO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D1 = CLBLM_R_X5Y105_SLICE_X7Y105_AQ;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D2 = CLBLL_L_X2Y105_SLICE_X1Y105_CO6;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D3 = CLBLL_L_X4Y103_SLICE_X4Y103_AQ;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D4 = CLBLM_R_X3Y105_SLICE_X3Y105_AQ;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D5 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X4Y103_D6 = CLBLM_R_X5Y105_SLICE_X7Y105_BO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A2 = CLBLL_L_X4Y103_SLICE_X5Y103_BQ;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A3 = CLBLL_L_X4Y103_SLICE_X5Y103_AQ;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A5 = CLBLL_L_X4Y104_SLICE_X4Y104_CO5;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_A6 = CLBLL_L_X4Y105_SLICE_X5Y105_BQ;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B1 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B2 = CLBLL_L_X4Y103_SLICE_X5Y103_BQ;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B3 = CLBLL_L_X4Y103_SLICE_X5Y103_AQ;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_B6 = CLBLL_L_X4Y104_SLICE_X4Y104_CO5;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A1 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A2 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A6 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C2 = CLBLL_L_X4Y104_SLICE_X5Y104_CO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C3 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C4 = CLBLM_R_X3Y103_SLICE_X3Y103_BQ;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C5 = CLBLL_L_X4Y103_SLICE_X5Y103_CQ;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B3 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B4 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B5 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B6 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_C6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B1 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_B2 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C2 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C3 = 1'b1;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D1 = CLBLL_L_X4Y104_SLICE_X5Y104_DO6;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D2 = CLBLL_L_X4Y103_SLICE_X5Y103_CQ;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D3 = CLBLL_L_X2Y105_SLICE_X0Y105_CQ;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D4 = CLBLM_R_X3Y103_SLICE_X3Y103_BQ;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D5 = CLBLL_L_X4Y105_SLICE_X5Y105_CQ;
  assign CLBLL_L_X4Y103_SLICE_X5Y103_D6 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C4 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C5 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C6 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D1 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D2 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D3 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D4 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D5 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_D6 = 1'b1;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_D = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A1 = CLBLM_R_X3Y106_SLICE_X3Y106_DO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A2 = CLBLL_L_X2Y108_SLICE_X0Y108_BQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A3 = CLBLM_R_X5Y107_SLICE_X6Y107_AQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A4 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_A6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_D = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B1 = CLBLM_R_X3Y106_SLICE_X3Y106_DO6;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B2 = CLBLL_L_X2Y108_SLICE_X0Y108_BQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B3 = CLBLM_R_X5Y107_SLICE_X6Y107_AQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_B6 = CLBLM_R_X5Y107_SLICE_X6Y107_BQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C2 = CLBLM_R_X5Y107_SLICE_X6Y107_CQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C3 = CLBLM_R_X5Y107_SLICE_X6Y107_BQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C4 = CLBLM_R_X5Y106_SLICE_X6Y106_AO5;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C5 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_C6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D2 = CLBLM_R_X5Y107_SLICE_X6Y107_CQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D3 = CLBLM_R_X5Y107_SLICE_X6Y107_DQ;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D4 = CLBLM_R_X5Y106_SLICE_X6Y106_AO5;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D5 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X6Y107_D6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C4 = CLBLM_R_X5Y105_SLICE_X7Y105_BO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C5 = CLBLM_R_X3Y105_SLICE_X3Y105_AQ;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_C6 = CLBLM_R_X5Y103_SLICE_X6Y103_BQ;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D3 = CLBLL_L_X4Y104_SLICE_X5Y104_BO6;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D5 = CLBLM_R_X3Y105_SLICE_X3Y105_AQ;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D4 = CLBLM_R_X3Y104_SLICE_X2Y104_BQ;
  assign CLBLM_R_X5Y104_SLICE_X7Y104_D6 = CLBLM_R_X5Y103_SLICE_X6Y103_BQ;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A2 = CLBLL_L_X4Y104_SLICE_X4Y104_BQ;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A3 = CLBLL_L_X4Y104_SLICE_X4Y104_AQ;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A5 = CLBLM_R_X3Y104_SLICE_X3Y104_BQ;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A6 = CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B2 = CLBLL_L_X4Y104_SLICE_X4Y104_BQ;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B3 = CLBLL_L_X4Y104_SLICE_X4Y104_AQ;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B5 = CLBLM_R_X3Y104_SLICE_X3Y104_BQ;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B6 = CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_A1 = CLBLL_L_X2Y104_SLICE_X0Y104_AQ;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_A2 = CLBLL_L_X2Y104_SLICE_X0Y104_CO6;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_A6 = CLBLL_L_X2Y103_SLICE_X0Y103_CO6;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C1 = CLBLL_L_X4Y103_SLICE_X4Y103_BO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C2 = CLBLL_L_X4Y105_SLICE_X5Y105_BQ;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C3 = CLBLL_L_X4Y104_SLICE_X4Y104_BQ;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C4 = CLBLM_R_X5Y104_SLICE_X7Y104_BQ;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C5 = CLBLL_L_X2Y105_SLICE_X0Y105_CQ;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C6 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_A5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_B1 = CLBLL_L_X2Y103_SLICE_X0Y103_DO6;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_B2 = CLBLL_L_X2Y104_SLICE_X0Y104_CO6;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_B3 = CLBLL_L_X2Y103_SLICE_X0Y103_AQ;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_B4 = CLBLL_L_X2Y106_SLICE_X1Y106_BQ;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D1 = CLBLL_L_X4Y104_SLICE_X5Y104_AQ;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D2 = CLBLL_L_X4Y104_SLICE_X4Y104_CO5;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_B6 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D5 = CLBLL_L_X4Y103_SLICE_X5Y103_BQ;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_C1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_C2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_C3 = CLBLL_L_X2Y106_SLICE_X1Y106_BQ;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D6 = CLBLL_L_X4Y105_SLICE_X4Y105_BO6;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_C4 = CLBLL_L_X2Y104_SLICE_X0Y104_CO5;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_C5 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_C6 = CLBLL_L_X2Y103_SLICE_X0Y103_AQ;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_D1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_D2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_D3 = CLBLL_L_X2Y106_SLICE_X1Y106_BQ;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_D4 = CLBLL_L_X2Y104_SLICE_X0Y104_CO5;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_D5 = CLBLL_L_X2Y103_SLICE_X0Y103_BQ;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_D6 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A1 = CLBLL_L_X4Y104_SLICE_X4Y104_CO5;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A3 = CLBLL_L_X4Y104_SLICE_X5Y104_AQ;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A4 = CLBLL_L_X4Y103_SLICE_X5Y103_BQ;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A6 = 1'b1;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B2 = CLBLM_R_X5Y104_SLICE_X6Y104_BQ;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_B3 = CLBLM_R_X5Y104_SLICE_X6Y104_AQ;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B1 = CLBLL_L_X4Y105_SLICE_X5Y105_AQ;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B2 = CLBLM_R_X5Y104_SLICE_X6Y104_CO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B3 = CLBLL_L_X4Y105_SLICE_X4Y105_AQ;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B4 = CLBLM_R_X3Y104_SLICE_X2Y104_AQ;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_A1 = CLBLM_R_X3Y103_SLICE_X2Y103_CQ;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_A2 = CLBLM_R_X3Y103_SLICE_X3Y103_CO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_A3 = CLBLL_L_X2Y103_SLICE_X1Y103_AQ;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_A5 = CLBLL_L_X2Y103_SLICE_X1Y103_CO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_A6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B5 = CLBLL_L_X4Y105_SLICE_X5Y105_CQ;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B6 = CLBLL_L_X2Y105_SLICE_X0Y105_BQ;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C2 = CLBLM_R_X5Y104_SLICE_X6Y104_CO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_B2 = CLBLL_L_X2Y103_SLICE_X1Y103_BQ;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_B3 = CLBLL_L_X2Y103_SLICE_X1Y103_AQ;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_B4 = CLBLL_L_X2Y104_SLICE_X1Y104_AO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_B6 = CLBLL_L_X2Y103_SLICE_X1Y103_CO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C3 = CLBLL_L_X4Y105_SLICE_X5Y105_CQ;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C5 = CLBLL_L_X4Y105_SLICE_X5Y105_AQ;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_C1 = CLBLL_L_X2Y103_SLICE_X1Y103_BQ;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_C2 = CLBLL_L_X2Y103_SLICE_X1Y103_DO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_C3 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_C4 = CLBLL_L_X2Y103_SLICE_X1Y103_AQ;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_C5 = CLBLL_L_X2Y104_SLICE_X0Y104_BQ;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_C6 = CLBLL_L_X2Y103_SLICE_X0Y103_BQ;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D1 = CLBLL_L_X4Y105_SLICE_X4Y105_AQ;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D2 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D3 = CLBLM_R_X5Y105_SLICE_X7Y105_AQ;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D4 = CLBLM_R_X3Y105_SLICE_X3Y105_AQ;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D5 = CLBLL_L_X4Y105_SLICE_X5Y105_AQ;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D6 = CLBLM_R_X5Y105_SLICE_X7Y105_BO6;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_D1 = CLBLL_L_X2Y103_SLICE_X0Y103_AQ;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_D2 = 1'b1;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_D3 = CLBLL_L_X2Y104_SLICE_X0Y104_AQ;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_D4 = CLBLM_R_X3Y103_SLICE_X2Y103_CQ;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_D5 = CLBLL_L_X2Y104_SLICE_X0Y104_BQ;
  assign CLBLL_L_X2Y103_SLICE_X1Y103_D6 = CLBLL_L_X2Y103_SLICE_X0Y103_BQ;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C3 = CLBLM_R_X5Y104_SLICE_X6Y104_AQ;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C4 = CLBLM_R_X5Y105_SLICE_X7Y105_AQ;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C5 = CLBLM_R_X3Y105_SLICE_X3Y105_AQ;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_C6 = CLBLM_R_X5Y105_SLICE_X6Y105_BQ;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_D = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_D = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A4 = CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D4 = CLBLM_R_X5Y103_SLICE_X6Y103_DO6;
  assign CLBLM_R_X5Y104_SLICE_X6Y104_D6 = CLBLM_R_X5Y104_SLICE_X7Y104_BQ;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C1 = CLBLL_L_X4Y105_SLICE_X4Y105_AQ;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C4 = CLBLL_L_X2Y105_SLICE_X0Y105_CQ;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C6 = CLBLM_R_X3Y103_SLICE_X3Y103_BQ;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B5 = CLBLL_L_X2Y104_SLICE_X0Y104_BQ;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B6 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C2 = CLBLL_L_X2Y105_SLICE_X0Y105_BQ;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A1 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A3 = CLBLL_L_X4Y105_SLICE_X4Y105_AQ;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A4 = CLBLM_R_X5Y104_SLICE_X6Y104_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A5 = CLBLL_L_X4Y103_SLICE_X4Y103_AQ;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B1 = CLBLM_R_X5Y107_SLICE_X6Y107_DQ;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B2 = CLBLM_R_X5Y105_SLICE_X7Y105_BO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B3 = CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B4 = CLBLL_L_X2Y105_SLICE_X0Y105_DQ;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A1 = CLBLL_L_X2Y104_SLICE_X1Y104_AO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A2 = CLBLL_L_X2Y103_SLICE_X1Y103_CO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A3 = CLBLL_L_X2Y104_SLICE_X0Y104_AQ;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A4 = CLBLL_L_X2Y103_SLICE_X1Y103_BQ;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_A6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C1 = CLBLL_L_X4Y103_SLICE_X4Y103_AQ;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C2 = CLBLL_L_X4Y103_SLICE_X5Y103_DO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B5 = CLBLM_R_X5Y105_SLICE_X7Y105_AQ;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C4 = CLBLL_L_X2Y105_SLICE_X1Y105_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C5 = CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C6 = CLBLM_R_X3Y105_SLICE_X3Y105_AQ;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B1 = CLBLL_L_X2Y104_SLICE_X0Y104_DO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B3 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B4 = CLBLL_L_X2Y106_SLICE_X1Y106_BQ;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B5 = CLBLL_L_X2Y103_SLICE_X0Y103_BQ;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_B6 = CLBLL_L_X2Y104_SLICE_X0Y104_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D2 = CLBLL_L_X4Y105_SLICE_X4Y105_AQ;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D1 = CLBLL_L_X4Y105_SLICE_X5Y105_AQ;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C2 = CLBLL_L_X2Y103_SLICE_X1Y103_CO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C3 = CLBLL_L_X2Y105_SLICE_X0Y105_BQ;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D4 = CLBLM_R_X3Y104_SLICE_X3Y104_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D5 = CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D6 = CLBLM_R_X5Y104_SLICE_X6Y104_CO6;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C5 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_C6 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D1 = CLBLL_L_X2Y104_SLICE_X0Y104_CO5;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D2 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D5 = CLBLL_L_X2Y104_SLICE_X0Y104_BQ;
  assign CLBLL_L_X2Y104_SLICE_X0Y104_D6 = CLBLL_L_X2Y106_SLICE_X1Y106_BQ;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A1 = CLBLL_L_X4Y105_SLICE_X5Y105_AQ;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A2 = CLBLM_R_X5Y104_SLICE_X6Y104_CO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A5 = CLBLL_L_X4Y105_SLICE_X4Y105_AQ;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A6 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B1 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B2 = CLBLL_L_X4Y105_SLICE_X5Y105_BQ;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B3 = CLBLL_L_X4Y103_SLICE_X4Y103_BO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B4 = CLBLM_R_X5Y104_SLICE_X7Y104_BQ;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A1 = CLBLM_R_X3Y103_SLICE_X2Y103_CQ;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A2 = CLBLM_R_X3Y103_SLICE_X3Y103_CO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A3 = CLBLL_L_X2Y103_SLICE_X1Y103_AQ;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A4 = 1'b1;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A5 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C3 = CLBLM_R_X5Y104_SLICE_X6Y104_CO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C5 = CLBLL_L_X4Y105_SLICE_X5Y105_AQ;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C2 = CLBLL_L_X4Y105_SLICE_X5Y105_CQ;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_A6 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C4 = CLBLL_L_X4Y105_SLICE_X4Y105_AQ;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B1 = CLBLM_R_X3Y103_SLICE_X2Y103_CQ;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B2 = CLBLM_R_X3Y103_SLICE_X3Y103_CO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B3 = CLBLM_R_X3Y103_SLICE_X3Y103_DO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B4 = CLBLL_L_X2Y103_SLICE_X1Y103_BQ;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D1 = CLBLL_L_X4Y105_SLICE_X4Y105_AQ;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B5 = CLBLL_L_X2Y103_SLICE_X1Y103_AQ;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_B6 = CLBLM_R_X5Y104_SLICE_X6Y104_DO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C1 = CLBLL_L_X2Y103_SLICE_X1Y103_BQ;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D2 = CLBLL_L_X4Y105_SLICE_X5Y105_CQ;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C2 = CLBLM_R_X3Y103_SLICE_X3Y103_CO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D4 = CLBLL_L_X2Y105_SLICE_X0Y105_CQ;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C3 = CLBLL_L_X2Y105_SLICE_X1Y105_AO5;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D6 = CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C4 = CLBLL_L_X2Y104_SLICE_X1Y104_AO5;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_C5 = CLBLM_R_X5Y104_SLICE_X6Y104_DO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D1 = CLBLL_L_X2Y105_SLICE_X1Y105_AO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D2 = CLBLM_R_X3Y103_SLICE_X3Y103_CO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D3 = CLBLL_L_X2Y103_SLICE_X1Y103_BQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B5 = CLBLL_L_X4Y106_SLICE_X4Y106_BO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D4 = CLBLL_L_X2Y104_SLICE_X1Y104_AO5;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D5 = CLBLM_R_X5Y104_SLICE_X6Y104_DO6;
  assign CLBLL_L_X2Y104_SLICE_X1Y104_D6 = CLBLM_R_X3Y103_SLICE_X3Y103_DO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B6 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A3 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A4 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_A5 = 1'b1;
  assign CLBLM_R_X5Y107_SLICE_X7Y107_C1 = 1'b1;
  assign LIOI3_X0Y117_ILOGIC_X0Y118_D = LIOB33_X0Y117_IOB_X0Y118_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_D = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A1 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A2 = CLBLL_L_X2Y105_SLICE_X0Y105_BQ;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A3 = CLBLM_R_X3Y106_SLICE_X2Y106_BQ;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A4 = CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A5 = CLBLL_L_X4Y106_SLICE_X5Y106_AQ;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A6 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_AX = CLBLL_L_X4Y106_SLICE_X4Y106_BO5;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B1 = CLBLM_R_X3Y106_SLICE_X2Y106_CO5;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B3 = CLBLL_L_X4Y106_SLICE_X4Y106_AQ;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B4 = CLBLM_R_X3Y104_SLICE_X2Y104_DO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A1 = CLBLL_L_X2Y106_SLICE_X1Y106_A5Q;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A3 = CLBLL_L_X2Y105_SLICE_X0Y105_AQ;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A4 = CLBLL_L_X2Y103_SLICE_X1Y103_CO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A5 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B5 = CLBLL_L_X4Y106_SLICE_X5Y106_AQ;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B6 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C4 = CLBLL_L_X2Y105_SLICE_X0Y105_BQ;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B1 = CLBLM_R_X3Y105_SLICE_X2Y105_CO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B2 = CLBLL_L_X2Y105_SLICE_X0Y105_BQ;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B4 = CLBLM_R_X3Y105_SLICE_X2Y105_B5Q;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B6 = CLBLM_R_X3Y104_SLICE_X2Y104_BQ;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C3 = CLBLM_R_X3Y106_SLICE_X2Y106_AQ;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C2 = CLBLL_L_X2Y105_SLICE_X0Y105_CQ;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C3 = CLBLM_R_X3Y105_SLICE_X2Y105_CO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C4 = CLBLM_R_X3Y105_SLICE_X2Y105_B5Q;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C5 = CLBLL_L_X2Y105_SLICE_X0Y105_BQ;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D1 = CLBLL_L_X4Y106_SLICE_X4Y106_CO5;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D2 = CLBLL_L_X4Y106_SLICE_X4Y106_AQ;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D3 = CLBLL_L_X2Y106_SLICE_X1Y106_DO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D4 = CLBLL_L_X4Y106_SLICE_X4Y106_AO5;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D5 = CLBLL_L_X4Y106_SLICE_X5Y106_AQ;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D6 = CLBLM_R_X3Y106_SLICE_X2Y106_DO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D3 = CLBLL_L_X2Y105_SLICE_X0Y105_DQ;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D4 = CLBLM_R_X3Y104_SLICE_X2Y104_BQ;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D6 = CLBLL_L_X2Y105_SLICE_X1Y105_BQ;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A1 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A2 = CLBLM_R_X3Y104_SLICE_X2Y104_DO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A3 = CLBLL_L_X4Y106_SLICE_X5Y106_AQ;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A4 = CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A6 = CLBLL_L_X4Y105_SLICE_X5Y105_CQ;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B1 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B2 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B3 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B4 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A1 = CLBLM_R_X3Y106_SLICE_X3Y106_CO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A2 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A3 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A4 = CLBLM_R_X3Y105_SLICE_X2Y105_AQ;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A5 = CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A6 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C1 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C2 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B1 = CLBLL_L_X2Y105_SLICE_X1Y105_DO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B2 = CLBLL_L_X2Y104_SLICE_X1Y104_DO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B3 = CLBLL_L_X2Y106_SLICE_X0Y106_CO5;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B4 = CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B5 = CLBLL_L_X2Y104_SLICE_X1Y104_CO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B6 = CLBLL_L_X2Y105_SLICE_X1Y105_CO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C3 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C1 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D1 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C2 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C3 = CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C4 = CLBLL_L_X2Y105_SLICE_X0Y105_BQ;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C5 = CLBLL_L_X2Y105_SLICE_X0Y105_AQ;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D6 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C6 = CLBLM_R_X3Y105_SLICE_X2Y105_AQ;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D2 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D3 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D4 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D5 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D2 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D3 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D4 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D5 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D6 = CLBLL_L_X2Y105_SLICE_X0Y105_BQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C2 = CLBLM_R_X3Y107_SLICE_X2Y107_AQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C3 = CLBLL_L_X4Y107_SLICE_X5Y107_BQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C5 = CLBLL_L_X2Y107_SLICE_X1Y107_BQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D6 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A1 = CLBLL_L_X4Y107_SLICE_X4Y107_AQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A2 = CLBLL_L_X4Y107_SLICE_X4Y107_BQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A3 = CLBLM_R_X3Y106_SLICE_X2Y106_CO5;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A5 = CLBLL_L_X4Y106_SLICE_X4Y106_BO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A6 = 1'b1;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_D = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B1 = CLBLL_L_X4Y106_SLICE_X4Y106_AQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B2 = CLBLL_L_X4Y107_SLICE_X4Y107_BQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B4 = CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A1 = CLBLL_L_X2Y107_SLICE_X0Y107_CQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A2 = CLBLL_L_X2Y107_SLICE_X0Y107_BQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A3 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A4 = CLBLL_L_X2Y105_SLICE_X0Y105_BQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A5 = CLBLL_L_X2Y106_SLICE_X1Y106_AQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C1 = CLBLL_L_X4Y106_SLICE_X4Y106_BO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C2 = CLBLL_L_X4Y107_SLICE_X4Y107_CQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C3 = CLBLL_L_X4Y107_SLICE_X4Y107_AQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C5 = CLBLL_L_X4Y107_SLICE_X4Y107_BQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A6 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C6 = CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B1 = CLBLL_L_X2Y106_SLICE_X0Y106_DO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B2 = CLBLL_L_X2Y104_SLICE_X1Y104_BO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B4 = CLBLL_L_X2Y105_SLICE_X0Y105_DQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B5 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D1 = CLBLL_L_X4Y107_SLICE_X5Y107_AQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D2 = CLBLM_R_X3Y106_SLICE_X2Y106_BQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D3 = CLBLL_L_X2Y107_SLICE_X1Y107_AQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B6 = CLBLL_L_X2Y106_SLICE_X0Y106_AO5;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D5 = CLBLL_L_X4Y107_SLICE_X5Y107_BQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D4 = CLBLM_R_X3Y106_SLICE_X2Y106_AQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C2 = CLBLL_L_X2Y108_SLICE_X0Y108_BQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D6 = CLBLM_R_X3Y107_SLICE_X2Y107_AQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C3 = CLBLM_R_X3Y106_SLICE_X3Y106_DO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C4 = CLBLL_L_X2Y108_SLICE_X0Y108_A5Q;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C6 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D1 = CLBLM_R_X3Y105_SLICE_X2Y105_AQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D2 = CLBLL_L_X2Y106_SLICE_X1Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D3 = CLBLL_L_X2Y106_SLICE_X1Y106_AQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D4 = CLBLL_L_X2Y105_SLICE_X0Y105_BQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D5 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D6 = CLBLL_L_X2Y107_SLICE_X0Y107_BQ;
  assign LIOB33_X0Y119_IOB_X0Y120_O = CLBLL_L_X4Y104_SLICE_X4Y104_DO6;
  assign LIOB33_X0Y119_IOB_X0Y119_O = CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A1 = CLBLL_L_X2Y107_SLICE_X0Y107_DO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A2 = CLBLL_L_X2Y107_SLICE_X0Y107_DO5;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A4 = CLBLL_L_X4Y107_SLICE_X5Y107_AQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A6 = CLBLL_L_X2Y107_SLICE_X1Y107_CQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B1 = CLBLL_L_X2Y107_SLICE_X0Y107_DO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B2 = CLBLL_L_X2Y107_SLICE_X0Y107_DO5;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B4 = CLBLL_L_X4Y107_SLICE_X5Y107_AQ;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A1 = CLBLL_L_X2Y106_SLICE_X1Y106_AQ;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A2 = CLBLL_L_X2Y106_SLICE_X1Y106_BQ;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A4 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A6 = CLBLL_L_X2Y103_SLICE_X1Y103_CO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C1 = CLBLL_L_X2Y107_SLICE_X1Y107_CQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B5 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B6 = CLBLL_L_X4Y107_SLICE_X5Y107_BQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C4 = CLBLM_R_X3Y107_SLICE_X2Y107_BQ;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_AX = CLBLL_L_X2Y106_SLICE_X1Y106_CO5;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C6 = CLBLL_L_X4Y107_SLICE_X5Y107_AQ;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B1 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B2 = CLBLL_L_X2Y106_SLICE_X1Y106_BQ;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B3 = CLBLL_L_X4Y104_SLICE_X5Y104_AQ;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B4 = CLBLL_L_X2Y104_SLICE_X1Y104_BO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C2 = CLBLL_L_X2Y103_SLICE_X1Y103_CO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C4 = CLBLL_L_X2Y106_SLICE_X1Y106_A5Q;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C5 = CLBLL_L_X2Y106_SLICE_X1Y106_AQ;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C6 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D1 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D2 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D3 = CLBLL_L_X4Y107_SLICE_X4Y107_DO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D4 = CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D5 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D1 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D2 = CLBLL_L_X2Y105_SLICE_X0Y105_BQ;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D3 = CLBLL_L_X2Y107_SLICE_X0Y107_CQ;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D5 = CLBLL_L_X2Y106_SLICE_X1Y106_AQ;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D6 = CLBLL_L_X2Y107_SLICE_X0Y107_BQ;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = CLBLL_L_X2Y107_SLICE_X0Y107_AO5;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = CLBLL_L_X2Y105_SLICE_X1Y105_BQ;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A1 = CLBLL_L_X2Y103_SLICE_X1Y103_CO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A4 = CLBLL_L_X2Y105_SLICE_X0Y105_BQ;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A5 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A6 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B1 = CLBLL_L_X2Y107_SLICE_X0Y107_DO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B2 = CLBLL_L_X2Y107_SLICE_X0Y107_BQ;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B3 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B4 = CLBLL_L_X2Y107_SLICE_X0Y107_DO5;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B5 = CLBLM_R_X3Y105_SLICE_X2Y105_AQ;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C2 = CLBLL_L_X2Y107_SLICE_X0Y107_CQ;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C4 = CLBLL_L_X2Y107_SLICE_X0Y107_BQ;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C5 = CLBLL_L_X2Y107_SLICE_X0Y107_DO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C6 = CLBLL_L_X2Y107_SLICE_X0Y107_DO5;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D2 = CLBLL_L_X2Y103_SLICE_X1Y103_CO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D4 = CLBLL_L_X2Y105_SLICE_X0Y105_CQ;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D6 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A2 = CLBLM_R_X3Y106_SLICE_X2Y106_AO5;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A3 = CLBLL_L_X2Y107_SLICE_X1Y107_AQ;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A4 = CLBLL_L_X2Y107_SLICE_X1Y107_DO5;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A6 = CLBLL_L_X2Y107_SLICE_X1Y107_BQ;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B1 = CLBLL_L_X2Y107_SLICE_X1Y107_DO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B2 = CLBLM_R_X3Y106_SLICE_X2Y106_AO5;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B3 = CLBLM_R_X3Y106_SLICE_X2Y106_AQ;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B6 = CLBLL_L_X2Y107_SLICE_X1Y107_BQ;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C2 = CLBLM_R_X3Y106_SLICE_X2Y106_AO5;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C3 = CLBLL_L_X2Y107_SLICE_X1Y107_BQ;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C4 = CLBLL_L_X2Y107_SLICE_X1Y107_AQ;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C5 = CLBLL_L_X2Y107_SLICE_X1Y107_DO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C6 = CLBLL_L_X2Y107_SLICE_X1Y107_CQ;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D1 = CLBLL_L_X2Y105_SLICE_X0Y105_BQ;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D2 = CLBLL_L_X2Y103_SLICE_X1Y103_CO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D3 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D6 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B6 = CLBLM_R_X3Y105_SLICE_X2Y105_BQ;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C3 = CLBLM_R_X5Y105_SLICE_X6Y105_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D3 = CLBLM_R_X3Y107_SLICE_X3Y107_AO5;
  assign CLBLL_L_X2Y103_SLICE_X0Y103_A4 = CLBLL_L_X2Y106_SLICE_X1Y106_BQ;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A1 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A2 = CLBLM_R_X3Y104_SLICE_X2Y104_CO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A4 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_AX = CLBLL_L_X2Y108_SLICE_X0Y108_BO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B1 = CLBLL_L_X2Y108_SLICE_X0Y108_A5Q;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B2 = CLBLM_R_X3Y104_SLICE_X2Y104_CO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B3 = CLBLL_L_X2Y108_SLICE_X0Y108_AQ;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B5 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_BX = CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C3 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D1 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D3 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A1 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A3 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B1 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B3 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C1 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C3 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D1 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D3 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D6 = 1'b1;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_D = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A2 = CLBLM_R_X3Y104_SLICE_X3Y104_AQ;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A3 = CLBLM_R_X3Y103_SLICE_X3Y103_AQ;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A4 = CLBLL_L_X2Y105_SLICE_X0Y105_CQ;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A5 = CLBLM_R_X5Y103_SLICE_X7Y103_AO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_A6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_D = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B1 = CLBLL_L_X4Y105_SLICE_X5Y105_DO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B2 = CLBLM_R_X3Y103_SLICE_X3Y103_BQ;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B3 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_B6 = CLBLM_R_X3Y105_SLICE_X2Y105_A5Q;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C1 = CLBLL_L_X4Y105_SLICE_X5Y105_BQ;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C2 = CLBLL_L_X2Y105_SLICE_X0Y105_BQ;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C3 = CLBLL_L_X4Y103_SLICE_X4Y103_CO6;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C4 = CLBLL_L_X4Y104_SLICE_X5Y104_AO5;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C5 = CLBLL_L_X2Y105_SLICE_X0Y105_CQ;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_C6 = CLBLL_L_X4Y104_SLICE_X4Y104_BQ;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D1 = CLBLL_L_X4Y103_SLICE_X4Y103_AQ;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D2 = CLBLM_R_X5Y105_SLICE_X7Y105_AQ;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D3 = CLBLM_R_X3Y105_SLICE_X3Y105_AQ;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D4 = CLBLM_R_X3Y105_SLICE_X2Y105_A5Q;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D5 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X3Y103_D6 = CLBLL_L_X2Y105_SLICE_X1Y105_CO6;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A2 = CLBLM_R_X5Y103_SLICE_X7Y103_AO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A3 = CLBLM_R_X3Y103_SLICE_X2Y103_AQ;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A5 = CLBLM_R_X3Y103_SLICE_X3Y103_AQ;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_A6 = CLBLL_L_X2Y105_SLICE_X0Y105_CQ;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B1 = CLBLM_R_X3Y103_SLICE_X2Y103_BQ;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B2 = CLBLM_R_X5Y103_SLICE_X7Y103_AO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B3 = CLBLM_R_X3Y103_SLICE_X2Y103_AQ;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_B6 = CLBLL_L_X2Y105_SLICE_X0Y105_CQ;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C1 = CLBLL_L_X2Y105_SLICE_X0Y105_AQ;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C2 = CLBLM_R_X3Y103_SLICE_X3Y103_CO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C4 = CLBLL_L_X2Y103_SLICE_X1Y103_CO6;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C5 = CLBLM_R_X3Y103_SLICE_X2Y103_CQ;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_C6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D1 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D2 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D3 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D4 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D5 = 1'b1;
  assign CLBLM_R_X3Y103_SLICE_X2Y103_D6 = 1'b1;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_D = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = CLBLL_L_X2Y106_SLICE_X0Y106_BQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = CLBLL_L_X2Y106_SLICE_X0Y106_BQ;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D3 = CLBLM_R_X3Y105_SLICE_X3Y105_AQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D5 = CLBLL_L_X4Y105_SLICE_X5Y105_AQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = CLBLL_L_X4Y104_SLICE_X4Y104_DO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A1 = CLBLL_L_X4Y107_SLICE_X4Y107_CQ;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A3 = CLBLM_R_X3Y104_SLICE_X3Y104_AQ;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A6 = CLBLM_R_X5Y104_SLICE_X7Y104_CO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B2 = CLBLM_R_X3Y104_SLICE_X3Y104_BQ;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B3 = CLBLM_R_X3Y103_SLICE_X2Y103_BQ;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B4 = CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B6 = CLBLL_L_X4Y104_SLICE_X4Y104_BQ;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C1 = CLBLM_R_X3Y104_SLICE_X2Y104_AQ;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C2 = CLBLL_L_X2Y105_SLICE_X0Y105_BQ;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C3 = CLBLL_L_X2Y104_SLICE_X0Y104_AQ;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C4 = CLBLL_L_X4Y105_SLICE_X5Y105_CQ;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C5 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C6 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D1 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D2 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D3 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D4 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D5 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A3 = CLBLM_R_X3Y104_SLICE_X2Y104_AQ;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A4 = CLBLM_R_X3Y105_SLICE_X2Y105_BQ;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A6 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B2 = CLBLM_R_X3Y104_SLICE_X2Y104_BQ;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B3 = CLBLM_R_X3Y104_SLICE_X2Y104_AQ;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B4 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C1 = CLBLM_R_X3Y104_SLICE_X3Y104_AQ;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C2 = CLBLM_R_X3Y103_SLICE_X2Y103_AQ;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C3 = CLBLL_L_X2Y108_SLICE_X0Y108_AQ;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C4 = CLBLM_R_X3Y103_SLICE_X2Y103_BQ;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C5 = CLBLM_R_X3Y103_SLICE_X3Y103_AQ;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C6 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D1 = CLBLM_R_X3Y104_SLICE_X3Y104_AQ;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D2 = CLBLM_R_X3Y103_SLICE_X2Y103_AQ;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D3 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D4 = CLBLL_L_X2Y108_SLICE_X0Y108_BO5;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D5 = CLBLM_R_X3Y103_SLICE_X3Y103_AQ;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D6 = CLBLM_R_X3Y103_SLICE_X2Y103_BQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A1 = CLBLL_L_X2Y105_SLICE_X0Y105_CQ;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A3 = CLBLM_R_X3Y105_SLICE_X2Y105_CO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A4 = CLBLM_R_X3Y105_SLICE_X2Y105_B5Q;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A5 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A6 = CLBLM_R_X3Y105_SLICE_X3Y105_AQ;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B1 = CLBLL_L_X2Y105_SLICE_X0Y105_CQ;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B2 = CLBLL_L_X2Y105_SLICE_X1Y105_CO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B3 = CLBLM_R_X3Y105_SLICE_X2Y105_A5Q;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B4 = CLBLL_L_X4Y104_SLICE_X5Y104_AQ;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B5 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B6 = CLBLL_L_X4Y105_SLICE_X5Y105_BQ;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C1 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C4 = CLBLL_L_X2Y105_SLICE_X0Y105_BQ;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C5 = CLBLM_R_X3Y105_SLICE_X3Y105_AQ;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C6 = CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D1 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D2 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D3 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D4 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D5 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D6 = 1'b1;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_D = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A1 = CLBLM_R_X3Y105_SLICE_X2Y105_DO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A2 = CLBLL_L_X2Y104_SLICE_X1Y104_BO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A3 = CLBLM_R_X3Y105_SLICE_X2Y105_AQ;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A4 = CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A5 = CLBLL_L_X2Y107_SLICE_X1Y107_DO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A6 = CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_AX = CLBLM_R_X3Y105_SLICE_X2Y105_CO5;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B2 = CLBLM_R_X3Y105_SLICE_X2Y105_BQ;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B4 = CLBLL_L_X2Y105_SLICE_X0Y105_DQ;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B5 = CLBLM_R_X3Y105_SLICE_X2Y105_B5Q;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_BX = CLBLM_R_X3Y105_SLICE_X2Y105_DO5;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C1 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C3 = CLBLM_R_X5Y105_SLICE_X7Y105_AQ;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C4 = CLBLM_R_X3Y105_SLICE_X2Y105_A5Q;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C6 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_C4 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D1 = CLBLM_R_X3Y107_SLICE_X2Y107_AQ;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_C5 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D4 = CLBLL_L_X2Y107_SLICE_X0Y107_CQ;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D6 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_C6 = 1'b1;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_D = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_D = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_D1 = 1'b1;
  assign CLBLM_R_X5Y103_SLICE_X7Y103_D6 = 1'b1;
endmodule
