module top(
  input LIOB33_SING_X0Y100_IOB_X0Y100_IPAD,
  input LIOB33_X0Y101_IOB_X0Y101_IPAD,
  input LIOB33_X0Y101_IOB_X0Y102_IPAD,
  input LIOB33_X0Y103_IOB_X0Y103_IPAD,
  input LIOB33_X0Y103_IOB_X0Y104_IPAD,
  input LIOB33_X0Y105_IOB_X0Y105_IPAD,
  input LIOB33_X0Y105_IOB_X0Y106_IPAD,
  input LIOB33_X0Y107_IOB_X0Y107_IPAD,
  input LIOB33_X0Y107_IOB_X0Y108_IPAD,
  input LIOB33_X0Y109_IOB_X0Y109_IPAD,
  input LIOB33_X0Y109_IOB_X0Y110_IPAD,
  input LIOB33_X0Y111_IOB_X0Y111_IPAD,
  input LIOB33_X0Y111_IOB_X0Y112_IPAD,
  input LIOB33_X0Y113_IOB_X0Y113_IPAD,
  input LIOB33_X0Y113_IOB_X0Y114_IPAD,
  input LIOB33_X0Y115_IOB_X0Y115_IPAD,
  input LIOB33_X0Y115_IOB_X0Y116_IPAD,
  input LIOB33_X0Y117_IOB_X0Y117_IPAD,
  input LIOB33_X0Y117_IOB_X0Y118_IPAD,
  input LIOB33_X0Y127_IOB_X0Y128_IPAD,
  output LIOB33_X0Y119_IOB_X0Y119_OPAD,
  output LIOB33_X0Y119_IOB_X0Y120_OPAD,
  output LIOB33_X0Y121_IOB_X0Y121_OPAD,
  output LIOB33_X0Y121_IOB_X0Y122_OPAD,
  output LIOB33_X0Y123_IOB_X0Y123_OPAD,
  output LIOB33_X0Y123_IOB_X0Y124_OPAD
  );
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_AO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_AO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_A_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_BO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_BO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_B_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_CO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_CO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_C_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_DO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_DO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X0Y105_D_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_AO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_AO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_AQ;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_A_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_BO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_BO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_B_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_CLK;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_CO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_CO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_C_XOR;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D1;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D2;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D3;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D4;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_DO5;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_DO6;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D_CY;
  wire [0:0] CLBLL_L_X2Y105_SLICE_X1Y105_D_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_AO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_AQ;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_A_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_BO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_BQ;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_B_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_CLK;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_CO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_CQ;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_C_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_DO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_DO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_DQ;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X0Y106_D_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A5Q;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_AMUX;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_AO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_AQ;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_AX;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_A_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_BO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_BQ;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_B_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_CLK;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_CMUX;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_CO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_CO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_C_XOR;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D1;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D2;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D3;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D4;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_DO5;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_DO6;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D_CY;
  wire [0:0] CLBLL_L_X2Y106_SLICE_X1Y106_D_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_AO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_AQ;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_A_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_BO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_BO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_B_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_CLK;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_CO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_CO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_C_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_DO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_DO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X0Y107_D_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_AO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_AQ;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_A_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_BO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_BO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_BQ;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_B_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_CLK;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_CO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_CO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_CQ;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_C_XOR;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D1;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D2;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D3;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D4;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_DO5;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_DO6;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_DQ;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D_CY;
  wire [0:0] CLBLL_L_X2Y107_SLICE_X1Y107_D_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_AO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_A_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_BO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_BO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_B_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_CO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_C_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_DO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_DO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X0Y108_D_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_AMUX;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_AO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_A_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_BMUX;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_BO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_B_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_CO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_CO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_C_XOR;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D1;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D2;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D3;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D4;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_DMUX;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_DO5;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D_CY;
  wire [0:0] CLBLL_L_X2Y108_SLICE_X1Y108_D_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_AO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_AQ;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_A_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_BMUX;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_BO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_B_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_CLK;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_CO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_C_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_DO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_DO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X0Y109_D_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_AO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_AO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_AQ;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_A_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_BO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_BO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_BQ;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_B_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_CLK;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_CMUX;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_CO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_CO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_C_XOR;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D1;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D2;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D3;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D4;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_DMUX;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_DO5;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_DO6;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D_CY;
  wire [0:0] CLBLL_L_X2Y109_SLICE_X1Y109_D_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_AO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_AQ;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_A_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_BO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_BO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_BQ;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_B_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_CLK;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_CO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_CO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_CQ;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_C_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_DO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_DO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X0Y110_D_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_AO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_AO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_AQ;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_A_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_BO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_BO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_B_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_CLK;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_CO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_CO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_C_XOR;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D1;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D2;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D3;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D4;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_DO5;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D_CY;
  wire [0:0] CLBLL_L_X2Y110_SLICE_X1Y110_D_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_AO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_AO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_AQ;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_A_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_BO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_BO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_BQ;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_B_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_CLK;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_CO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_C_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_DO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_DO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X4Y104_D_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_AO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_AO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_AQ;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_A_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_BO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_BO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_BQ;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_B_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_CLK;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_CO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_CO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_C_XOR;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D1;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D2;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D3;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D4;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_DO5;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_DO6;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D_CY;
  wire [0:0] CLBLL_L_X4Y104_SLICE_X5Y104_D_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_AO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_AO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_AQ;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_A_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_BO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_BO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_BQ;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_B_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_CLK;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_CO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_CQ;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_C_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_DO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_DO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_DQ;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X4Y105_D_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_AO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_AO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_AQ;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_A_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_BO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_B_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_CLK;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_CO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_CO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_C_XOR;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D1;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D2;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D3;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D4;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_DO5;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_DO6;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D_CY;
  wire [0:0] CLBLL_L_X4Y105_SLICE_X5Y105_D_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_AO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_AO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_AQ;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_A_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_BO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_BO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_BQ;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_B_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_CLK;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_CO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_CQ;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_C_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_DO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_DO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X4Y106_D_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_AO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_AO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_AQ;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_A_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_BO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_BO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_BQ;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_B_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_CLK;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_CO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_CO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_C_XOR;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D1;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D2;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D3;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D4;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_DO5;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_DO6;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D_CY;
  wire [0:0] CLBLL_L_X4Y106_SLICE_X5Y106_D_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_AO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_AQ;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_A_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B5Q;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_BMUX;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_BO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_BQ;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_B_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_CLK;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_CO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_C_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_DO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_DO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X4Y107_D_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A5Q;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_AMUX;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_AO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_AO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_AQ;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_AX;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_A_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_BMUX;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_BO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_B_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_CLK;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_CMUX;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_CO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_C_XOR;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D1;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D2;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D3;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D4;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_DO5;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D_CY;
  wire [0:0] CLBLL_L_X4Y107_SLICE_X5Y107_D_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_A_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_BO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_B_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_CO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_C_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_DO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X4Y108_D_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_AO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_A_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_BO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_B_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_CO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_C_XOR;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D1;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D2;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D3;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D4;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_DO5;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_DO6;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D_CY;
  wire [0:0] CLBLL_L_X4Y108_SLICE_X5Y108_D_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A5Q;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AMUX;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_AX;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_A_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_BQ;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_B_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CLK;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CMUX;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_C_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_DMUX;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_DO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X4Y109_D_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_A_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_BO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_BQ;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_B_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CLK;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_C_XOR;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D1;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D2;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D3;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D4;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_DO5;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D_CY;
  wire [0:0] CLBLL_L_X4Y109_SLICE_X5Y109_D_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_AO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_AO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_AQ;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_A_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_BO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_BO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_BQ;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_B_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_CLK;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_CO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_CO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_CQ;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_C_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_DO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_DO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_DQ;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X2Y104_D_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_AO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_AO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_AQ;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_A_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_BO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_BQ;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_B_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_CLK;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_CO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_CO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_C_XOR;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D1;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D2;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D3;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D4;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_DO5;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_DO6;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D_CY;
  wire [0:0] CLBLM_R_X3Y104_SLICE_X3Y104_D_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_AO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_AQ;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_A_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_BO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_BO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_BQ;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_B_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_CLK;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_CMUX;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_CO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_CO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_C_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_DMUX;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_DO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_DO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X2Y105_D_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A5Q;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_AMUX;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_AO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_AO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_AQ;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_AX;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_A_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_BMUX;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_BO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_B_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_CLK;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_CO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_C_XOR;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D1;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D2;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D3;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D4;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_DO5;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_DO6;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D_CY;
  wire [0:0] CLBLM_R_X3Y105_SLICE_X3Y105_D_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_AO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_AO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_AQ;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_A_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_BO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_BO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_B_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_CLK;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_CMUX;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_CO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_C_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_DO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_DO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X2Y106_D_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_AO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_AO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_A_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_BO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_B_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_CO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_CO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_C_XOR;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D1;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D2;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D3;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D4;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_DO5;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_DO6;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D_CY;
  wire [0:0] CLBLM_R_X3Y106_SLICE_X3Y106_D_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_AO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_AQ;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_A_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_BO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_BO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_B_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_CLK;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_CO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_C_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_DO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_DO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X2Y107_D_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_AO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_AO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_A_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_BO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_BO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_B_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_CO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_C_XOR;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D1;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D2;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D3;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D4;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_DO5;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_DO6;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D_CY;
  wire [0:0] CLBLM_R_X3Y107_SLICE_X3Y107_D_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_AO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_AO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_AQ;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_A_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_BO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_BO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_BQ;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_B_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_CLK;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_CMUX;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_CO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_CO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_C_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_DO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X2Y108_D_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_AMUX;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_AO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_A_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_BMUX;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_BO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_B_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_CMUX;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_CO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_C_XOR;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D1;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D2;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D3;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D4;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_DO5;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D_CY;
  wire [0:0] CLBLM_R_X3Y108_SLICE_X3Y108_D_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_AQ;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_A_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B5Q;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_BMUX;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_BO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_BO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_BQ;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_B_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CLK;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CMUX;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_C_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_DO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_DO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X2Y109_D_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AMUX;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_A_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_BO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_BQ;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_B_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CLK;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_C_XOR;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D1;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D2;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D3;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D4;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_DO5;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D_CY;
  wire [0:0] CLBLM_R_X3Y109_SLICE_X3Y109_D_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A5Q;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AMUX;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AQ;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_AX;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_A_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_BO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_BQ;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_B_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_CLK;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_CO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_CQ;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_C_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_DMUX;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_DO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X2Y110_D_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A5Q;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AMUX;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_AQ;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_A_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_BO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_B_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_CLK;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_CMUX;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_CO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_C_XOR;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D1;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D2;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D3;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D4;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_DO5;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D_CY;
  wire [0:0] CLBLM_R_X3Y110_SLICE_X3Y110_D_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_AO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_AQ;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_A_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_BO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_BO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_BQ;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_B_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_CLK;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_CO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_CO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_CQ;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_C_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_DO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_DO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X6Y105_D_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A5Q;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_AMUX;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_AO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_AO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_AQ;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_AX;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_A_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_BMUX;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_BO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_BO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_B_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_CLK;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_CO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_C_XOR;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D1;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D2;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D3;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D4;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_DO5;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_DO6;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D_CY;
  wire [0:0] CLBLM_R_X5Y105_SLICE_X7Y105_D_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A5Q;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_AMUX;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_AO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_AQ;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_A_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B5Q;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_BMUX;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_BO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_BQ;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_B_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_CLK;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_CO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_CQ;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_C_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_DMUX;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_DO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X6Y106_D_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_AO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_AO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_A_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_BO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_B_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_CO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_CO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_C_XOR;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D1;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D2;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D3;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D4;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_DO5;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_DO6;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D_CY;
  wire [0:0] CLBLM_R_X5Y106_SLICE_X7Y106_D_XOR;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I;
  wire [0:0] CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  wire [0:0] LIOB33_SING_X0Y100_IOB_X0Y100_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y101_I;
  wire [0:0] LIOB33_X0Y101_IOB_X0Y102_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y103_I;
  wire [0:0] LIOB33_X0Y103_IOB_X0Y104_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y105_I;
  wire [0:0] LIOB33_X0Y105_IOB_X0Y106_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y107_I;
  wire [0:0] LIOB33_X0Y107_IOB_X0Y108_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y109_I;
  wire [0:0] LIOB33_X0Y109_IOB_X0Y110_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_I;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y113_I;
  wire [0:0] LIOB33_X0Y113_IOB_X0Y114_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y115_I;
  wire [0:0] LIOB33_X0Y115_IOB_X0Y116_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y117_I;
  wire [0:0] LIOB33_X0Y117_IOB_X0Y118_I;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y119_O;
  wire [0:0] LIOB33_X0Y119_IOB_X0Y120_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y121_O;
  wire [0:0] LIOB33_X0Y121_IOB_X0Y122_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y123_O;
  wire [0:0] LIOB33_X0Y123_IOB_X0Y124_O;
  wire [0:0] LIOB33_X0Y127_IOB_X0Y128_I;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_D;
  wire [0:0] LIOI3_SING_X0Y100_ILOGIC_X0Y100_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y101_O;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_D;
  wire [0:0] LIOI3_X0Y101_ILOGIC_X0Y102_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y103_O;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_D;
  wire [0:0] LIOI3_X0Y103_ILOGIC_X0Y104_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y105_O;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_D;
  wire [0:0] LIOI3_X0Y105_ILOGIC_X0Y106_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y109_O;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_D;
  wire [0:0] LIOI3_X0Y109_ILOGIC_X0Y110_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y111_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y115_O;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_D;
  wire [0:0] LIOI3_X0Y115_ILOGIC_X0Y116_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y117_O;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y118_D;
  wire [0:0] LIOI3_X0Y117_ILOGIC_X0Y118_O;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y121_TQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_D1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_OQ;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_T1;
  wire [0:0] LIOI3_X0Y121_OLOGIC_X0Y122_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y123_TQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_D1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_OQ;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_T1;
  wire [0:0] LIOI3_X0Y123_OLOGIC_X0Y124_TQ;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_D;
  wire [0:0] LIOI3_X0Y127_ILOGIC_X0Y128_O;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y105_SLICE_X0Y105_DO5),
.O6(CLBLL_L_X2Y105_SLICE_X0Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y105_SLICE_X0Y105_CO5),
.O6(CLBLL_L_X2Y105_SLICE_X0Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y105_SLICE_X0Y105_BO5),
.O6(CLBLL_L_X2Y105_SLICE_X0Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y105_SLICE_X0Y105_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y105_SLICE_X0Y105_AO5),
.O6(CLBLL_L_X2Y105_SLICE_X0Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y105_SLICE_X1Y105_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y105_SLICE_X1Y105_AO6),
.Q(CLBLL_L_X2Y105_SLICE_X1Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y105_SLICE_X1Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y105_SLICE_X1Y105_DO5),
.O6(CLBLL_L_X2Y105_SLICE_X1Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y105_SLICE_X1Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y105_SLICE_X1Y105_CO5),
.O6(CLBLL_L_X2Y105_SLICE_X1Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y105_SLICE_X1Y105_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y105_SLICE_X1Y105_BO5),
.O6(CLBLL_L_X2Y105_SLICE_X1Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaaf5005aaaa0000)
  ) CLBLL_L_X2Y105_SLICE_X1Y105_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(1'b1),
.I2(CLBLL_L_X2Y105_SLICE_X1Y105_AQ),
.I3(CLBLM_R_X3Y105_SLICE_X2Y105_CO5),
.I4(CLBLM_R_X3Y104_SLICE_X2Y104_BQ),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLL_L_X2Y105_SLICE_X1Y105_AO5),
.O6(CLBLL_L_X2Y105_SLICE_X1Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y106_SLICE_X0Y106_AO6),
.Q(CLBLL_L_X2Y106_SLICE_X0Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y106_SLICE_X0Y106_BO6),
.Q(CLBLL_L_X2Y106_SLICE_X0Y106_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y106_SLICE_X0Y106_CO6),
.Q(CLBLL_L_X2Y106_SLICE_X0Y106_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y106_SLICE_X0Y106_DO6),
.Q(CLBLL_L_X2Y106_SLICE_X0Y106_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h99d8dddd8888dddd)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_DLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLL_L_X2Y106_SLICE_X0Y106_CQ),
.I2(CLBLL_L_X2Y106_SLICE_X0Y106_DQ),
.I3(LIOB33_X0Y101_IOB_X0Y102_I),
.I4(CLBLL_L_X2Y106_SLICE_X1Y106_CO6),
.I5(CLBLL_L_X2Y107_SLICE_X0Y107_AQ),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_DO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdf0ffff0d000f0f)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_CLUT (
.I0(CLBLL_L_X2Y106_SLICE_X0Y106_CQ),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLL_L_X2Y107_SLICE_X0Y107_AQ),
.I4(CLBLL_L_X2Y106_SLICE_X1Y106_CO6),
.I5(CLBLL_L_X2Y106_SLICE_X0Y106_AQ),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_CO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f7f0d5f055f055)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_BLUT (
.I0(CLBLL_L_X2Y106_SLICE_X1Y106_CO6),
.I1(LIOB33_X0Y101_IOB_X0Y102_I),
.I2(CLBLL_L_X2Y106_SLICE_X0Y106_DQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLL_L_X2Y106_SLICE_X0Y106_BQ),
.I5(CLBLL_L_X2Y107_SLICE_X0Y107_AQ),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_BO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00cc00cc00fc30)
  ) CLBLL_L_X2Y106_SLICE_X0Y106_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLL_L_X2Y106_SLICE_X0Y106_AQ),
.I3(CLBLL_L_X2Y106_SLICE_X1Y106_BQ),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLL_L_X2Y106_SLICE_X0Y106_AO5),
.O6(CLBLL_L_X2Y106_SLICE_X0Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y106_SLICE_X1Y106_CO5),
.Q(CLBLL_L_X2Y106_SLICE_X1Y106_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y106_SLICE_X1Y106_AO6),
.Q(CLBLL_L_X2Y106_SLICE_X1Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y106_SLICE_X1Y106_BO6),
.Q(CLBLL_L_X2Y106_SLICE_X1Y106_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f0fcc00cf0f)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y105_SLICE_X5Y105_DO6),
.I2(CLBLL_L_X4Y106_SLICE_X4Y106_DO6),
.I3(CLBLL_L_X2Y106_SLICE_X1Y106_AQ),
.I4(CLBLL_L_X2Y107_SLICE_X1Y107_DQ),
.I5(CLBLL_L_X4Y105_SLICE_X4Y105_AQ),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_DO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c0aaaa000f)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_CLUT (
.I0(CLBLL_L_X4Y105_SLICE_X4Y105_AQ),
.I1(LIOB33_X0Y105_IOB_X0Y105_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLL_L_X2Y106_SLICE_X1Y106_A5Q),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_CO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaa0aaa0aa0caa0c)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_BLUT (
.I0(CLBLL_L_X2Y106_SLICE_X1Y106_AQ),
.I1(CLBLL_L_X2Y106_SLICE_X1Y106_BQ),
.I2(LIOB33_X0Y103_IOB_X0Y103_I),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(1'b1),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_BO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc55cc00cc00ccf0)
  ) CLBLL_L_X2Y106_SLICE_X1Y106_ALUT (
.I0(CLBLL_L_X2Y107_SLICE_X1Y107_DQ),
.I1(CLBLL_L_X2Y107_SLICE_X0Y107_AQ),
.I2(CLBLL_L_X2Y106_SLICE_X1Y106_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y103_IOB_X0Y103_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLL_L_X2Y106_SLICE_X1Y106_AO5),
.O6(CLBLL_L_X2Y106_SLICE_X1Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y107_SLICE_X0Y107_AO6),
.Q(CLBLL_L_X2Y107_SLICE_X0Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_DO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_CO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_BO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hee22ee22cc00cc00)
  ) CLBLL_L_X2Y107_SLICE_X0Y107_ALUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(1'b1),
.I3(CLBLL_L_X2Y107_SLICE_X1Y107_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y105_IOB_X0Y105_I),
.O5(CLBLL_L_X2Y107_SLICE_X0Y107_AO5),
.O6(CLBLL_L_X2Y107_SLICE_X0Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y107_SLICE_X1Y107_AO6),
.Q(CLBLL_L_X2Y107_SLICE_X1Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y107_SLICE_X1Y107_BO6),
.Q(CLBLL_L_X2Y107_SLICE_X1Y107_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y107_SLICE_X1Y107_CO6),
.Q(CLBLL_L_X2Y107_SLICE_X1Y107_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y107_SLICE_X1Y107_DO6),
.Q(CLBLL_L_X2Y107_SLICE_X1Y107_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000044304430)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_DLUT (
.I0(CLBLL_L_X2Y106_SLICE_X0Y106_AQ),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(CLBLL_L_X2Y107_SLICE_X1Y107_DQ),
.I3(LIOB33_X0Y103_IOB_X0Y103_I),
.I4(CLBLM_R_X3Y109_SLICE_X2Y109_B5Q),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_DO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0faf0f000aa0000)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_CLUT (
.I0(CLBLM_R_X3Y107_SLICE_X2Y107_BO6),
.I1(1'b1),
.I2(CLBLL_L_X2Y107_SLICE_X1Y107_DQ),
.I3(CLBLM_R_X3Y106_SLICE_X3Y106_DO6),
.I4(CLBLL_L_X2Y108_SLICE_X1Y108_BO5),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_CO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfeeefaaafcccf000)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_BLUT (
.I0(LIOB33_X0Y103_IOB_X0Y103_I),
.I1(CLBLL_L_X2Y107_SLICE_X1Y107_BQ),
.I2(CLBLL_L_X2Y107_SLICE_X1Y107_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLL_L_X2Y108_SLICE_X1Y108_AO6),
.I5(CLBLL_L_X2Y108_SLICE_X1Y108_AO5),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_BO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefaeeaafcf0cc00)
  ) CLBLL_L_X2Y107_SLICE_X1Y107_ALUT (
.I0(LIOB33_X0Y101_IOB_X0Y102_I),
.I1(CLBLL_L_X2Y109_SLICE_X1Y109_BQ),
.I2(CLBLL_L_X2Y107_SLICE_X1Y107_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLL_L_X2Y108_SLICE_X1Y108_AO6),
.I5(CLBLL_L_X2Y108_SLICE_X1Y108_AO5),
.O5(CLBLL_L_X2Y107_SLICE_X1Y107_AO5),
.O6(CLBLL_L_X2Y107_SLICE_X1Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_DO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_CO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_BO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y108_SLICE_X0Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X0Y108_AO5),
.O6(CLBLL_L_X2Y108_SLICE_X0Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf1f10101f1fd010d)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_DLUT (
.I0(CLBLL_L_X2Y107_SLICE_X1Y107_AQ),
.I1(CLBLM_R_X3Y108_SLICE_X2Y108_BQ),
.I2(CLBLL_L_X2Y106_SLICE_X0Y106_CQ),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(LIOB33_X0Y101_IOB_X0Y101_I),
.I5(CLBLL_L_X2Y107_SLICE_X1Y107_BQ),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_DO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0e0e00000e020000)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_CLUT (
.I0(CLBLL_L_X2Y107_SLICE_X1Y107_AQ),
.I1(CLBLM_R_X3Y108_SLICE_X2Y108_BQ),
.I2(CLBLL_L_X2Y106_SLICE_X0Y106_CQ),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(CLBLM_R_X3Y109_SLICE_X3Y109_CQ),
.I5(CLBLL_L_X2Y107_SLICE_X1Y107_BQ),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_CO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000fad8ccccffdd)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_BLUT (
.I0(CLBLM_R_X3Y108_SLICE_X2Y108_BQ),
.I1(CLBLL_L_X2Y107_SLICE_X1Y107_BQ),
.I2(CLBLL_L_X2Y107_SLICE_X1Y107_AQ),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(CLBLL_L_X2Y106_SLICE_X0Y106_CQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_BO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h1030103023032303)
  ) CLBLL_L_X2Y108_SLICE_X1Y108_ALUT (
.I0(CLBLL_L_X2Y106_SLICE_X0Y106_DQ),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLL_L_X4Y108_SLICE_X4Y108_AO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y108_SLICE_X1Y108_AO5),
.O6(CLBLL_L_X2Y108_SLICE_X1Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y109_SLICE_X0Y109_AO6),
.Q(CLBLL_L_X2Y109_SLICE_X0Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_DO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_CO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f00030f0f0005)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_BLUT (
.I0(LIOB33_X0Y115_IOB_X0Y116_I),
.I1(LIOB33_X0Y113_IOB_X0Y114_I),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLL_L_X4Y108_SLICE_X4Y108_AO6),
.I4(CLBLL_L_X2Y106_SLICE_X0Y106_CQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_BO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa0ffa082a082a0)
  ) CLBLL_L_X2Y109_SLICE_X0Y109_ALUT (
.I0(CLBLL_L_X2Y109_SLICE_X0Y109_BO5),
.I1(CLBLM_R_X3Y107_SLICE_X2Y107_CO6),
.I2(CLBLL_L_X2Y109_SLICE_X0Y109_AQ),
.I3(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I4(1'b1),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLL_L_X2Y109_SLICE_X0Y109_AO5),
.O6(CLBLL_L_X2Y109_SLICE_X0Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y109_SLICE_X1Y109_AO6),
.Q(CLBLL_L_X2Y109_SLICE_X1Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y109_SLICE_X1Y109_BO6),
.Q(CLBLL_L_X2Y109_SLICE_X1Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h8f8f8888ff000000)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_DLUT (
.I0(CLBLL_L_X2Y108_SLICE_X1Y108_BO6),
.I1(CLBLL_L_X2Y109_SLICE_X1Y109_AQ),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(CLBLL_L_X4Y108_SLICE_X4Y108_AO6),
.I4(CLBLL_L_X2Y106_SLICE_X0Y106_CQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_DO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h708f7788008f0088)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_CLUT (
.I0(CLBLL_L_X2Y108_SLICE_X1Y108_BO6),
.I1(CLBLL_L_X2Y109_SLICE_X1Y109_AQ),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(CLBLM_R_X3Y110_SLICE_X2Y110_CQ),
.I4(CLBLL_L_X2Y106_SLICE_X0Y106_CQ),
.I5(1'b1),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_CO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff4f004f004f00)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_BLUT (
.I0(CLBLM_R_X3Y106_SLICE_X2Y106_CO6),
.I1(CLBLL_L_X2Y109_SLICE_X1Y109_BQ),
.I2(CLBLM_R_X3Y106_SLICE_X3Y106_BO6),
.I3(CLBLL_L_X2Y109_SLICE_X0Y109_BO5),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLL_L_X2Y110_SLICE_X0Y110_CQ),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_BO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfabef0f0aaaa0000)
  ) CLBLL_L_X2Y109_SLICE_X1Y109_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I2(CLBLL_L_X2Y109_SLICE_X1Y109_AQ),
.I3(CLBLM_R_X3Y107_SLICE_X2Y107_CO6),
.I4(CLBLL_L_X2Y109_SLICE_X0Y109_AQ),
.I5(CLBLL_L_X2Y109_SLICE_X0Y109_BO5),
.O5(CLBLL_L_X2Y109_SLICE_X1Y109_AO5),
.O6(CLBLL_L_X2Y109_SLICE_X1Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y110_SLICE_X0Y110_AO6),
.Q(CLBLL_L_X2Y110_SLICE_X0Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y110_SLICE_X0Y110_BO6),
.Q(CLBLL_L_X2Y110_SLICE_X0Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y110_SLICE_X0Y110_CO6),
.Q(CLBLL_L_X2Y110_SLICE_X0Y110_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0f0f0f0f0f)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_DO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff888f888f888)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_CLUT (
.I0(CLBLL_L_X2Y108_SLICE_X1Y108_AO6),
.I1(CLBLL_L_X2Y110_SLICE_X0Y110_CQ),
.I2(CLBLL_L_X2Y110_SLICE_X0Y110_BQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y115_IOB_X0Y116_I),
.I5(CLBLL_L_X2Y108_SLICE_X1Y108_AO5),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_CO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffeca0eca0eca0)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_BLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(LIOB33_X0Y115_IOB_X0Y115_I),
.I2(CLBLL_L_X2Y110_SLICE_X0Y110_AQ),
.I3(CLBLL_L_X2Y108_SLICE_X1Y108_AO5),
.I4(CLBLL_L_X2Y108_SLICE_X1Y108_AO6),
.I5(CLBLL_L_X2Y110_SLICE_X0Y110_BQ),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_BO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfff8ff88f8f88888)
  ) CLBLL_L_X2Y110_SLICE_X0Y110_ALUT (
.I0(CLBLL_L_X2Y110_SLICE_X1Y110_AQ),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLL_L_X2Y110_SLICE_X0Y110_AQ),
.I3(LIOB33_X0Y113_IOB_X0Y114_I),
.I4(CLBLL_L_X2Y108_SLICE_X1Y108_AO6),
.I5(CLBLL_L_X2Y108_SLICE_X1Y108_AO5),
.O5(CLBLL_L_X2Y110_SLICE_X0Y110_AO5),
.O6(CLBLL_L_X2Y110_SLICE_X0Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X2Y110_SLICE_X1Y110_AO6),
.Q(CLBLL_L_X2Y110_SLICE_X1Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffff00ff00)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X2Y110_SLICE_X1Y110_CO6),
.I4(1'b1),
.I5(CLBLL_L_X2Y110_SLICE_X1Y110_BO6),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_DO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffe3c3c3c3d)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_CLUT (
.I0(CLBLL_L_X2Y110_SLICE_X0Y110_AQ),
.I1(CLBLL_L_X2Y110_SLICE_X0Y110_BQ),
.I2(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I3(CLBLL_L_X2Y110_SLICE_X0Y110_CQ),
.I4(CLBLL_L_X2Y110_SLICE_X1Y110_AQ),
.I5(CLBLL_L_X2Y109_SLICE_X1Y109_AQ),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_CO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h7bffff7bdeffffde)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_BLUT (
.I0(CLBLM_R_X3Y109_SLICE_X3Y109_CQ),
.I1(CLBLL_L_X2Y109_SLICE_X0Y109_AQ),
.I2(CLBLL_L_X2Y110_SLICE_X1Y110_AQ),
.I3(CLBLL_L_X4Y109_SLICE_X5Y109_BQ),
.I4(CLBLL_L_X2Y110_SLICE_X0Y110_AQ),
.I5(CLBLL_L_X2Y110_SLICE_X0Y110_CQ),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_BO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfefafcf0eeaacc00)
  ) CLBLL_L_X2Y110_SLICE_X1Y110_ALUT (
.I0(CLBLL_L_X2Y110_SLICE_X1Y110_AQ),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y113_IOB_X0Y113_I),
.I3(CLBLL_L_X2Y109_SLICE_X1Y109_AQ),
.I4(CLBLL_L_X2Y108_SLICE_X1Y108_AO6),
.I5(CLBLL_L_X2Y108_SLICE_X1Y108_AO5),
.O5(CLBLL_L_X2Y110_SLICE_X1Y110_AO5),
.O6(CLBLL_L_X2Y110_SLICE_X1Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y104_SLICE_X4Y104_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y104_SLICE_X4Y104_AO6),
.Q(CLBLL_L_X4Y104_SLICE_X4Y104_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y104_SLICE_X4Y104_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y104_SLICE_X4Y104_BO6),
.Q(CLBLL_L_X4Y104_SLICE_X4Y104_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y104_SLICE_X4Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y104_SLICE_X4Y104_DO5),
.O6(CLBLL_L_X4Y104_SLICE_X4Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y104_SLICE_X4Y104_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y104_SLICE_X4Y104_CO5),
.O6(CLBLL_L_X4Y104_SLICE_X4Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaac030c030)
  ) CLBLL_L_X4Y104_SLICE_X4Y104_BLUT (
.I0(CLBLM_R_X5Y105_SLICE_X6Y105_CQ),
.I1(CLBLL_L_X4Y104_SLICE_X4Y104_BQ),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLL_L_X4Y105_SLICE_X5Y105_BO6),
.I4(1'b1),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLL_L_X4Y104_SLICE_X4Y104_BO5),
.O6(CLBLL_L_X4Y104_SLICE_X4Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'habbaabba01100110)
  ) CLBLL_L_X4Y104_SLICE_X4Y104_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(CLBLL_L_X4Y104_SLICE_X4Y104_AQ),
.I3(CLBLL_L_X4Y104_SLICE_X5Y104_CO6),
.I4(1'b1),
.I5(CLBLL_L_X2Y106_SLICE_X1Y106_A5Q),
.O5(CLBLL_L_X4Y104_SLICE_X4Y104_AO5),
.O6(CLBLL_L_X4Y104_SLICE_X4Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y104_SLICE_X5Y104_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y104_SLICE_X5Y104_AO6),
.Q(CLBLL_L_X4Y104_SLICE_X5Y104_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y104_SLICE_X5Y104_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y104_SLICE_X5Y104_BO6),
.Q(CLBLL_L_X4Y104_SLICE_X5Y104_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y104_SLICE_X5Y104_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y104_SLICE_X5Y104_DO5),
.O6(CLBLL_L_X4Y104_SLICE_X5Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333333b333b)
  ) CLBLL_L_X4Y104_SLICE_X5Y104_CLUT (
.I0(CLBLL_L_X4Y104_SLICE_X5Y104_BQ),
.I1(CLBLL_L_X2Y106_SLICE_X0Y106_DQ),
.I2(CLBLM_R_X3Y105_SLICE_X3Y105_AQ),
.I3(CLBLL_L_X4Y104_SLICE_X5Y104_AQ),
.I4(1'b1),
.I5(CLBLL_L_X4Y105_SLICE_X5Y105_BO6),
.O5(CLBLL_L_X4Y104_SLICE_X5Y104_CO5),
.O6(CLBLL_L_X4Y104_SLICE_X5Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000fe0001)
  ) CLBLL_L_X4Y104_SLICE_X5Y104_BLUT (
.I0(CLBLM_R_X3Y105_SLICE_X3Y105_AQ),
.I1(CLBLL_L_X4Y105_SLICE_X5Y105_BO6),
.I2(CLBLL_L_X4Y104_SLICE_X5Y104_AQ),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(CLBLL_L_X4Y104_SLICE_X5Y104_BQ),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLL_L_X4Y104_SLICE_X5Y104_BO5),
.O6(CLBLL_L_X4Y104_SLICE_X5Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa30213021)
  ) CLBLL_L_X4Y104_SLICE_X5Y104_ALUT (
.I0(CLBLM_R_X3Y105_SLICE_X3Y105_AQ),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(CLBLL_L_X4Y104_SLICE_X5Y104_AQ),
.I3(CLBLL_L_X4Y105_SLICE_X5Y105_BO6),
.I4(1'b1),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLL_L_X4Y104_SLICE_X5Y104_AO5),
.O6(CLBLL_L_X4Y104_SLICE_X5Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y105_SLICE_X4Y105_AO6),
.Q(CLBLL_L_X4Y105_SLICE_X4Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y105_SLICE_X4Y105_BO6),
.Q(CLBLL_L_X4Y105_SLICE_X4Y105_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y105_SLICE_X4Y105_CO6),
.Q(CLBLL_L_X4Y105_SLICE_X4Y105_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y105_SLICE_X4Y105_DO6),
.Q(CLBLL_L_X4Y105_SLICE_X4Y105_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc88508850)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_DLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLL_L_X4Y105_SLICE_X4Y105_CQ),
.I2(CLBLL_L_X4Y105_SLICE_X4Y105_DQ),
.I3(CLBLM_R_X3Y104_SLICE_X3Y104_DO6),
.I4(1'b1),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLL_L_X4Y105_SLICE_X4Y105_DO5),
.O6(CLBLL_L_X4Y105_SLICE_X4Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00a404a404)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLL_L_X4Y105_SLICE_X4Y105_CQ),
.I2(CLBLM_R_X3Y104_SLICE_X3Y104_DO6),
.I3(CLBLL_L_X4Y105_SLICE_X4Y105_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLL_L_X4Y105_SLICE_X4Y105_CO5),
.O6(CLBLL_L_X4Y105_SLICE_X4Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0a0a04444)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_BLUT (
.I0(CLBLM_R_X3Y104_SLICE_X3Y104_DO6),
.I1(CLBLL_L_X4Y105_SLICE_X4Y105_BQ),
.I2(CLBLM_R_X3Y104_SLICE_X3Y104_AQ),
.I3(1'b1),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLL_L_X4Y105_SLICE_X4Y105_BO5),
.O6(CLBLL_L_X4Y105_SLICE_X4Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000003c003c)
  ) CLBLL_L_X4Y105_SLICE_X4Y105_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y105_SLICE_X5Y105_DO6),
.I2(CLBLL_L_X4Y105_SLICE_X4Y105_AQ),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(CLBLL_L_X4Y105_SLICE_X5Y105_AQ),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLL_L_X4Y105_SLICE_X4Y105_AO5),
.O6(CLBLL_L_X4Y105_SLICE_X4Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y105_SLICE_X5Y105_AO6),
.Q(CLBLL_L_X4Y105_SLICE_X5Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a000000000000)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_DLUT (
.I0(CLBLM_R_X5Y105_SLICE_X7Y105_AQ),
.I1(1'b1),
.I2(CLBLL_L_X4Y106_SLICE_X5Y106_DO6),
.I3(1'b1),
.I4(CLBLL_L_X4Y105_SLICE_X5Y105_AQ),
.I5(CLBLM_R_X5Y105_SLICE_X7Y105_A5Q),
.O5(CLBLL_L_X4Y105_SLICE_X5Y105_DO5),
.O6(CLBLL_L_X4Y105_SLICE_X5Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010000003333)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_CLUT (
.I0(CLBLL_L_X4Y105_SLICE_X4Y105_AQ),
.I1(CLBLM_R_X3Y105_SLICE_X3Y105_AQ),
.I2(CLBLL_L_X4Y106_SLICE_X5Y106_CO6),
.I3(CLBLL_L_X4Y105_SLICE_X5Y105_AQ),
.I4(CLBLL_L_X4Y104_SLICE_X5Y104_AQ),
.I5(CLBLL_L_X2Y106_SLICE_X0Y106_BQ),
.O5(CLBLL_L_X4Y105_SLICE_X5Y105_CO5),
.O6(CLBLL_L_X4Y105_SLICE_X5Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffbfff00000000)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_BLUT (
.I0(CLBLL_L_X4Y106_SLICE_X5Y106_DO6),
.I1(CLBLM_R_X5Y105_SLICE_X7Y105_A5Q),
.I2(CLBLL_L_X4Y105_SLICE_X5Y105_AQ),
.I3(CLBLM_R_X5Y105_SLICE_X7Y105_AQ),
.I4(CLBLL_L_X4Y105_SLICE_X4Y105_AQ),
.I5(CLBLL_L_X2Y106_SLICE_X0Y106_BQ),
.O5(CLBLL_L_X4Y105_SLICE_X5Y105_BO5),
.O6(CLBLL_L_X4Y105_SLICE_X5Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccb4f00000)
  ) CLBLL_L_X4Y105_SLICE_X5Y105_ALUT (
.I0(CLBLL_L_X4Y106_SLICE_X5Y106_DO6),
.I1(CLBLM_R_X5Y105_SLICE_X7Y105_A5Q),
.I2(CLBLL_L_X4Y105_SLICE_X5Y105_AQ),
.I3(CLBLM_R_X5Y105_SLICE_X7Y105_AQ),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLL_L_X4Y105_SLICE_X5Y105_AO5),
.O6(CLBLL_L_X4Y105_SLICE_X5Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y106_SLICE_X4Y106_AO6),
.Q(CLBLL_L_X4Y106_SLICE_X4Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y106_SLICE_X4Y106_BO6),
.Q(CLBLL_L_X4Y106_SLICE_X4Y106_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y106_SLICE_X4Y106_CO6),
.Q(CLBLL_L_X4Y106_SLICE_X4Y106_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hfbffffffffffffff)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_DLUT (
.I0(CLBLL_L_X4Y107_SLICE_X5Y107_AQ),
.I1(CLBLL_L_X4Y106_SLICE_X4Y106_CQ),
.I2(CLBLL_L_X4Y107_SLICE_X4Y107_B5Q),
.I3(CLBLL_L_X4Y107_SLICE_X4Y107_AQ),
.I4(CLBLL_L_X4Y106_SLICE_X4Y106_BQ),
.I5(CLBLM_R_X3Y109_SLICE_X3Y109_DO6),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_DO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f01144f0f01144)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_CLUT (
.I0(LIOB33_X0Y105_IOB_X0Y106_I),
.I1(CLBLL_L_X4Y106_SLICE_X4Y106_CQ),
.I2(CLBLL_L_X4Y107_SLICE_X4Y107_B5Q),
.I3(CLBLL_L_X4Y107_SLICE_X4Y107_DO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_CO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hedeecccc22220000)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_BLUT (
.I0(CLBLL_L_X4Y106_SLICE_X4Y106_BQ),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLL_L_X4Y107_SLICE_X5Y107_AQ),
.I3(CLBLM_R_X3Y109_SLICE_X3Y109_DO6),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLL_L_X4Y107_SLICE_X4Y107_AQ),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_BO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00fc30cc00ff33)
  ) CLBLL_L_X4Y106_SLICE_X4Y106_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLL_L_X4Y106_SLICE_X4Y106_AQ),
.I3(CLBLM_R_X3Y106_SLICE_X2Y106_AQ),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLM_R_X3Y106_SLICE_X3Y106_DO6),
.O5(CLBLL_L_X4Y106_SLICE_X4Y106_AO5),
.O6(CLBLL_L_X4Y106_SLICE_X4Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y106_SLICE_X5Y106_AO6),
.Q(CLBLL_L_X4Y106_SLICE_X5Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y106_SLICE_X5Y106_BO6),
.Q(CLBLL_L_X4Y106_SLICE_X5Y106_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff77ffffff5555)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_DLUT (
.I0(CLBLL_L_X4Y106_SLICE_X5Y106_BQ),
.I1(CLBLL_L_X4Y107_SLICE_X4Y107_DO6),
.I2(1'b1),
.I3(CLBLL_L_X4Y106_SLICE_X4Y106_CQ),
.I4(CLBLL_L_X4Y106_SLICE_X5Y106_AQ),
.I5(CLBLL_L_X2Y106_SLICE_X0Y106_BQ),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_DO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff7fffffff5f5)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_CLUT (
.I0(CLBLL_L_X4Y106_SLICE_X5Y106_BQ),
.I1(CLBLL_L_X4Y107_SLICE_X4Y107_DO6),
.I2(CLBLL_L_X4Y106_SLICE_X5Y106_AQ),
.I3(CLBLL_L_X4Y106_SLICE_X4Y106_CQ),
.I4(CLBLM_R_X5Y105_SLICE_X7Y105_BO5),
.I5(CLBLL_L_X2Y106_SLICE_X0Y106_BQ),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_CO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaac0909090)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_BLUT (
.I0(CLBLL_L_X4Y106_SLICE_X5Y106_AQ),
.I1(CLBLL_L_X4Y106_SLICE_X5Y106_BQ),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLL_L_X4Y106_SLICE_X4Y106_DO6),
.I4(CLBLL_L_X2Y106_SLICE_X0Y106_BQ),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_BO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff090500000905)
  ) CLBLL_L_X4Y106_SLICE_X5Y106_ALUT (
.I0(CLBLL_L_X4Y106_SLICE_X5Y106_AQ),
.I1(CLBLL_L_X2Y106_SLICE_X0Y106_BQ),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLL_L_X4Y106_SLICE_X4Y106_DO6),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLL_L_X4Y106_SLICE_X4Y106_CQ),
.O5(CLBLL_L_X4Y106_SLICE_X5Y106_AO5),
.O6(CLBLL_L_X4Y106_SLICE_X5Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y107_SLICE_X4Y107_BO5),
.Q(CLBLL_L_X4Y107_SLICE_X4Y107_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y107_SLICE_X4Y107_AO6),
.Q(CLBLL_L_X4Y107_SLICE_X4Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y107_SLICE_X4Y107_BO6),
.Q(CLBLL_L_X4Y107_SLICE_X4Y107_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000404400000000)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_DLUT (
.I0(CLBLL_L_X4Y107_SLICE_X5Y107_AQ),
.I1(CLBLL_L_X4Y107_SLICE_X4Y107_AQ),
.I2(CLBLL_L_X2Y109_SLICE_X1Y109_CO5),
.I3(CLBLL_L_X4Y108_SLICE_X4Y108_CO6),
.I4(CLBLL_L_X4Y107_SLICE_X4Y107_B5Q),
.I5(CLBLL_L_X4Y106_SLICE_X4Y106_BQ),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_DO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb0f04000f0f00000)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_CLUT (
.I0(CLBLL_L_X4Y107_SLICE_X5Y107_AQ),
.I1(CLBLL_L_X4Y107_SLICE_X4Y107_AQ),
.I2(CLBLM_R_X3Y107_SLICE_X2Y107_AO6),
.I3(CLBLL_L_X4Y106_SLICE_X4Y106_BQ),
.I4(CLBLL_L_X4Y107_SLICE_X4Y107_B5Q),
.I5(CLBLM_R_X3Y109_SLICE_X3Y109_DO6),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_CO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfa50fa50eeeecccc)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_BLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLL_L_X4Y107_SLICE_X4Y107_CO6),
.I2(CLBLL_L_X4Y107_SLICE_X5Y107_CO6),
.I3(LIOB33_X0Y117_IOB_X0Y118_I),
.I4(CLBLL_L_X4Y106_SLICE_X4Y106_BQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_BO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heaea1040eaea1040)
  ) CLBLL_L_X4Y107_SLICE_X4Y107_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLL_L_X4Y107_SLICE_X4Y107_AQ),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_R_X3Y109_SLICE_X3Y109_DO6),
.I4(CLBLL_L_X4Y107_SLICE_X5Y107_AQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X4Y107_AO5),
.O6(CLBLL_L_X4Y107_SLICE_X4Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y107_SLICE_X5Y107_BO5),
.Q(CLBLL_L_X4Y107_SLICE_X5Y107_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y107_SLICE_X5Y107_AO6),
.Q(CLBLL_L_X4Y107_SLICE_X5Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000088000000)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_DLUT (
.I0(CLBLL_L_X4Y105_SLICE_X4Y105_BQ),
.I1(CLBLL_L_X4Y105_SLICE_X4Y105_CQ),
.I2(1'b1),
.I3(CLBLL_L_X4Y105_SLICE_X4Y105_DQ),
.I4(CLBLM_R_X3Y104_SLICE_X3Y104_AQ),
.I5(CLBLL_L_X4Y107_SLICE_X5Y107_BO6),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_DO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffe08000000)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_CLUT (
.I0(CLBLL_L_X4Y105_SLICE_X4Y105_BQ),
.I1(CLBLL_L_X4Y105_SLICE_X4Y105_CQ),
.I2(LIOB33_X0Y107_IOB_X0Y107_I),
.I3(CLBLM_R_X3Y104_SLICE_X3Y104_AQ),
.I4(CLBLL_L_X4Y105_SLICE_X4Y105_DQ),
.I5(CLBLL_L_X4Y107_SLICE_X4Y107_BQ),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_CO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'heeee4444fe0ef404)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_BLUT (
.I0(LIOB33_X0Y107_IOB_X0Y107_I),
.I1(CLBLL_L_X4Y107_SLICE_X5Y107_A5Q),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLL_L_X4Y107_SLICE_X4Y107_BQ),
.I4(CLBLL_L_X4Y107_SLICE_X5Y107_CO6),
.I5(1'b1),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_BO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff3c0000003c)
  ) CLBLL_L_X4Y107_SLICE_X5Y107_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y109_SLICE_X3Y109_DO6),
.I2(CLBLL_L_X4Y107_SLICE_X5Y107_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLL_L_X4Y107_SLICE_X5Y107_A5Q),
.O5(CLBLL_L_X4Y107_SLICE_X5Y107_AO5),
.O6(CLBLL_L_X4Y107_SLICE_X5Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffffffffdcff)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_DLUT (
.I0(CLBLM_R_X3Y110_SLICE_X2Y110_BQ),
.I1(CLBLM_R_X3Y108_SLICE_X3Y108_BO6),
.I2(CLBLL_L_X4Y109_SLICE_X4Y109_DO6),
.I3(CLBLM_R_X3Y109_SLICE_X2Y109_CO6),
.I4(CLBLL_L_X2Y109_SLICE_X1Y109_CO6),
.I5(CLBLM_R_X3Y108_SLICE_X2Y108_CO6),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_DO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff8e0affffaf0a)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_CLUT (
.I0(CLBLM_R_X3Y110_SLICE_X2Y110_BQ),
.I1(CLBLL_L_X4Y109_SLICE_X5Y109_CO6),
.I2(CLBLL_L_X4Y109_SLICE_X4Y109_DO6),
.I3(CLBLM_R_X3Y109_SLICE_X2Y109_CO6),
.I4(CLBLL_L_X2Y109_SLICE_X1Y109_CO6),
.I5(CLBLM_R_X3Y108_SLICE_X3Y108_CO6),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_CO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000009000009)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_BLUT (
.I0(CLBLM_R_X3Y110_SLICE_X3Y110_A5Q),
.I1(CLBLL_L_X4Y109_SLICE_X4Y109_A5Q),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_R_X3Y109_SLICE_X2Y109_BQ),
.I4(CLBLL_L_X4Y109_SLICE_X4Y109_BQ),
.I5(CLBLM_R_X3Y110_SLICE_X3Y110_BO6),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_BO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ffff9009ffff)
  ) CLBLL_L_X4Y108_SLICE_X4Y108_ALUT (
.I0(CLBLM_R_X3Y110_SLICE_X3Y110_A5Q),
.I1(CLBLL_L_X4Y109_SLICE_X4Y109_A5Q),
.I2(CLBLL_L_X4Y109_SLICE_X4Y109_BQ),
.I3(CLBLM_R_X3Y109_SLICE_X2Y109_BQ),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLM_R_X3Y110_SLICE_X3Y110_BO6),
.O5(CLBLL_L_X4Y108_SLICE_X4Y108_AO5),
.O6(CLBLL_L_X4Y108_SLICE_X4Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_DO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_CO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_BO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y108_SLICE_X5Y108_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y108_SLICE_X5Y108_AO5),
.O6(CLBLL_L_X4Y108_SLICE_X5Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y109_SLICE_X4Y109_CO6),
.Q(CLBLL_L_X4Y109_SLICE_X4Y109_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y109_SLICE_X4Y109_AO6),
.Q(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y109_SLICE_X4Y109_BO6),
.Q(CLBLL_L_X4Y109_SLICE_X4Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hb3b3a0a0ff00ffff)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_DLUT (
.I0(CLBLL_L_X2Y108_SLICE_X1Y108_BO6),
.I1(LIOB33_X0Y109_IOB_X0Y110_I),
.I2(CLBLL_L_X2Y109_SLICE_X0Y109_AQ),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(CLBLL_L_X2Y106_SLICE_X0Y106_CQ),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_DO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f015400fff0fff)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_CLUT (
.I0(CLBLL_L_X4Y108_SLICE_X4Y108_AO6),
.I1(CLBLM_R_X3Y106_SLICE_X3Y106_CO6),
.I2(CLBLM_R_X3Y109_SLICE_X3Y109_BQ),
.I3(CLBLL_L_X4Y109_SLICE_X4Y109_A5Q),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_CO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'habae0404aeae0404)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_BLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLL_L_X4Y109_SLICE_X4Y109_BQ),
.I2(CLBLL_L_X4Y108_SLICE_X4Y108_AO6),
.I3(CLBLM_R_X3Y109_SLICE_X3Y109_BQ),
.I4(CLBLL_L_X4Y109_SLICE_X4Y109_A5Q),
.I5(CLBLM_R_X3Y106_SLICE_X3Y106_CO6),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_BO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h88d8889c88d888d8)
  ) CLBLL_L_X4Y109_SLICE_X4Y109_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLL_L_X4Y109_SLICE_X4Y109_BQ),
.I2(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.I3(CLBLL_L_X4Y108_SLICE_X4Y108_AO6),
.I4(CLBLL_L_X4Y109_SLICE_X4Y109_CO5),
.I5(CLBLM_R_X3Y106_SLICE_X3Y106_CO6),
.O5(CLBLL_L_X4Y109_SLICE_X4Y109_AO5),
.O6(CLBLL_L_X4Y109_SLICE_X4Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y109_SLICE_X5Y109_AO6),
.Q(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLL_L_X4Y109_SLICE_X5Y109_BO6),
.Q(CLBLL_L_X4Y109_SLICE_X5Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_DO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c005d55dd55dd55)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_CLUT (
.I0(CLBLM_R_X3Y109_SLICE_X3Y109_AO5),
.I1(CLBLM_R_X3Y110_SLICE_X2Y110_A5Q),
.I2(CLBLL_L_X4Y109_SLICE_X5Y109_BQ),
.I3(CLBLL_L_X4Y109_SLICE_X4Y109_DO5),
.I4(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I5(CLBLL_L_X2Y108_SLICE_X1Y108_BO6),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_CO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffc0c0c030c0c0)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y109_SLICE_X5Y109_BQ),
.I2(CLBLL_L_X2Y109_SLICE_X0Y109_BO5),
.I3(CLBLM_R_X3Y106_SLICE_X3Y106_BO6),
.I4(CLBLM_R_X3Y109_SLICE_X3Y109_CQ),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_BO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hececececa060a0a0)
  ) CLBLL_L_X4Y109_SLICE_X5Y109_ALUT (
.I0(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I1(CLBLL_L_X4Y109_SLICE_X5Y109_BQ),
.I2(CLBLL_L_X2Y109_SLICE_X0Y109_BO5),
.I3(CLBLM_R_X3Y106_SLICE_X3Y106_BO6),
.I4(CLBLM_R_X3Y109_SLICE_X3Y109_CQ),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLL_L_X4Y109_SLICE_X5Y109_AO5),
.O6(CLBLL_L_X4Y109_SLICE_X5Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y104_SLICE_X2Y104_AO6),
.Q(CLBLM_R_X3Y104_SLICE_X2Y104_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y104_SLICE_X2Y104_BO6),
.Q(CLBLM_R_X3Y104_SLICE_X2Y104_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y104_SLICE_X2Y104_CO6),
.Q(CLBLM_R_X3Y104_SLICE_X2Y104_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_D_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y104_SLICE_X2Y104_DO6),
.Q(CLBLM_R_X3Y104_SLICE_X2Y104_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00a1f0ff000000)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_DLUT (
.I0(CLBLL_L_X4Y105_SLICE_X5Y105_BO6),
.I1(CLBLM_R_X3Y104_SLICE_X2Y104_CQ),
.I2(CLBLM_R_X3Y104_SLICE_X2Y104_DQ),
.I3(CLBLL_L_X4Y104_SLICE_X4Y104_BQ),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_R_X3Y104_SLICE_X2Y104_DO5),
.O6(CLBLM_R_X3Y104_SLICE_X2Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f098ccf0f00000)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_CLUT (
.I0(CLBLL_L_X4Y105_SLICE_X5Y105_BO6),
.I1(CLBLM_R_X3Y104_SLICE_X2Y104_CQ),
.I2(CLBLM_R_X3Y104_SLICE_X2Y104_DQ),
.I3(CLBLL_L_X4Y104_SLICE_X4Y104_BQ),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_R_X3Y104_SLICE_X2Y104_CO5),
.O6(CLBLM_R_X3Y104_SLICE_X2Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f098009800)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_BLUT (
.I0(CLBLM_R_X3Y105_SLICE_X2Y105_CO6),
.I1(CLBLM_R_X3Y104_SLICE_X2Y104_BQ),
.I2(CLBLM_R_X3Y104_SLICE_X2Y104_AQ),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(1'b1),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X3Y104_SLICE_X2Y104_BO5),
.O6(CLBLM_R_X3Y104_SLICE_X2Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000a100a100)
  ) CLBLM_R_X3Y104_SLICE_X2Y104_ALUT (
.I0(CLBLM_R_X3Y105_SLICE_X2Y105_CO6),
.I1(CLBLM_R_X3Y104_SLICE_X2Y104_BQ),
.I2(CLBLM_R_X3Y104_SLICE_X2Y104_AQ),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(CLBLM_R_X3Y104_SLICE_X2Y104_CQ),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X3Y104_SLICE_X2Y104_AO5),
.O6(CLBLM_R_X3Y104_SLICE_X2Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y104_SLICE_X3Y104_AO6),
.Q(CLBLM_R_X3Y104_SLICE_X3Y104_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y104_SLICE_X3Y104_BO6),
.Q(CLBLM_R_X3Y104_SLICE_X3Y104_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h4f0f4f0f4f0f4f0f)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_DLUT (
.I0(CLBLL_L_X4Y105_SLICE_X5Y105_BO6),
.I1(CLBLL_L_X4Y104_SLICE_X4Y104_BQ),
.I2(CLBLL_L_X2Y106_SLICE_X0Y106_DQ),
.I3(CLBLM_R_X3Y104_SLICE_X2Y104_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y104_SLICE_X3Y104_DO5),
.O6(CLBLM_R_X3Y104_SLICE_X3Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff0f0ffffe0f0)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_CLUT (
.I0(CLBLL_L_X4Y105_SLICE_X5Y105_BO6),
.I1(CLBLM_R_X3Y105_SLICE_X3Y105_AQ),
.I2(CLBLL_L_X2Y106_SLICE_X0Y106_DQ),
.I3(CLBLL_L_X4Y104_SLICE_X5Y104_BQ),
.I4(CLBLL_L_X4Y104_SLICE_X4Y104_AQ),
.I5(CLBLL_L_X4Y104_SLICE_X5Y104_AQ),
.O5(CLBLM_R_X3Y104_SLICE_X3Y104_CO5),
.O6(CLBLM_R_X3Y104_SLICE_X3Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'he4a0e4a0b1a0b1a0)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_BLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_R_X3Y104_SLICE_X3Y104_BQ),
.I2(CLBLL_L_X4Y104_SLICE_X4Y104_AQ),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(1'b1),
.I5(CLBLM_R_X3Y104_SLICE_X3Y104_CO6),
.O5(CLBLM_R_X3Y104_SLICE_X3Y104_BO5),
.O6(CLBLM_R_X3Y104_SLICE_X3Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff981000009810)
  ) CLBLM_R_X3Y104_SLICE_X3Y104_ALUT (
.I0(CLBLM_R_X3Y104_SLICE_X3Y104_DO6),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(CLBLM_R_X3Y104_SLICE_X3Y104_AQ),
.I3(LIOB33_X0Y103_IOB_X0Y104_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_R_X3Y110_SLICE_X2Y110_CQ),
.O5(CLBLM_R_X3Y104_SLICE_X3Y104_AO5),
.O6(CLBLM_R_X3Y104_SLICE_X3Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y105_SLICE_X2Y105_AO6),
.Q(CLBLM_R_X3Y105_SLICE_X2Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y105_SLICE_X2Y105_BO6),
.Q(CLBLM_R_X3Y105_SLICE_X2Y105_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0f0f04c4c0c0c)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_DLUT (
.I0(CLBLM_R_X3Y105_SLICE_X2Y105_CO5),
.I1(CLBLM_R_X5Y105_SLICE_X6Y105_CQ),
.I2(CLBLL_L_X2Y106_SLICE_X0Y106_DQ),
.I3(1'b1),
.I4(CLBLL_L_X2Y105_SLICE_X1Y105_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y105_SLICE_X2Y105_DO5),
.O6(CLBLM_R_X3Y105_SLICE_X2Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00f3f3ff55f7f7)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_CLUT (
.I0(CLBLM_R_X3Y104_SLICE_X2Y104_BQ),
.I1(CLBLM_R_X3Y105_SLICE_X3Y105_A5Q),
.I2(CLBLM_R_X3Y105_SLICE_X3Y105_DO6),
.I3(CLBLL_L_X4Y105_SLICE_X5Y105_BO6),
.I4(CLBLM_R_X3Y108_SLICE_X3Y108_DO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y105_SLICE_X2Y105_CO5),
.O6(CLBLM_R_X3Y105_SLICE_X2Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hb0e4b0e4a0a0a0a0)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_BLUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_R_X3Y105_SLICE_X2Y105_BQ),
.I2(CLBLM_R_X3Y105_SLICE_X2Y105_AQ),
.I3(CLBLM_R_X3Y105_SLICE_X2Y105_DO5),
.I4(1'b1),
.I5(LIOB33_X0Y105_IOB_X0Y106_I),
.O5(CLBLM_R_X3Y105_SLICE_X2Y105_BO5),
.O6(CLBLM_R_X3Y105_SLICE_X2Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'habfaaaaa01500000)
  ) CLBLM_R_X3Y105_SLICE_X2Y105_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLM_R_X3Y105_SLICE_X2Y105_BQ),
.I2(CLBLM_R_X3Y105_SLICE_X2Y105_AQ),
.I3(CLBLM_R_X3Y105_SLICE_X2Y105_DO5),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLL_L_X2Y105_SLICE_X1Y105_AQ),
.O5(CLBLM_R_X3Y105_SLICE_X2Y105_AO5),
.O6(CLBLM_R_X3Y105_SLICE_X2Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y105_SLICE_X3Y105_BO6),
.Q(CLBLM_R_X3Y105_SLICE_X3Y105_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y105_SLICE_X3Y105_AO6),
.Q(CLBLM_R_X3Y105_SLICE_X3Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3fff0f0ffffffff)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y104_SLICE_X5Y104_BQ),
.I2(CLBLL_L_X4Y104_SLICE_X4Y104_AQ),
.I3(CLBLL_L_X4Y105_SLICE_X5Y105_CO6),
.I4(CLBLL_L_X2Y106_SLICE_X0Y106_DQ),
.I5(CLBLM_R_X3Y104_SLICE_X3Y104_BQ),
.O5(CLBLM_R_X3Y105_SLICE_X3Y105_DO5),
.O6(CLBLM_R_X3Y105_SLICE_X3Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h440044000000c000)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_CLUT (
.I0(CLBLL_L_X4Y105_SLICE_X5Y105_BO6),
.I1(CLBLL_L_X2Y105_SLICE_X1Y105_AQ),
.I2(CLBLM_R_X3Y105_SLICE_X3Y105_A5Q),
.I3(CLBLM_R_X3Y104_SLICE_X2Y104_BQ),
.I4(CLBLM_R_X3Y105_SLICE_X3Y105_DO6),
.I5(CLBLM_R_X3Y108_SLICE_X3Y108_DO6),
.O5(CLBLM_R_X3Y105_SLICE_X3Y105_CO5),
.O6(CLBLM_R_X3Y105_SLICE_X3Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hce02cd01ffffaaaa)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_BLUT (
.I0(CLBLM_R_X3Y105_SLICE_X3Y105_DO6),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_R_X3Y104_SLICE_X3Y104_BQ),
.I4(CLBLM_R_X3Y105_SLICE_X3Y105_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y105_SLICE_X3Y105_BO5),
.O6(CLBLM_R_X3Y105_SLICE_X3Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff30ff0300300003)
  ) CLBLM_R_X3Y105_SLICE_X3Y105_ALUT (
.I0(1'b1),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(CLBLM_R_X3Y105_SLICE_X3Y105_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLL_L_X4Y105_SLICE_X5Y105_BO6),
.I5(CLBLM_R_X3Y105_SLICE_X3Y105_A5Q),
.O5(CLBLM_R_X3Y105_SLICE_X3Y105_AO5),
.O6(CLBLM_R_X3Y105_SLICE_X3Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y106_SLICE_X2Y106_AO6),
.Q(CLBLM_R_X3Y106_SLICE_X2Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7000ffff7000ffff)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_DLUT (
.I0(CLBLL_L_X4Y105_SLICE_X5Y105_DO6),
.I1(CLBLL_L_X4Y105_SLICE_X4Y105_AQ),
.I2(CLBLM_R_X3Y108_SLICE_X3Y108_DO6),
.I3(CLBLL_L_X2Y106_SLICE_X0Y106_BQ),
.I4(CLBLL_L_X2Y110_SLICE_X1Y110_DO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_DO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000808f0000b0bf)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_CLUT (
.I0(CLBLL_L_X4Y105_SLICE_X4Y105_AQ),
.I1(CLBLL_L_X2Y106_SLICE_X0Y106_BQ),
.I2(CLBLM_R_X3Y108_SLICE_X3Y108_DO6),
.I3(CLBLM_R_X3Y105_SLICE_X3Y105_A5Q),
.I4(CLBLL_L_X2Y110_SLICE_X1Y110_DO6),
.I5(CLBLL_L_X2Y106_SLICE_X1Y106_A5Q),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_CO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0007000f000f000f)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_BLUT (
.I0(CLBLM_R_X3Y106_SLICE_X2Y106_AQ),
.I1(CLBLM_R_X3Y105_SLICE_X2Y105_DO5),
.I2(CLBLM_R_X3Y106_SLICE_X3Y106_AO6),
.I3(CLBLL_L_X2Y106_SLICE_X1Y106_DO6),
.I4(CLBLL_L_X2Y106_SLICE_X0Y106_AQ),
.I5(CLBLM_R_X3Y105_SLICE_X2Y105_BQ),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_BO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff3c000000f000)
  ) CLBLM_R_X3Y106_SLICE_X2Y106_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y105_SLICE_X2Y105_DO5),
.I2(CLBLM_R_X3Y106_SLICE_X2Y106_AQ),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_R_X3Y105_SLICE_X2Y105_BQ),
.O5(CLBLM_R_X3Y106_SLICE_X2Y106_AO5),
.O6(CLBLM_R_X3Y106_SLICE_X2Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc505f535c505f535)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_DLUT (
.I0(CLBLM_R_X3Y105_SLICE_X3Y105_A5Q),
.I1(CLBLL_L_X2Y106_SLICE_X0Y106_BQ),
.I2(CLBLM_R_X3Y108_SLICE_X3Y108_DO6),
.I3(CLBLL_L_X4Y105_SLICE_X4Y105_AQ),
.I4(CLBLL_L_X2Y106_SLICE_X1Y106_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_DO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff8f0fffff0000)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_CLUT (
.I0(CLBLM_R_X3Y106_SLICE_X2Y106_AQ),
.I1(CLBLM_R_X5Y105_SLICE_X6Y105_CQ),
.I2(CLBLL_L_X2Y106_SLICE_X0Y106_DQ),
.I3(CLBLM_R_X3Y105_SLICE_X2Y105_BQ),
.I4(CLBLL_L_X2Y106_SLICE_X0Y106_CQ),
.I5(CLBLM_R_X3Y105_SLICE_X3Y105_CO6),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_CO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2eff22ffeeff22ff)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_BLUT (
.I0(CLBLM_R_X3Y105_SLICE_X3Y105_BO5),
.I1(CLBLM_R_X3Y108_SLICE_X3Y108_DO6),
.I2(CLBLL_L_X4Y105_SLICE_X5Y105_DO6),
.I3(CLBLL_L_X2Y110_SLICE_X1Y110_DO6),
.I4(CLBLL_L_X2Y106_SLICE_X0Y106_BQ),
.I5(CLBLL_L_X4Y105_SLICE_X4Y105_AQ),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_BO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333337333333333)
  ) CLBLM_R_X3Y106_SLICE_X3Y106_ALUT (
.I0(CLBLL_L_X4Y104_SLICE_X5Y104_AQ),
.I1(CLBLL_L_X2Y106_SLICE_X0Y106_CQ),
.I2(CLBLL_L_X2Y106_SLICE_X1Y106_BQ),
.I3(CLBLL_L_X4Y105_SLICE_X5Y105_BO6),
.I4(CLBLM_R_X3Y105_SLICE_X3Y105_AQ),
.I5(CLBLL_L_X4Y104_SLICE_X5Y104_BQ),
.O5(CLBLM_R_X3Y106_SLICE_X3Y106_AO5),
.O6(CLBLM_R_X3Y106_SLICE_X3Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y107_SLICE_X2Y107_AO5),
.Q(CLBLM_R_X3Y107_SLICE_X2Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0808000000000000)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_DLUT (
.I0(CLBLL_L_X4Y106_SLICE_X4Y106_AQ),
.I1(CLBLL_L_X4Y107_SLICE_X5Y107_DO6),
.I2(CLBLM_R_X3Y105_SLICE_X3Y105_DO6),
.I3(1'b1),
.I4(CLBLM_R_X3Y109_SLICE_X2Y109_AQ),
.I5(CLBLL_L_X4Y108_SLICE_X4Y108_BO6),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_DO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff5f5dffffffff)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_CLUT (
.I0(CLBLL_L_X4Y109_SLICE_X5Y109_BQ),
.I1(CLBLM_R_X3Y105_SLICE_X3Y105_DO6),
.I2(CLBLM_R_X3Y108_SLICE_X3Y108_DO6),
.I3(CLBLM_R_X3Y105_SLICE_X3Y105_A5Q),
.I4(CLBLM_R_X3Y106_SLICE_X2Y106_DO6),
.I5(CLBLM_R_X3Y109_SLICE_X3Y109_CQ),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_CO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0000020e00000)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_BLUT (
.I0(CLBLM_R_X3Y108_SLICE_X2Y108_BQ),
.I1(CLBLL_L_X2Y106_SLICE_X0Y106_CQ),
.I2(CLBLL_L_X2Y109_SLICE_X1Y109_BQ),
.I3(LIOB33_X0Y115_IOB_X0Y115_I),
.I4(CLBLM_R_X3Y107_SLICE_X2Y107_AO6),
.I5(CLBLL_L_X2Y107_SLICE_X1Y107_AQ),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_BO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00003333bbb8bb88)
  ) CLBLM_R_X3Y107_SLICE_X2Y107_ALUT (
.I0(CLBLM_R_X3Y108_SLICE_X2Y108_BQ),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_R_X3Y107_SLICE_X2Y107_AQ),
.I3(CLBLL_L_X4Y108_SLICE_X4Y108_BO6),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(1'b1),
.O5(CLBLM_R_X3Y107_SLICE_X2Y107_AO5),
.O6(CLBLM_R_X3Y107_SLICE_X2Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000044554444)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_DLUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(CLBLM_R_X3Y106_SLICE_X3Y106_DO6),
.I2(1'b1),
.I3(LIOB33_X0Y111_IOB_X0Y112_I),
.I4(CLBLL_L_X4Y108_SLICE_X4Y108_DO6),
.I5(CLBLL_L_X2Y106_SLICE_X0Y106_CQ),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_DO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c0d0c0c0c0d0c0c)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_CLUT (
.I0(CLBLL_L_X2Y110_SLICE_X1Y110_DO6),
.I1(CLBLM_R_X3Y106_SLICE_X3Y106_DO6),
.I2(CLBLM_R_X3Y108_SLICE_X3Y108_DO6),
.I3(CLBLL_L_X2Y109_SLICE_X1Y109_BQ),
.I4(CLBLL_L_X4Y108_SLICE_X4Y108_DO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_CO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffffff008800a0)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_BLUT (
.I0(CLBLM_R_X3Y108_SLICE_X3Y108_DO6),
.I1(CLBLM_R_X3Y106_SLICE_X2Y106_AQ),
.I2(CLBLL_L_X2Y105_SLICE_X1Y105_AQ),
.I3(CLBLL_L_X2Y106_SLICE_X0Y106_CQ),
.I4(CLBLL_L_X2Y106_SLICE_X0Y106_DQ),
.I5(CLBLM_R_X3Y108_SLICE_X3Y108_AO5),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_BO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3030300030203000)
  ) CLBLM_R_X3Y107_SLICE_X3Y107_ALUT (
.I0(CLBLM_R_X3Y107_SLICE_X3Y107_DO6),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLM_R_X3Y107_SLICE_X3Y107_BO6),
.I4(CLBLM_R_X3Y109_SLICE_X3Y109_DO6),
.I5(CLBLM_R_X3Y107_SLICE_X3Y107_CO6),
.O5(CLBLM_R_X3Y107_SLICE_X3Y107_AO5),
.O6(CLBLM_R_X3Y107_SLICE_X3Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y108_SLICE_X2Y108_AO6),
.Q(CLBLM_R_X3Y108_SLICE_X2Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y108_SLICE_X2Y108_BO6),
.Q(CLBLM_R_X3Y108_SLICE_X2Y108_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hea80ea80ffffffff)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_DLUT (
.I0(CLBLM_R_X3Y108_SLICE_X2Y108_CO5),
.I1(CLBLM_R_X3Y109_SLICE_X2Y109_AQ),
.I2(CLBLM_R_X3Y108_SLICE_X3Y108_BO6),
.I3(CLBLM_R_X3Y110_SLICE_X2Y110_A5Q),
.I4(1'b1),
.I5(CLBLM_R_X3Y109_SLICE_X2Y109_CO5),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_DO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h080f080877007777)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_CLUT (
.I0(CLBLL_L_X2Y108_SLICE_X1Y108_BO6),
.I1(CLBLL_L_X4Y109_SLICE_X5Y109_BQ),
.I2(CLBLM_R_X3Y110_SLICE_X2Y110_A5Q),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(CLBLL_L_X2Y106_SLICE_X0Y106_CQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_CO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ff0c0c0c)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y108_SLICE_X2Y108_BQ),
.I2(CLBLL_L_X4Y108_SLICE_X4Y108_AO6),
.I3(CLBLL_L_X4Y106_SLICE_X4Y106_AQ),
.I4(CLBLL_L_X4Y108_SLICE_X4Y108_BO6),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_BO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ccfc00f0)
  ) CLBLM_R_X3Y108_SLICE_X2Y108_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X4Y108_SLICE_X4Y108_BO6),
.I2(CLBLM_R_X3Y108_SLICE_X2Y108_AQ),
.I3(CLBLL_L_X4Y108_SLICE_X4Y108_AO6),
.I4(CLBLM_R_X3Y107_SLICE_X2Y107_AQ),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X3Y108_SLICE_X2Y108_AO5),
.O6(CLBLM_R_X3Y108_SLICE_X2Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff01ff01ff00ff00)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_DLUT (
.I0(CLBLM_R_X3Y108_SLICE_X2Y108_AQ),
.I1(CLBLL_L_X2Y109_SLICE_X1Y109_BQ),
.I2(CLBLL_L_X2Y110_SLICE_X1Y110_DO6),
.I3(CLBLL_L_X2Y106_SLICE_X0Y106_CQ),
.I4(1'b1),
.I5(LIOB33_X0Y107_IOB_X0Y108_I),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_DO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffff5f5fffff5f7)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_CLUT (
.I0(CLBLM_R_X3Y109_SLICE_X2Y109_AQ),
.I1(CLBLM_R_X3Y109_SLICE_X3Y109_AO6),
.I2(CLBLL_L_X2Y108_SLICE_X1Y108_CO6),
.I3(CLBLM_R_X3Y110_SLICE_X2Y110_A5Q),
.I4(CLBLM_R_X3Y108_SLICE_X3Y108_BO5),
.I5(CLBLL_L_X2Y108_SLICE_X1Y108_DO6),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_CO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0dddf22222222222)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_BLUT (
.I0(CLBLL_L_X2Y106_SLICE_X0Y106_CQ),
.I1(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.I2(CLBLL_L_X2Y108_SLICE_X1Y108_BO6),
.I3(CLBLM_R_X3Y109_SLICE_X3Y109_CQ),
.I4(CLBLM_R_X3Y109_SLICE_X2Y109_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_BO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0fcfcf0000aa00)
  ) CLBLM_R_X3Y108_SLICE_X3Y108_ALUT (
.I0(LIOB33_X0Y113_IOB_X0Y113_I),
.I1(CLBLL_L_X4Y108_SLICE_X4Y108_AO6),
.I2(LIOB33_X0Y105_IOB_X0Y106_I),
.I3(CLBLL_L_X2Y106_SLICE_X1Y106_A5Q),
.I4(CLBLL_L_X2Y106_SLICE_X0Y106_CQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y108_SLICE_X3Y108_AO5),
.O6(CLBLM_R_X3Y108_SLICE_X3Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y109_SLICE_X2Y109_BO5),
.Q(CLBLM_R_X3Y109_SLICE_X2Y109_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y109_SLICE_X2Y109_AO6),
.Q(CLBLM_R_X3Y109_SLICE_X2Y109_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y109_SLICE_X2Y109_BO6),
.Q(CLBLM_R_X3Y109_SLICE_X2Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaf0aaf0ffff0000)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_DLUT (
.I0(LIOB33_X0Y111_IOB_X0Y112_I),
.I1(1'b1),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(CLBLL_L_X4Y106_SLICE_X4Y106_AQ),
.I4(CLBLM_R_X3Y109_SLICE_X2Y109_BQ),
.I5(CLBLM_R_X3Y108_SLICE_X3Y108_AO6),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_DO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff70ff778fff88ff)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_CLUT (
.I0(CLBLL_L_X2Y108_SLICE_X1Y108_BO6),
.I1(CLBLL_L_X4Y109_SLICE_X5Y109_AQ),
.I2(LIOB33_X0Y109_IOB_X0Y109_I),
.I3(CLBLM_R_X3Y110_SLICE_X2Y110_AQ),
.I4(CLBLL_L_X2Y106_SLICE_X0Y106_CQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_CO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccaaccaafff0f0f0)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_BLUT (
.I0(CLBLM_R_X3Y109_SLICE_X2Y109_DO6),
.I1(CLBLM_R_X3Y110_SLICE_X3Y110_A5Q),
.I2(CLBLM_R_X3Y107_SLICE_X3Y107_AO6),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(CLBLL_L_X2Y106_SLICE_X0Y106_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_BO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hdeccdecc5a005a00)
  ) CLBLM_R_X3Y109_SLICE_X2Y109_ALUT (
.I0(CLBLL_L_X4Y107_SLICE_X5Y107_DO6),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLM_R_X3Y109_SLICE_X2Y109_AQ),
.I3(CLBLL_L_X2Y109_SLICE_X0Y109_BO6),
.I4(1'b1),
.I5(CLBLL_L_X4Y104_SLICE_X5Y104_BQ),
.O5(CLBLM_R_X3Y109_SLICE_X2Y109_AO5),
.O6(CLBLM_R_X3Y109_SLICE_X2Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y109_SLICE_X3Y109_BO6),
.Q(CLBLM_R_X3Y109_SLICE_X3Y109_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y109_SLICE_X3Y109_CO6),
.Q(CLBLM_R_X3Y109_SLICE_X3Y109_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7f55ff7f15005515)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_DLUT (
.I0(CLBLM_R_X3Y110_SLICE_X2Y110_CQ),
.I1(CLBLM_R_X3Y109_SLICE_X2Y109_CO6),
.I2(CLBLM_R_X3Y108_SLICE_X2Y108_DO6),
.I3(CLBLL_L_X4Y109_SLICE_X4Y109_DO6),
.I4(CLBLM_R_X3Y110_SLICE_X2Y110_BQ),
.I5(CLBLL_L_X2Y109_SLICE_X1Y109_DO6),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_DO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff82ff8282828282)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_CLUT (
.I0(CLBLL_L_X2Y109_SLICE_X0Y109_BO5),
.I1(CLBLM_R_X3Y109_SLICE_X3Y109_CQ),
.I2(CLBLM_R_X3Y106_SLICE_X3Y106_BO6),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(1'b1),
.I5(CLBLM_R_X3Y109_SLICE_X2Y109_BQ),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_CO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0003300cc)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y109_SLICE_X3Y109_BQ),
.I2(CLBLM_R_X3Y108_SLICE_X2Y108_AQ),
.I3(CLBLL_L_X4Y108_SLICE_X4Y108_AO6),
.I4(CLBLM_R_X3Y106_SLICE_X3Y106_CO6),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_BO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000ff0f73737373)
  ) CLBLM_R_X3Y109_SLICE_X3Y109_ALUT (
.I0(LIOB33_X0Y109_IOB_X0Y109_I),
.I1(CLBLM_R_X3Y110_SLICE_X2Y110_AQ),
.I2(CLBLL_L_X2Y106_SLICE_X0Y106_CQ),
.I3(LIOB33_X0Y101_IOB_X0Y101_I),
.I4(CLBLL_L_X4Y109_SLICE_X5Y109_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y109_SLICE_X3Y109_AO5),
.O6(CLBLM_R_X3Y109_SLICE_X3Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y110_SLICE_X2Y110_DO6),
.Q(CLBLM_R_X3Y110_SLICE_X2Y110_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y110_SLICE_X2Y110_AO6),
.Q(CLBLM_R_X3Y110_SLICE_X2Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y110_SLICE_X2Y110_BO6),
.Q(CLBLM_R_X3Y110_SLICE_X2Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y110_SLICE_X2Y110_CO6),
.Q(CLBLM_R_X3Y110_SLICE_X2Y110_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd8a8f88855ffffff)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_DLUT (
.I0(CLBLM_R_X3Y109_SLICE_X2Y109_AQ),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLL_L_X2Y109_SLICE_X0Y109_BO6),
.I3(CLBLM_R_X3Y110_SLICE_X2Y110_A5Q),
.I4(CLBLL_L_X4Y107_SLICE_X5Y107_DO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_DO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffa0a0a0f7a0a8a0)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_CLUT (
.I0(CLBLM_R_X3Y110_SLICE_X2Y110_BQ),
.I1(CLBLM_R_X3Y110_SLICE_X2Y110_AQ),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLL_L_X2Y109_SLICE_X0Y109_BO6),
.I4(CLBLM_R_X3Y110_SLICE_X2Y110_CQ),
.I5(CLBLM_R_X3Y110_SLICE_X2Y110_DO5),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_CO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfcfcf0f0cc0c00c0)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X2Y109_SLICE_X0Y109_BO6),
.I2(CLBLM_R_X3Y110_SLICE_X2Y110_AQ),
.I3(CLBLM_R_X3Y110_SLICE_X2Y110_DO5),
.I4(CLBLM_R_X3Y110_SLICE_X2Y110_BQ),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_BO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'heaaeeaaec00cc00c)
  ) CLBLM_R_X3Y110_SLICE_X2Y110_ALUT (
.I0(LIOB33_X0Y117_IOB_X0Y117_I),
.I1(CLBLL_L_X2Y109_SLICE_X0Y109_BO6),
.I2(CLBLM_R_X3Y110_SLICE_X2Y110_AQ),
.I3(CLBLM_R_X3Y110_SLICE_X2Y110_DO5),
.I4(1'b1),
.I5(CLBLM_R_X3Y110_SLICE_X2Y110_A5Q),
.O5(CLBLM_R_X3Y110_SLICE_X2Y110_AO5),
.O6(CLBLM_R_X3Y110_SLICE_X2Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y110_SLICE_X3Y110_AO5),
.Q(CLBLM_R_X3Y110_SLICE_X3Y110_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X3Y110_SLICE_X3Y110_AO6),
.Q(CLBLM_R_X3Y110_SLICE_X3Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he4e4ff00e4e4ff00)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_DLUT (
.I0(CLBLL_L_X4Y106_SLICE_X4Y106_AQ),
.I1(LIOB33_X0Y101_IOB_X0Y101_I),
.I2(LIOB33_X0Y111_IOB_X0Y111_I),
.I3(CLBLM_R_X3Y110_SLICE_X3Y110_A5Q),
.I4(CLBLM_R_X3Y108_SLICE_X3Y108_AO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_DO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hfc5cfc5cac0cac0c)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_CLUT (
.I0(CLBLL_L_X4Y106_SLICE_X4Y106_AQ),
.I1(CLBLM_R_X3Y110_SLICE_X3Y110_AQ),
.I2(CLBLM_R_X3Y108_SLICE_X3Y108_AO6),
.I3(LIOB33_X0Y109_IOB_X0Y110_I),
.I4(1'b1),
.I5(LIOB33_SING_X0Y100_IOB_X0Y100_I),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_CO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5faf5faf5ebf5eb)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_BLUT (
.I0(CLBLM_R_X3Y109_SLICE_X3Y109_BQ),
.I1(CLBLM_R_X3Y109_SLICE_X2Y109_BQ),
.I2(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.I3(CLBLM_R_X3Y110_SLICE_X3Y110_AQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y110_SLICE_X3Y110_A5Q),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_BO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0c0ee22ee22)
  ) CLBLM_R_X3Y110_SLICE_X3Y110_ALUT (
.I0(CLBLM_R_X3Y110_SLICE_X3Y110_DO6),
.I1(LIOB33_X0Y117_IOB_X0Y117_I),
.I2(CLBLL_L_X4Y109_SLICE_X4Y109_AQ),
.I3(CLBLM_R_X3Y110_SLICE_X3Y110_AQ),
.I4(CLBLM_R_X3Y110_SLICE_X3Y110_CO6),
.I5(1'b1),
.O5(CLBLM_R_X3Y110_SLICE_X3Y110_AO5),
.O6(CLBLM_R_X3Y110_SLICE_X3Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y105_SLICE_X6Y105_AO6),
.Q(CLBLM_R_X5Y105_SLICE_X6Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y105_SLICE_X6Y105_BO6),
.Q(CLBLM_R_X5Y105_SLICE_X6Y105_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y105_SLICE_X6Y105_CO6),
.Q(CLBLM_R_X5Y105_SLICE_X6Y105_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f000c030f00040b)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_DLUT (
.I0(CLBLL_L_X2Y106_SLICE_X0Y106_DQ),
.I1(CLBLM_R_X5Y105_SLICE_X6Y105_CQ),
.I2(LIOB33_X0Y117_IOB_X0Y117_I),
.I3(CLBLM_R_X5Y106_SLICE_X6Y106_AQ),
.I4(LIOB33_X0Y105_IOB_X0Y106_I),
.I5(CLBLM_R_X3Y105_SLICE_X3Y105_CO6),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_DO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffaaaaaaff080000)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_CLUT (
.I0(CLBLM_R_X5Y105_SLICE_X6Y105_BQ),
.I1(CLBLM_R_X5Y105_SLICE_X6Y105_AQ),
.I2(CLBLM_R_X3Y105_SLICE_X2Y105_DO6),
.I3(CLBLM_R_X5Y105_SLICE_X6Y105_CQ),
.I4(CLBLM_R_X5Y105_SLICE_X6Y105_DO6),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_CO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00088f0f0009c)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_BLUT (
.I0(CLBLM_R_X3Y105_SLICE_X2Y105_DO6),
.I1(CLBLM_R_X5Y105_SLICE_X6Y105_BQ),
.I2(CLBLM_R_X5Y105_SLICE_X6Y105_AQ),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(CLBLM_R_X5Y105_SLICE_X6Y105_CQ),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_BO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff84ff8484848484)
  ) CLBLM_R_X5Y105_SLICE_X6Y105_ALUT (
.I0(CLBLM_R_X3Y105_SLICE_X2Y105_DO6),
.I1(CLBLM_R_X5Y105_SLICE_X6Y105_DO6),
.I2(CLBLM_R_X5Y105_SLICE_X6Y105_AQ),
.I3(LIOB33_X0Y117_IOB_X0Y117_I),
.I4(1'b1),
.I5(CLBLL_L_X4Y105_SLICE_X4Y105_DQ),
.O5(CLBLM_R_X5Y105_SLICE_X6Y105_AO5),
.O6(CLBLM_R_X5Y105_SLICE_X6Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y105_SLICE_X7Y105_BO6),
.Q(CLBLM_R_X5Y105_SLICE_X7Y105_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y105_SLICE_X7Y105_AO6),
.Q(CLBLM_R_X5Y105_SLICE_X7Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_DO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_CO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f09c003f3f3f3f)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_BLUT (
.I0(CLBLL_L_X4Y106_SLICE_X5Y106_DO6),
.I1(CLBLM_R_X5Y105_SLICE_X7Y105_A5Q),
.I2(CLBLM_R_X5Y105_SLICE_X7Y105_AQ),
.I3(LIOB33_X0Y105_IOB_X0Y106_I),
.I4(LIOB33_X0Y117_IOB_X0Y117_I),
.I5(1'b1),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_BO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0021212121)
  ) CLBLM_R_X5Y105_SLICE_X7Y105_ALUT (
.I0(CLBLL_L_X4Y106_SLICE_X5Y106_DO6),
.I1(LIOB33_X0Y105_IOB_X0Y106_I),
.I2(CLBLM_R_X5Y105_SLICE_X7Y105_AQ),
.I3(CLBLL_L_X4Y106_SLICE_X5Y106_BQ),
.I4(1'b1),
.I5(LIOB33_X0Y117_IOB_X0Y117_I),
.O5(CLBLM_R_X5Y105_SLICE_X7Y105_AO5),
.O6(CLBLM_R_X5Y105_SLICE_X7Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_A5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y106_SLICE_X6Y106_AO5),
.Q(CLBLM_R_X5Y106_SLICE_X6Y106_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_B5_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y106_SLICE_X6Y106_BO5),
.Q(CLBLM_R_X5Y106_SLICE_X6Y106_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_A_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y106_SLICE_X6Y106_AO6),
.Q(CLBLM_R_X5Y106_SLICE_X6Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_B_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y106_SLICE_X6Y106_BO6),
.Q(CLBLM_R_X5Y106_SLICE_X6Y106_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_C_FDRE (
.C(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O),
.CE(1'b1),
.D(CLBLM_R_X5Y106_SLICE_X6Y106_CO6),
.Q(CLBLM_R_X5Y106_SLICE_X6Y106_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fff7fffffffffff)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_DLUT (
.I0(CLBLM_R_X3Y106_SLICE_X2Y106_AQ),
.I1(CLBLM_R_X5Y105_SLICE_X6Y105_CQ),
.I2(CLBLM_R_X3Y107_SLICE_X2Y107_DO6),
.I3(CLBLM_R_X3Y105_SLICE_X2Y105_BQ),
.I4(1'b1),
.I5(CLBLM_R_X3Y105_SLICE_X3Y105_CO6),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_DO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h9333333333333333)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_CLUT (
.I0(CLBLM_R_X3Y106_SLICE_X2Y106_AQ),
.I1(CLBLM_R_X5Y106_SLICE_X6Y106_CQ),
.I2(CLBLM_R_X3Y107_SLICE_X2Y107_DO6),
.I3(CLBLM_R_X5Y105_SLICE_X6Y105_CQ),
.I4(CLBLM_R_X3Y105_SLICE_X3Y105_CO6),
.I5(CLBLM_R_X3Y105_SLICE_X2Y105_BQ),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_CO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hc3cccccc56aa55aa)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_BLUT (
.I0(CLBLM_R_X5Y106_SLICE_X6Y106_B5Q),
.I1(CLBLM_R_X5Y106_SLICE_X6Y106_BQ),
.I2(CLBLM_R_X5Y106_SLICE_X6Y106_CQ),
.I3(CLBLM_R_X5Y106_SLICE_X6Y106_DO6),
.I4(CLBLM_R_X5Y106_SLICE_X6Y106_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_BO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h010100000ffff000)
  ) CLBLM_R_X5Y106_SLICE_X6Y106_ALUT (
.I0(CLBLM_R_X5Y106_SLICE_X6Y106_B5Q),
.I1(CLBLM_R_X5Y106_SLICE_X6Y106_BQ),
.I2(CLBLM_R_X5Y106_SLICE_X6Y106_CQ),
.I3(CLBLM_R_X5Y106_SLICE_X6Y106_DO6),
.I4(CLBLM_R_X5Y106_SLICE_X6Y106_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X6Y106_AO5),
.O6(CLBLM_R_X5Y106_SLICE_X6Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_DO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_CO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_BO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y106_SLICE_X7Y106_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y106_SLICE_X7Y106_AO5),
.O6(CLBLM_R_X5Y106_SLICE_X7Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(LIOB33_X0Y127_IOB_X0Y128_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y101_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y101_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y101_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y101_IOB_X0Y102_IBUF (
.I(LIOB33_X0Y101_IOB_X0Y102_IPAD),
.O(LIOB33_X0Y101_IOB_X0Y102_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y103_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y103_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y103_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y103_IOB_X0Y104_IBUF (
.I(LIOB33_X0Y103_IOB_X0Y104_IPAD),
.O(LIOB33_X0Y103_IOB_X0Y104_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y105_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y105_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y105_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y105_IOB_X0Y106_IBUF (
.I(LIOB33_X0Y105_IOB_X0Y106_IPAD),
.O(LIOB33_X0Y105_IOB_X0Y106_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y107_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y107_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y107_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y107_IOB_X0Y108_IBUF (
.I(LIOB33_X0Y107_IOB_X0Y108_IPAD),
.O(LIOB33_X0Y107_IOB_X0Y108_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y109_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y109_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y109_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y109_IOB_X0Y110_IBUF (
.I(LIOB33_X0Y109_IOB_X0Y110_IPAD),
.O(LIOB33_X0Y109_IOB_X0Y110_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y111_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y111_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y111_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y111_IOB_X0Y112_IBUF (
.I(LIOB33_X0Y111_IOB_X0Y112_IPAD),
.O(LIOB33_X0Y111_IOB_X0Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y113_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y113_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y113_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y113_IOB_X0Y114_IBUF (
.I(LIOB33_X0Y113_IOB_X0Y114_IPAD),
.O(LIOB33_X0Y113_IOB_X0Y114_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y115_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y115_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y115_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y115_IOB_X0Y116_IBUF (
.I(LIOB33_X0Y115_IOB_X0Y116_IPAD),
.O(LIOB33_X0Y115_IOB_X0Y116_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y117_IOB_X0Y117_IBUF (
.I(LIOB33_X0Y117_IOB_X0Y117_IPAD),
.O(LIOB33_X0Y117_IOB_X0Y117_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y117_IOB_X0Y118_IBUF (
.I(LIOB33_X0Y117_IOB_X0Y118_IPAD),
.O(LIOB33_X0Y117_IOB_X0Y118_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y119_OBUF (
.I(CLBLL_L_X2Y110_SLICE_X0Y110_DO6),
.O(LIOB33_X0Y119_IOB_X0Y119_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y119_IOB_X0Y120_OBUF (
.I(CLBLM_R_X3Y106_SLICE_X2Y106_BO6),
.O(LIOB33_X0Y119_IOB_X0Y120_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y121_OBUF (
.I(CLBLM_R_X3Y109_SLICE_X2Y109_B5Q),
.O(LIOB33_X0Y121_IOB_X0Y121_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y121_IOB_X0Y122_OBUF (
.I(CLBLL_L_X2Y109_SLICE_X1Y109_DO5),
.O(LIOB33_X0Y121_IOB_X0Y122_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y123_OBUF (
.I(CLBLL_L_X2Y107_SLICE_X1Y107_CQ),
.O(LIOB33_X0Y123_IOB_X0Y123_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .SLEW("SLOW")
  ) LIOB33_X0Y123_IOB_X0Y124_OBUF (
.I(CLBLL_L_X2Y107_SLICE_X1Y107_CQ),
.O(LIOB33_X0Y123_IOB_X0Y124_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_X0Y127_IOB_X0Y128_IBUF (
.I(LIOB33_X0Y127_IOB_X0Y128_IPAD),
.O(LIOB33_X0Y127_IOB_X0Y128_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
  ) LIOB33_SING_X0Y100_IOB_X0Y100_IBUF (
.I(LIOB33_SING_X0Y100_IOB_X0Y100_IPAD),
.O(LIOB33_SING_X0Y100_IOB_X0Y100_I)
  );
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A = CLBLL_L_X2Y105_SLICE_X0Y105_AO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B = CLBLL_L_X2Y105_SLICE_X0Y105_BO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C = CLBLL_L_X2Y105_SLICE_X0Y105_CO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D = CLBLL_L_X2Y105_SLICE_X0Y105_DO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A = CLBLL_L_X2Y105_SLICE_X1Y105_AO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B = CLBLL_L_X2Y105_SLICE_X1Y105_BO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C = CLBLL_L_X2Y105_SLICE_X1Y105_CO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D = CLBLL_L_X2Y105_SLICE_X1Y105_DO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A = CLBLL_L_X2Y106_SLICE_X0Y106_AO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B = CLBLL_L_X2Y106_SLICE_X0Y106_BO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C = CLBLL_L_X2Y106_SLICE_X0Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D = CLBLL_L_X2Y106_SLICE_X0Y106_DO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A = CLBLL_L_X2Y106_SLICE_X1Y106_AO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B = CLBLL_L_X2Y106_SLICE_X1Y106_BO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C = CLBLL_L_X2Y106_SLICE_X1Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D = CLBLL_L_X2Y106_SLICE_X1Y106_DO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_AMUX = CLBLL_L_X2Y106_SLICE_X1Y106_A5Q;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_CMUX = CLBLL_L_X2Y106_SLICE_X1Y106_CO5;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A = CLBLL_L_X2Y107_SLICE_X0Y107_AO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B = CLBLL_L_X2Y107_SLICE_X0Y107_BO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C = CLBLL_L_X2Y107_SLICE_X0Y107_CO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D = CLBLL_L_X2Y107_SLICE_X0Y107_DO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A = CLBLL_L_X2Y107_SLICE_X1Y107_AO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B = CLBLL_L_X2Y107_SLICE_X1Y107_BO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C = CLBLL_L_X2Y107_SLICE_X1Y107_CO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D = CLBLL_L_X2Y107_SLICE_X1Y107_DO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A = CLBLL_L_X2Y108_SLICE_X0Y108_AO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B = CLBLL_L_X2Y108_SLICE_X0Y108_BO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C = CLBLL_L_X2Y108_SLICE_X0Y108_CO6;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D = CLBLL_L_X2Y108_SLICE_X0Y108_DO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A = CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B = CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C = CLBLL_L_X2Y108_SLICE_X1Y108_CO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D = CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_AMUX = CLBLL_L_X2Y108_SLICE_X1Y108_AO5;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_BMUX = CLBLL_L_X2Y108_SLICE_X1Y108_BO5;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_DMUX = CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A = CLBLL_L_X2Y109_SLICE_X0Y109_AO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B = CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C = CLBLL_L_X2Y109_SLICE_X0Y109_CO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D = CLBLL_L_X2Y109_SLICE_X0Y109_DO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_BMUX = CLBLL_L_X2Y109_SLICE_X0Y109_BO5;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A = CLBLL_L_X2Y109_SLICE_X1Y109_AO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B = CLBLL_L_X2Y109_SLICE_X1Y109_BO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C = CLBLL_L_X2Y109_SLICE_X1Y109_CO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D = CLBLL_L_X2Y109_SLICE_X1Y109_DO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_CMUX = CLBLL_L_X2Y109_SLICE_X1Y109_CO5;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_DMUX = CLBLL_L_X2Y109_SLICE_X1Y109_DO5;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A = CLBLL_L_X2Y110_SLICE_X0Y110_AO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B = CLBLL_L_X2Y110_SLICE_X0Y110_BO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C = CLBLL_L_X2Y110_SLICE_X0Y110_CO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D = CLBLL_L_X2Y110_SLICE_X0Y110_DO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A = CLBLL_L_X2Y110_SLICE_X1Y110_AO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B = CLBLL_L_X2Y110_SLICE_X1Y110_BO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C = CLBLL_L_X2Y110_SLICE_X1Y110_CO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D = CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A = CLBLL_L_X4Y104_SLICE_X4Y104_AO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B = CLBLL_L_X4Y104_SLICE_X4Y104_BO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C = CLBLL_L_X4Y104_SLICE_X4Y104_CO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D = CLBLL_L_X4Y104_SLICE_X4Y104_DO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A = CLBLL_L_X4Y104_SLICE_X5Y104_AO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B = CLBLL_L_X4Y104_SLICE_X5Y104_BO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C = CLBLL_L_X4Y104_SLICE_X5Y104_CO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D = CLBLL_L_X4Y104_SLICE_X5Y104_DO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A = CLBLL_L_X4Y105_SLICE_X4Y105_AO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B = CLBLL_L_X4Y105_SLICE_X4Y105_BO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C = CLBLL_L_X4Y105_SLICE_X4Y105_CO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D = CLBLL_L_X4Y105_SLICE_X4Y105_DO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A = CLBLL_L_X4Y105_SLICE_X5Y105_AO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C = CLBLL_L_X4Y105_SLICE_X5Y105_CO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D = CLBLL_L_X4Y105_SLICE_X5Y105_DO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A = CLBLL_L_X4Y106_SLICE_X4Y106_AO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B = CLBLL_L_X4Y106_SLICE_X4Y106_BO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C = CLBLL_L_X4Y106_SLICE_X4Y106_CO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D = CLBLL_L_X4Y106_SLICE_X4Y106_DO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A = CLBLL_L_X4Y106_SLICE_X5Y106_AO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B = CLBLL_L_X4Y106_SLICE_X5Y106_BO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C = CLBLL_L_X4Y106_SLICE_X5Y106_CO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D = CLBLL_L_X4Y106_SLICE_X5Y106_DO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A = CLBLL_L_X4Y107_SLICE_X4Y107_AO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B = CLBLL_L_X4Y107_SLICE_X4Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C = CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D = CLBLL_L_X4Y107_SLICE_X4Y107_DO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_BMUX = CLBLL_L_X4Y107_SLICE_X4Y107_B5Q;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A = CLBLL_L_X4Y107_SLICE_X5Y107_AO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B = CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C = CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D = CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_AMUX = CLBLL_L_X4Y107_SLICE_X5Y107_A5Q;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_BMUX = CLBLL_L_X4Y107_SLICE_X5Y107_BO5;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_CMUX = CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B = CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D = CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A = CLBLL_L_X4Y108_SLICE_X5Y108_AO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B = CLBLL_L_X4Y108_SLICE_X5Y108_BO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C = CLBLL_L_X4Y108_SLICE_X5Y108_CO6;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D = CLBLL_L_X4Y108_SLICE_X5Y108_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A = CLBLL_L_X4Y109_SLICE_X4Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B = CLBLL_L_X4Y109_SLICE_X4Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_AMUX = CLBLL_L_X4Y109_SLICE_X4Y109_A5Q;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_CMUX = CLBLL_L_X4Y109_SLICE_X4Y109_CO5;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_DMUX = CLBLL_L_X4Y109_SLICE_X4Y109_DO5;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A = CLBLL_L_X4Y109_SLICE_X5Y109_AO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B = CLBLL_L_X4Y109_SLICE_X5Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C = CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D = CLBLL_L_X4Y109_SLICE_X5Y109_DO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A = CLBLM_R_X3Y104_SLICE_X2Y104_AO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B = CLBLM_R_X3Y104_SLICE_X2Y104_BO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C = CLBLM_R_X3Y104_SLICE_X2Y104_CO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D = CLBLM_R_X3Y104_SLICE_X2Y104_DO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A = CLBLM_R_X3Y104_SLICE_X3Y104_AO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B = CLBLM_R_X3Y104_SLICE_X3Y104_BO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C = CLBLM_R_X3Y104_SLICE_X3Y104_CO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D = CLBLM_R_X3Y104_SLICE_X3Y104_DO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A = CLBLM_R_X3Y105_SLICE_X2Y105_AO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B = CLBLM_R_X3Y105_SLICE_X2Y105_BO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C = CLBLM_R_X3Y105_SLICE_X2Y105_CO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D = CLBLM_R_X3Y105_SLICE_X2Y105_DO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_CMUX = CLBLM_R_X3Y105_SLICE_X2Y105_CO5;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_DMUX = CLBLM_R_X3Y105_SLICE_X2Y105_DO5;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A = CLBLM_R_X3Y105_SLICE_X3Y105_AO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B = CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C = CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D = CLBLM_R_X3Y105_SLICE_X3Y105_DO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_AMUX = CLBLM_R_X3Y105_SLICE_X3Y105_A5Q;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_BMUX = CLBLM_R_X3Y105_SLICE_X3Y105_BO5;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A = CLBLM_R_X3Y106_SLICE_X2Y106_AO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B = CLBLM_R_X3Y106_SLICE_X2Y106_BO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C = CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D = CLBLM_R_X3Y106_SLICE_X2Y106_DO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_CMUX = CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A = CLBLM_R_X3Y106_SLICE_X3Y106_AO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B = CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C = CLBLM_R_X3Y106_SLICE_X3Y106_CO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D = CLBLM_R_X3Y106_SLICE_X3Y106_DO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A = CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B = CLBLM_R_X3Y107_SLICE_X2Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C = CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D = CLBLM_R_X3Y107_SLICE_X2Y107_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A = CLBLM_R_X3Y107_SLICE_X3Y107_AO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B = CLBLM_R_X3Y107_SLICE_X3Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C = CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D = CLBLM_R_X3Y107_SLICE_X3Y107_DO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A = CLBLM_R_X3Y108_SLICE_X2Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B = CLBLM_R_X3Y108_SLICE_X2Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C = CLBLM_R_X3Y108_SLICE_X2Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D = CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_CMUX = CLBLM_R_X3Y108_SLICE_X2Y108_CO5;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A = CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B = CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C = CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_AMUX = CLBLM_R_X3Y108_SLICE_X3Y108_AO5;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_BMUX = CLBLM_R_X3Y108_SLICE_X3Y108_BO5;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_CMUX = CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A = CLBLM_R_X3Y109_SLICE_X2Y109_AO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B = CLBLM_R_X3Y109_SLICE_X2Y109_BO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D = CLBLM_R_X3Y109_SLICE_X2Y109_DO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_BMUX = CLBLM_R_X3Y109_SLICE_X2Y109_B5Q;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_CMUX = CLBLM_R_X3Y109_SLICE_X2Y109_CO5;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A = CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B = CLBLM_R_X3Y109_SLICE_X3Y109_BO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C = CLBLM_R_X3Y109_SLICE_X3Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D = CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_AMUX = CLBLM_R_X3Y109_SLICE_X3Y109_AO5;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A = CLBLM_R_X3Y110_SLICE_X2Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B = CLBLM_R_X3Y110_SLICE_X2Y110_BO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C = CLBLM_R_X3Y110_SLICE_X2Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_AMUX = CLBLM_R_X3Y110_SLICE_X2Y110_A5Q;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_DMUX = CLBLM_R_X3Y110_SLICE_X2Y110_DO5;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A = CLBLM_R_X3Y110_SLICE_X3Y110_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B = CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C = CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_AMUX = CLBLM_R_X3Y110_SLICE_X3Y110_A5Q;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_CMUX = CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A = CLBLM_R_X5Y105_SLICE_X6Y105_AO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B = CLBLM_R_X5Y105_SLICE_X6Y105_BO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C = CLBLM_R_X5Y105_SLICE_X6Y105_CO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D = CLBLM_R_X5Y105_SLICE_X6Y105_DO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A = CLBLM_R_X5Y105_SLICE_X7Y105_AO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B = CLBLM_R_X5Y105_SLICE_X7Y105_BO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C = CLBLM_R_X5Y105_SLICE_X7Y105_CO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D = CLBLM_R_X5Y105_SLICE_X7Y105_DO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_AMUX = CLBLM_R_X5Y105_SLICE_X7Y105_A5Q;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_BMUX = CLBLM_R_X5Y105_SLICE_X7Y105_BO5;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A = CLBLM_R_X5Y106_SLICE_X6Y106_AO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B = CLBLM_R_X5Y106_SLICE_X6Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C = CLBLM_R_X5Y106_SLICE_X6Y106_CO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D = CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_AMUX = CLBLM_R_X5Y106_SLICE_X6Y106_A5Q;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_BMUX = CLBLM_R_X5Y106_SLICE_X6Y106_B5Q;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_DMUX = CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A = CLBLM_R_X5Y106_SLICE_X7Y106_AO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B = CLBLM_R_X5Y106_SLICE_X7Y106_BO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C = CLBLM_R_X5Y106_SLICE_X7Y106_CO6;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D = CLBLM_R_X5Y106_SLICE_X7Y106_DO6;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_O = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_O = LIOB33_X0Y101_IOB_X0Y101_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_O = LIOB33_X0Y103_IOB_X0Y104_I;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_O = LIOB33_X0Y103_IOB_X0Y103_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_O = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_O = LIOB33_X0Y105_IOB_X0Y105_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_O = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_O = LIOB33_X0Y109_IOB_X0Y109_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_O = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_O = LIOB33_X0Y111_IOB_X0Y111_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_O = LIOB33_X0Y115_IOB_X0Y116_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_O = LIOB33_X0Y115_IOB_X0Y115_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y118_O = LIOB33_X0Y117_IOB_X0Y118_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_O = LIOB33_X0Y117_IOB_X0Y117_I;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_OQ = CLBLL_L_X2Y109_SLICE_X1Y109_DO5;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_TQ = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_OQ = CLBLM_R_X3Y109_SLICE_X2Y109_B5Q;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_OQ = CLBLL_L_X2Y107_SLICE_X1Y107_CQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_TQ = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_OQ = CLBLL_L_X2Y107_SLICE_X1Y107_CQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_TQ = 1'b1;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_O = LIOB33_X0Y127_IOB_X0Y128_I;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_O = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_O = LIOB33_X0Y107_IOB_X0Y108_I;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_O = LIOB33_X0Y107_IOB_X0Y107_I;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_OQ = CLBLM_R_X3Y106_SLICE_X2Y106_BO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_OQ = CLBLL_L_X2Y110_SLICE_X0Y110_DO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_O = LIOB33_X0Y113_IOB_X0Y114_I;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_O = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C2 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C3 = CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C5 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A1 = CLBLL_L_X4Y104_SLICE_X5Y104_AQ;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A2 = CLBLL_L_X2Y106_SLICE_X0Y106_CQ;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A3 = CLBLL_L_X2Y106_SLICE_X1Y106_BQ;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A4 = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A5 = CLBLM_R_X3Y105_SLICE_X3Y105_AQ;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_A6 = CLBLL_L_X4Y104_SLICE_X5Y104_BQ;
  assign LIOB33_X0Y119_IOB_X0Y119_O = CLBLL_L_X2Y110_SLICE_X0Y110_DO6;
  assign LIOB33_X0Y119_IOB_X0Y120_O = CLBLM_R_X3Y106_SLICE_X2Y106_BO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C6 = CLBLM_R_X3Y109_SLICE_X2Y109_BQ;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B1 = CLBLM_R_X3Y105_SLICE_X3Y105_BO5;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B2 = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B3 = CLBLL_L_X4Y105_SLICE_X5Y105_DO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B4 = CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B5 = CLBLL_L_X2Y106_SLICE_X0Y106_BQ;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_B6 = CLBLL_L_X4Y105_SLICE_X4Y105_AQ;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_D1 = CLBLM_R_X3Y106_SLICE_X2Y106_BO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C1 = CLBLM_R_X3Y106_SLICE_X2Y106_AQ;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C2 = CLBLM_R_X5Y105_SLICE_X6Y105_CQ;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C3 = CLBLL_L_X2Y106_SLICE_X0Y106_DQ;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C4 = CLBLM_R_X3Y105_SLICE_X2Y105_BQ;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C5 = CLBLL_L_X2Y106_SLICE_X0Y106_CQ;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_C6 = CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y120_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_D1 = CLBLL_L_X2Y110_SLICE_X0Y110_DO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D1 = CLBLM_R_X3Y105_SLICE_X3Y105_A5Q;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D2 = CLBLL_L_X2Y106_SLICE_X0Y106_BQ;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D3 = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D4 = CLBLL_L_X4Y105_SLICE_X4Y105_AQ;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D5 = CLBLL_L_X2Y106_SLICE_X1Y106_A5Q;
  assign CLBLM_R_X3Y106_SLICE_X3Y106_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y119_OLOGIC_X0Y119_T1 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A1 = 1'b1;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A2 = CLBLM_R_X3Y105_SLICE_X2Y105_DO5;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A3 = CLBLM_R_X3Y106_SLICE_X2Y106_AQ;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_A6 = CLBLM_R_X3Y105_SLICE_X2Y105_BQ;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B1 = CLBLM_R_X3Y106_SLICE_X2Y106_AQ;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B2 = CLBLM_R_X3Y105_SLICE_X2Y105_DO5;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B3 = CLBLM_R_X3Y106_SLICE_X3Y106_AO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B4 = CLBLL_L_X2Y106_SLICE_X1Y106_DO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B5 = CLBLL_L_X2Y106_SLICE_X0Y106_AQ;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_B6 = CLBLM_R_X3Y105_SLICE_X2Y105_BQ;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C1 = CLBLL_L_X4Y105_SLICE_X4Y105_AQ;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C2 = CLBLL_L_X2Y106_SLICE_X0Y106_BQ;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C3 = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C4 = CLBLM_R_X3Y105_SLICE_X3Y105_A5Q;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C5 = CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_C6 = CLBLL_L_X2Y106_SLICE_X1Y106_A5Q;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D1 = CLBLL_L_X4Y105_SLICE_X5Y105_DO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D2 = CLBLL_L_X4Y105_SLICE_X4Y105_AQ;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D3 = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D4 = CLBLL_L_X2Y106_SLICE_X0Y106_BQ;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D5 = CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  assign CLBLM_R_X3Y106_SLICE_X2Y106_D6 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I0 = LIOB33_X0Y127_IOB_X0Y128_I;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign LIOB33_X0Y121_IOB_X0Y122_O = CLBLL_L_X2Y109_SLICE_X1Y109_DO5;
  assign LIOB33_X0Y121_IOB_X0Y121_O = CLBLM_R_X3Y109_SLICE_X2Y109_B5Q;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A1 = CLBLM_R_X3Y107_SLICE_X3Y107_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A4 = CLBLM_R_X3Y107_SLICE_X3Y107_BO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A5 = CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_A6 = CLBLM_R_X3Y107_SLICE_X3Y107_CO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B1 = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B2 = CLBLM_R_X3Y106_SLICE_X2Y106_AQ;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B3 = CLBLL_L_X2Y105_SLICE_X1Y105_AQ;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B4 = CLBLL_L_X2Y106_SLICE_X0Y106_CQ;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B5 = CLBLL_L_X2Y106_SLICE_X0Y106_DQ;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_B6 = CLBLM_R_X3Y108_SLICE_X3Y108_AO5;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C1 = CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C2 = CLBLM_R_X3Y106_SLICE_X3Y106_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C3 = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C4 = CLBLL_L_X2Y109_SLICE_X1Y109_BQ;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C5 = CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_C6 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B6 = CLBLL_L_X4Y107_SLICE_X4Y107_AQ;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D2 = CLBLM_R_X3Y106_SLICE_X3Y106_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D3 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D4 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D5 = CLBLL_L_X4Y108_SLICE_X4Y108_DO6;
  assign CLBLM_R_X3Y107_SLICE_X3Y107_D6 = CLBLL_L_X2Y106_SLICE_X0Y106_CQ;
  assign LIOI3_X0Y103_ILOGIC_X0Y103_D = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A1 = CLBLM_R_X3Y108_SLICE_X2Y108_BQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A3 = CLBLM_R_X3Y107_SLICE_X2Y107_AQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A4 = CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_A6 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B1 = CLBLM_R_X3Y108_SLICE_X2Y108_BQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B2 = CLBLL_L_X2Y106_SLICE_X0Y106_CQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B3 = CLBLL_L_X2Y109_SLICE_X1Y109_BQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B5 = CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_B6 = CLBLL_L_X2Y107_SLICE_X1Y107_AQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C1 = CLBLL_L_X4Y109_SLICE_X5Y109_BQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C2 = CLBLM_R_X3Y105_SLICE_X3Y105_DO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C3 = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C4 = CLBLM_R_X3Y105_SLICE_X3Y105_A5Q;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C5 = CLBLM_R_X3Y106_SLICE_X2Y106_DO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_C6 = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C6 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D1 = CLBLL_L_X4Y106_SLICE_X4Y106_AQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D2 = CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D3 = CLBLM_R_X3Y105_SLICE_X3Y105_DO6;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D4 = 1'b1;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D5 = CLBLM_R_X3Y109_SLICE_X2Y109_AQ;
  assign CLBLM_R_X3Y107_SLICE_X2Y107_D6 = CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C6 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B6 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_D = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_ILOGIC_X0Y111_D = LIOB33_X0Y111_IOB_X0Y111_I;
  assign LIOB33_X0Y123_IOB_X0Y124_O = CLBLL_L_X2Y107_SLICE_X1Y107_CQ;
  assign LIOB33_X0Y123_IOB_X0Y123_O = CLBLL_L_X2Y107_SLICE_X1Y107_CQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A1 = CLBLL_L_X4Y106_SLICE_X5Y106_DO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A3 = CLBLM_R_X5Y105_SLICE_X7Y105_AQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A4 = CLBLL_L_X4Y106_SLICE_X5Y106_BQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A5 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_A6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_AX = CLBLM_R_X5Y105_SLICE_X7Y105_BO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B1 = CLBLL_L_X4Y106_SLICE_X5Y106_DO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B2 = CLBLM_R_X5Y105_SLICE_X7Y105_A5Q;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B3 = CLBLM_R_X5Y105_SLICE_X7Y105_AQ;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_B6 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B4 = CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A1 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A2 = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A4 = CLBLL_L_X2Y106_SLICE_X1Y106_A5Q;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A5 = CLBLL_L_X2Y106_SLICE_X0Y106_CQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_A6 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C1 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C2 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C3 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B1 = CLBLL_L_X2Y106_SLICE_X0Y106_CQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B2 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B3 = CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B4 = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B5 = CLBLM_R_X3Y109_SLICE_X2Y109_AQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_B6 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D1 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D4 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C1 = CLBLM_R_X3Y109_SLICE_X2Y109_AQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C2 = CLBLM_R_X3Y109_SLICE_X3Y109_AO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C3 = CLBLL_L_X2Y108_SLICE_X1Y108_CO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C4 = CLBLM_R_X3Y110_SLICE_X2Y110_A5Q;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C5 = CLBLM_R_X3Y108_SLICE_X3Y108_BO5;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_C6 = CLBLL_L_X2Y108_SLICE_X1Y108_DO6;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D6 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A1 = CLBLM_R_X3Y105_SLICE_X2Y105_DO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A2 = CLBLM_R_X5Y105_SLICE_X6Y105_DO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A3 = CLBLM_R_X5Y105_SLICE_X6Y105_AQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D1 = CLBLM_R_X3Y108_SLICE_X2Y108_AQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D2 = CLBLL_L_X2Y109_SLICE_X1Y109_BQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D3 = CLBLL_L_X2Y110_SLICE_X1Y110_DO6;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D4 = CLBLL_L_X2Y106_SLICE_X0Y106_CQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B1 = CLBLM_R_X3Y105_SLICE_X2Y105_DO6;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B2 = CLBLM_R_X5Y105_SLICE_X6Y105_BQ;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X3Y108_D6 = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B3 = CLBLM_R_X5Y105_SLICE_X6Y105_AQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C2 = CLBLM_R_X5Y106_SLICE_X6Y106_CQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A1 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A2 = CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A3 = CLBLM_R_X3Y108_SLICE_X2Y108_AQ;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A4 = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A5 = CLBLM_R_X3Y107_SLICE_X2Y107_AQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_B6 = CLBLM_R_X5Y105_SLICE_X6Y105_CQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C1 = CLBLM_R_X5Y105_SLICE_X6Y105_BQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C5 = CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B1 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B2 = CLBLM_R_X3Y108_SLICE_X2Y108_BQ;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B3 = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B4 = CLBLL_L_X4Y106_SLICE_X4Y106_AQ;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B5 = CLBLL_L_X4Y108_SLICE_X4Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D1 = CLBLL_L_X2Y106_SLICE_X0Y106_DQ;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C1 = CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C2 = CLBLL_L_X4Y109_SLICE_X5Y109_BQ;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C3 = CLBLM_R_X3Y110_SLICE_X2Y110_A5Q;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C5 = CLBLL_L_X2Y106_SLICE_X0Y106_CQ;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_C6 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D2 = CLBLM_R_X5Y105_SLICE_X6Y105_CQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D4 = CLBLM_R_X5Y106_SLICE_X6Y106_AQ;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_D6 = CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D1 = CLBLM_R_X3Y108_SLICE_X2Y108_CO5;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D2 = CLBLM_R_X3Y109_SLICE_X2Y109_AQ;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D3 = CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D4 = CLBLM_R_X3Y110_SLICE_X2Y110_A5Q;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D5 = 1'b1;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_D6 = CLBLM_R_X3Y109_SLICE_X2Y109_CO5;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D1 = CLBLM_R_X3Y106_SLICE_X2Y106_AQ;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C6 = CLBLL_L_X2Y106_SLICE_X0Y106_BQ;
  assign CLBLM_R_X3Y108_SLICE_X2Y108_A6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D3 = CLBLM_R_X3Y107_SLICE_X2Y107_DO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y127_ILOGIC_X0Y128_D = LIOB33_X0Y127_IOB_X0Y128_I;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A1 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A2 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A3 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A4 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A5 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_A6 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B1 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B2 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B3 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B4 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B5 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_B6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A1 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A2 = CLBLM_R_X3Y110_SLICE_X2Y110_AQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A3 = CLBLL_L_X2Y106_SLICE_X0Y106_CQ;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C3 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C4 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A5 = CLBLL_L_X4Y109_SLICE_X5Y109_BQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_A6 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C1 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_C2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B1 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B2 = CLBLM_R_X3Y109_SLICE_X3Y109_BQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B3 = CLBLM_R_X3Y108_SLICE_X2Y108_AQ;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D1 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D2 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D3 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D4 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D5 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X7Y106_D6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B4 = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B5 = CLBLM_R_X3Y106_SLICE_X3Y106_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C1 = CLBLL_L_X2Y109_SLICE_X0Y109_BO5;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_C2 = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A1 = CLBLM_R_X5Y106_SLICE_X6Y106_B5Q;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A2 = CLBLM_R_X5Y106_SLICE_X6Y106_BQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A3 = CLBLM_R_X5Y106_SLICE_X6Y106_CQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A4 = CLBLM_R_X5Y106_SLICE_X6Y106_DO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A5 = CLBLM_R_X5Y106_SLICE_X6Y106_A5Q;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D1 = CLBLM_R_X3Y110_SLICE_X2Y110_CQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D2 = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D3 = CLBLM_R_X3Y108_SLICE_X2Y108_DO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D4 = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D5 = CLBLM_R_X3Y110_SLICE_X2Y110_BQ;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_D6 = CLBLL_L_X2Y109_SLICE_X1Y109_DO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_A6 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B5 = CLBLM_R_X5Y106_SLICE_X6Y106_A5Q;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B1 = CLBLM_R_X5Y106_SLICE_X6Y106_B5Q;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B2 = CLBLM_R_X5Y106_SLICE_X6Y106_BQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_B3 = CLBLM_R_X5Y106_SLICE_X6Y106_CQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A1 = CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A3 = CLBLM_R_X3Y109_SLICE_X2Y109_AQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A4 = CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A5 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C3 = CLBLM_R_X3Y107_SLICE_X2Y107_DO6;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C4 = CLBLM_R_X5Y105_SLICE_X6Y105_CQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_A6 = CLBLL_L_X4Y104_SLICE_X5Y104_BQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C1 = CLBLM_R_X3Y106_SLICE_X2Y106_AQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B1 = CLBLM_R_X3Y109_SLICE_X2Y109_DO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B2 = CLBLM_R_X3Y110_SLICE_X3Y110_A5Q;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B3 = CLBLM_R_X3Y107_SLICE_X3Y107_AO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B5 = CLBLL_L_X2Y106_SLICE_X0Y106_BQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_B6 = 1'b1;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_C6 = CLBLM_R_X3Y105_SLICE_X2Y105_BQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D2 = CLBLM_R_X5Y105_SLICE_X6Y105_CQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D4 = CLBLM_R_X3Y105_SLICE_X2Y105_BQ;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D5 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X5Y106_SLICE_X6Y106_D6 = CLBLM_R_X3Y105_SLICE_X3Y105_CO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C5 = CLBLL_L_X2Y106_SLICE_X0Y106_CQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C1 = CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C2 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C4 = CLBLM_R_X3Y110_SLICE_X2Y110_AQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_C6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D2 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D3 = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D4 = CLBLL_L_X4Y106_SLICE_X4Y106_AQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D5 = CLBLM_R_X3Y109_SLICE_X2Y109_BQ;
  assign CLBLM_R_X3Y109_SLICE_X2Y109_D6 = CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A1 = CLBLM_R_X3Y110_SLICE_X3Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A3 = CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A4 = CLBLM_R_X3Y110_SLICE_X3Y110_AQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A5 = CLBLM_R_X3Y110_SLICE_X3Y110_CO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_A6 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B1 = CLBLM_R_X3Y109_SLICE_X3Y109_BQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B2 = CLBLM_R_X3Y109_SLICE_X2Y109_BQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B3 = CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B4 = CLBLM_R_X3Y110_SLICE_X3Y110_AQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_B6 = CLBLM_R_X3Y110_SLICE_X3Y110_A5Q;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C1 = CLBLL_L_X4Y106_SLICE_X4Y106_AQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C2 = CLBLM_R_X3Y110_SLICE_X3Y110_AQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C3 = CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C4 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_C6 = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_X0Y115_ILOGIC_X0Y116_D = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign LIOI3_X0Y115_ILOGIC_X0Y115_D = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D1 = CLBLL_L_X4Y106_SLICE_X4Y106_AQ;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D2 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D4 = CLBLM_R_X3Y110_SLICE_X3Y110_A5Q;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D5 = CLBLM_R_X3Y108_SLICE_X3Y108_AO6;
  assign CLBLM_R_X3Y110_SLICE_X3Y110_D6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C1 = CLBLM_R_X3Y109_SLICE_X3Y109_AO5;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A2 = CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A3 = CLBLM_R_X3Y110_SLICE_X2Y110_AQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A4 = CLBLM_R_X3Y110_SLICE_X2Y110_DO5;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A5 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_A6 = CLBLM_R_X3Y110_SLICE_X2Y110_A5Q;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_AX = CLBLM_R_X3Y110_SLICE_X2Y110_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B1 = 1'b1;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B2 = CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C4 = CLBLL_L_X4Y109_SLICE_X4Y109_DO5;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B4 = CLBLM_R_X3Y110_SLICE_X2Y110_DO5;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B5 = CLBLM_R_X3Y110_SLICE_X2Y110_BQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_B3 = CLBLM_R_X3Y110_SLICE_X2Y110_AQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C1 = CLBLM_R_X3Y110_SLICE_X2Y110_BQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C6 = CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C2 = CLBLM_R_X3Y110_SLICE_X2Y110_AQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C4 = CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C5 = CLBLM_R_X3Y110_SLICE_X2Y110_CQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_C6 = CLBLM_R_X3Y110_SLICE_X2Y110_DO5;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D1 = CLBLM_R_X3Y109_SLICE_X2Y109_AQ;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D3 = CLBLL_L_X2Y109_SLICE_X0Y109_BO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D4 = CLBLM_R_X3Y110_SLICE_X2Y110_A5Q;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D5 = CLBLL_L_X4Y107_SLICE_X5Y107_DO6;
  assign CLBLM_R_X3Y110_SLICE_X2Y110_D6 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B5 = CLBLL_L_X2Y106_SLICE_X0Y106_BQ;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A3 = CLBLL_L_X4Y104_SLICE_X4Y104_AQ;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A4 = CLBLL_L_X4Y104_SLICE_X5Y104_CO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A5 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_A6 = CLBLL_L_X2Y106_SLICE_X1Y106_A5Q;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B1 = CLBLM_R_X5Y105_SLICE_X6Y105_CQ;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B2 = CLBLL_L_X4Y104_SLICE_X4Y104_BQ;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B4 = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B5 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C1 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C2 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C3 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C4 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C5 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_C6 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D1 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D2 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D3 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D4 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D5 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X4Y104_D6 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A1 = CLBLM_R_X3Y105_SLICE_X3Y105_AQ;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A3 = CLBLL_L_X4Y104_SLICE_X5Y104_AQ;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A4 = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A5 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_A6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_I = CLK_BUFG_BOT_R_X139Y152_BUFGCTRL_X0Y0_O;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B1 = CLBLM_R_X3Y105_SLICE_X3Y105_AQ;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B2 = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B3 = CLBLL_L_X4Y104_SLICE_X5Y104_AQ;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B5 = CLBLL_L_X4Y104_SLICE_X5Y104_BQ;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C1 = CLBLL_L_X4Y104_SLICE_X5Y104_BQ;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C2 = CLBLL_L_X2Y106_SLICE_X0Y106_DQ;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C3 = CLBLM_R_X3Y105_SLICE_X3Y105_AQ;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C4 = CLBLL_L_X4Y104_SLICE_X5Y104_AQ;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C5 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_C6 = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D1 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D2 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D3 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D4 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D5 = 1'b1;
  assign CLBLL_L_X4Y104_SLICE_X5Y104_D6 = 1'b1;
  assign LIOI3_X0Y101_ILOGIC_X0Y102_D = LIOB33_X0Y101_IOB_X0Y102_I;
  assign LIOI3_X0Y101_ILOGIC_X0Y101_D = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A1 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A2 = CLBLL_L_X4Y105_SLICE_X5Y105_DO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A3 = CLBLL_L_X4Y105_SLICE_X4Y105_AQ;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A5 = CLBLL_L_X4Y105_SLICE_X5Y105_AQ;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_A6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B1 = CLBLM_R_X3Y104_SLICE_X3Y104_DO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B2 = CLBLL_L_X4Y105_SLICE_X4Y105_BQ;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B3 = CLBLM_R_X3Y104_SLICE_X3Y104_AQ;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B4 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C2 = CLBLL_L_X4Y105_SLICE_X4Y105_CQ;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C3 = CLBLM_R_X3Y104_SLICE_X3Y104_DO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C4 = CLBLL_L_X4Y105_SLICE_X4Y105_BQ;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C5 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_C6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D2 = CLBLL_L_X4Y105_SLICE_X4Y105_CQ;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D3 = CLBLL_L_X4Y105_SLICE_X4Y105_DQ;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D4 = CLBLM_R_X3Y104_SLICE_X3Y104_DO6;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D5 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X4Y105_D6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A1 = CLBLL_L_X4Y106_SLICE_X5Y106_DO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A2 = CLBLM_R_X5Y105_SLICE_X7Y105_A5Q;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A3 = CLBLL_L_X4Y105_SLICE_X5Y105_AQ;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A4 = CLBLM_R_X5Y105_SLICE_X7Y105_AQ;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_A6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B1 = CLBLL_L_X4Y106_SLICE_X5Y106_DO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B2 = CLBLM_R_X5Y105_SLICE_X7Y105_A5Q;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B3 = CLBLL_L_X4Y105_SLICE_X5Y105_AQ;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B4 = CLBLM_R_X5Y105_SLICE_X7Y105_AQ;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B5 = CLBLL_L_X4Y105_SLICE_X4Y105_AQ;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_B6 = CLBLL_L_X2Y106_SLICE_X0Y106_BQ;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C1 = CLBLL_L_X4Y105_SLICE_X4Y105_AQ;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C2 = CLBLM_R_X3Y105_SLICE_X3Y105_AQ;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C3 = CLBLL_L_X4Y106_SLICE_X5Y106_CO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C4 = CLBLL_L_X4Y105_SLICE_X5Y105_AQ;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C5 = CLBLL_L_X4Y104_SLICE_X5Y104_AQ;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_C6 = CLBLL_L_X2Y106_SLICE_X0Y106_BQ;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D1 = CLBLM_R_X5Y105_SLICE_X7Y105_AQ;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D2 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D3 = CLBLL_L_X4Y106_SLICE_X5Y106_DO6;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D4 = 1'b1;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D5 = CLBLL_L_X4Y105_SLICE_X5Y105_AQ;
  assign CLBLL_L_X4Y105_SLICE_X5Y105_D6 = CLBLM_R_X5Y105_SLICE_X7Y105_A5Q;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B5 = CLBLL_L_X4Y106_SLICE_X4Y106_BQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B6 = 1'b1;
  assign LIOI3_X0Y117_ILOGIC_X0Y118_D = LIOB33_X0Y117_IOB_X0Y118_I;
  assign LIOI3_X0Y117_ILOGIC_X0Y117_D = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A1 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A3 = CLBLL_L_X4Y106_SLICE_X4Y106_AQ;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A4 = CLBLM_R_X3Y106_SLICE_X2Y106_AQ;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_A6 = CLBLM_R_X3Y106_SLICE_X3Y106_DO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B1 = CLBLL_L_X4Y106_SLICE_X4Y106_BQ;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B3 = CLBLL_L_X4Y107_SLICE_X5Y107_AQ;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B4 = CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A1 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A2 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A3 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A4 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A5 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_A6 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_B5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C2 = CLBLL_L_X4Y106_SLICE_X4Y106_CQ;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C3 = CLBLL_L_X4Y107_SLICE_X4Y107_B5Q;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B1 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B2 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B3 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B4 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B5 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_B6 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C4 = CLBLL_L_X4Y107_SLICE_X4Y107_DO6;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_C5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C1 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C2 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C3 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C4 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C5 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_C6 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D1 = CLBLL_L_X4Y107_SLICE_X5Y107_AQ;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D2 = CLBLL_L_X4Y106_SLICE_X4Y106_CQ;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D3 = CLBLL_L_X4Y107_SLICE_X4Y107_B5Q;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D4 = CLBLL_L_X4Y107_SLICE_X4Y107_AQ;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D5 = CLBLL_L_X4Y106_SLICE_X4Y106_BQ;
  assign CLBLL_L_X4Y106_SLICE_X4Y106_D6 = CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D1 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D2 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D3 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D4 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D5 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X0Y105_D6 = 1'b1;
  assign CLBLM_R_X3Y109_SLICE_X3Y109_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A1 = CLBLL_L_X4Y106_SLICE_X5Y106_AQ;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A2 = CLBLL_L_X2Y106_SLICE_X0Y106_BQ;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A4 = CLBLL_L_X4Y106_SLICE_X4Y106_DO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_A6 = CLBLL_L_X4Y106_SLICE_X4Y106_CQ;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B1 = CLBLL_L_X4Y106_SLICE_X5Y106_AQ;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B2 = CLBLL_L_X4Y106_SLICE_X5Y106_BQ;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_B4 = CLBLL_L_X4Y106_SLICE_X4Y106_DO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A2 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A3 = CLBLL_L_X2Y105_SLICE_X1Y105_AQ;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A4 = CLBLM_R_X3Y105_SLICE_X2Y105_CO5;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A5 = CLBLM_R_X3Y104_SLICE_X2Y104_BQ;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_A6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C1 = CLBLL_L_X4Y106_SLICE_X5Y106_BQ;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C2 = CLBLL_L_X4Y107_SLICE_X4Y107_DO6;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B1 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B2 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B3 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B4 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B5 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_B6 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C3 = CLBLL_L_X4Y106_SLICE_X5Y106_AQ;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C4 = CLBLL_L_X4Y106_SLICE_X4Y106_CQ;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_C5 = CLBLM_R_X5Y105_SLICE_X7Y105_BO5;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C1 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C2 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C3 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C4 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C5 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_C6 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D1 = CLBLL_L_X4Y106_SLICE_X5Y106_BQ;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D2 = CLBLL_L_X4Y107_SLICE_X4Y107_DO6;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D3 = 1'b1;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D4 = CLBLL_L_X4Y106_SLICE_X4Y106_CQ;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D5 = CLBLL_L_X4Y106_SLICE_X5Y106_AQ;
  assign CLBLL_L_X4Y106_SLICE_X5Y106_D6 = CLBLL_L_X2Y106_SLICE_X0Y106_BQ;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D1 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D2 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D3 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D4 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D5 = 1'b1;
  assign CLBLL_L_X2Y105_SLICE_X1Y105_D6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C2 = CLBLM_R_X3Y106_SLICE_X3Y106_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A2 = CLBLL_L_X4Y107_SLICE_X4Y107_AQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A4 = CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A5 = CLBLL_L_X4Y107_SLICE_X5Y107_AQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_A6 = 1'b1;
  assign LIOI3_X0Y103_ILOGIC_X0Y104_D = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B2 = CLBLL_L_X4Y107_SLICE_X4Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B3 = CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_B4 = LIOB33_X0Y117_IOB_X0Y118_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A1 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A3 = CLBLL_L_X2Y106_SLICE_X0Y106_AQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A4 = CLBLL_L_X2Y106_SLICE_X1Y106_BQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C1 = CLBLL_L_X4Y107_SLICE_X5Y107_AQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C2 = CLBLL_L_X4Y107_SLICE_X4Y107_AQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C3 = CLBLM_R_X3Y107_SLICE_X2Y107_AO6;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C4 = CLBLL_L_X4Y106_SLICE_X4Y106_BQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C5 = CLBLL_L_X4Y107_SLICE_X4Y107_B5Q;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_C6 = CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_A6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B1 = CLBLL_L_X2Y106_SLICE_X1Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B3 = CLBLL_L_X2Y106_SLICE_X0Y106_DQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C1 = CLBLL_L_X2Y106_SLICE_X0Y106_CQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D1 = CLBLL_L_X4Y107_SLICE_X5Y107_AQ;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D2 = CLBLL_L_X4Y107_SLICE_X4Y107_AQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C2 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D3 = CLBLL_L_X2Y109_SLICE_X1Y109_CO5;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D4 = CLBLL_L_X4Y108_SLICE_X4Y108_CO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D6 = CLBLL_L_X4Y106_SLICE_X4Y106_BQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C4 = CLBLL_L_X2Y107_SLICE_X0Y107_AQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C5 = CLBLL_L_X2Y106_SLICE_X1Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_C6 = CLBLL_L_X2Y106_SLICE_X0Y106_AQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y107_SLICE_X4Y107_D5 = CLBLL_L_X4Y107_SLICE_X4Y107_B5Q;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D2 = CLBLL_L_X2Y106_SLICE_X0Y106_CQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D3 = CLBLL_L_X2Y106_SLICE_X0Y106_DQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D4 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D5 = CLBLL_L_X2Y106_SLICE_X1Y106_CO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_D6 = CLBLL_L_X2Y107_SLICE_X0Y107_AQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A1 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A2 = CLBLM_R_X3Y109_SLICE_X3Y109_DO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A3 = CLBLL_L_X4Y107_SLICE_X5Y107_AQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_A6 = CLBLL_L_X4Y107_SLICE_X5Y107_A5Q;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_AX = CLBLL_L_X4Y107_SLICE_X5Y107_BO5;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B1 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B2 = CLBLL_L_X4Y107_SLICE_X5Y107_A5Q;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B4 = CLBLL_L_X4Y107_SLICE_X4Y107_BQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B5 = CLBLL_L_X4Y107_SLICE_X5Y107_CO6;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_B6 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A1 = CLBLL_L_X2Y107_SLICE_X1Y107_DQ;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A2 = CLBLL_L_X2Y107_SLICE_X0Y107_AQ;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A3 = CLBLL_L_X2Y106_SLICE_X1Y106_AQ;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A5 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_A6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C1 = CLBLL_L_X4Y105_SLICE_X4Y105_BQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C2 = CLBLL_L_X4Y105_SLICE_X4Y105_CQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C4 = CLBLM_R_X3Y104_SLICE_X3Y104_AQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C5 = CLBLL_L_X4Y105_SLICE_X4Y105_DQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_C6 = CLBLL_L_X4Y107_SLICE_X4Y107_BQ;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_AX = CLBLL_L_X2Y106_SLICE_X1Y106_CO5;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B1 = CLBLL_L_X2Y106_SLICE_X1Y106_AQ;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B2 = CLBLL_L_X2Y106_SLICE_X1Y106_BQ;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B3 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_B5 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D1 = CLBLL_L_X4Y105_SLICE_X4Y105_BQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D2 = CLBLL_L_X4Y105_SLICE_X4Y105_CQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D3 = 1'b1;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D4 = CLBLL_L_X4Y105_SLICE_X4Y105_DQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D5 = CLBLM_R_X3Y104_SLICE_X3Y104_AQ;
  assign CLBLL_L_X4Y107_SLICE_X5Y107_D6 = CLBLL_L_X4Y107_SLICE_X5Y107_BO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C1 = CLBLL_L_X4Y105_SLICE_X4Y105_AQ;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C4 = CLBLL_L_X2Y106_SLICE_X1Y106_A5Q;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_C6 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D1 = 1'b1;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D2 = CLBLL_L_X4Y105_SLICE_X5Y105_DO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D3 = CLBLL_L_X4Y106_SLICE_X4Y106_DO6;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D4 = CLBLL_L_X2Y106_SLICE_X1Y106_AQ;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D5 = CLBLL_L_X2Y107_SLICE_X1Y107_DQ;
  assign CLBLL_L_X2Y106_SLICE_X1Y106_D6 = CLBLL_L_X4Y105_SLICE_X4Y105_AQ;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_D1 = CLBLL_L_X2Y109_SLICE_X1Y109_DO5;
  assign LIOI3_X0Y121_OLOGIC_X0Y122_T1 = 1'b1;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_D1 = CLBLM_R_X3Y109_SLICE_X2Y109_B5Q;
  assign LIOI3_X0Y121_OLOGIC_X0Y121_T1 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A1 = CLBLM_R_X3Y110_SLICE_X3Y110_A5Q;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A2 = CLBLL_L_X4Y109_SLICE_X4Y109_A5Q;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A3 = CLBLL_L_X4Y109_SLICE_X4Y109_BQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A4 = CLBLM_R_X3Y109_SLICE_X2Y109_BQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_A6 = CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B1 = CLBLM_R_X3Y110_SLICE_X3Y110_A5Q;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B2 = CLBLL_L_X4Y109_SLICE_X4Y109_A5Q;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B4 = CLBLM_R_X3Y109_SLICE_X2Y109_BQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B5 = CLBLL_L_X4Y109_SLICE_X4Y109_BQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_B6 = CLBLM_R_X3Y110_SLICE_X3Y110_BO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A1 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A3 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C1 = CLBLM_R_X3Y110_SLICE_X2Y110_BQ;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C2 = CLBLL_L_X4Y109_SLICE_X5Y109_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C3 = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C4 = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C5 = CLBLL_L_X2Y109_SLICE_X1Y109_CO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_C6 = CLBLM_R_X3Y108_SLICE_X3Y108_CO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A4 = CLBLL_L_X2Y107_SLICE_X1Y107_BQ;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_A6 = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_B6 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D4 = CLBLM_R_X3Y109_SLICE_X2Y109_CO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C1 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D6 = CLBLM_R_X3Y108_SLICE_X2Y108_CO6;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_C6 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D1 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D3 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X0Y107_D6 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A1 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A2 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A3 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A4 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A5 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_A6 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B1 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B2 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B3 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B4 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A1 = LIOB33_X0Y101_IOB_X0Y102_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A2 = CLBLL_L_X2Y109_SLICE_X1Y109_BQ;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A3 = CLBLL_L_X2Y107_SLICE_X1Y107_AQ;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A5 = CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_A6 = CLBLL_L_X2Y108_SLICE_X1Y108_AO5;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B5 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_B6 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B1 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B2 = CLBLL_L_X2Y107_SLICE_X1Y107_BQ;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B3 = CLBLL_L_X2Y107_SLICE_X1Y107_AQ;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B5 = CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_B6 = CLBLL_L_X2Y108_SLICE_X1Y108_AO5;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C3 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C4 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C1 = CLBLM_R_X3Y107_SLICE_X2Y107_BO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C2 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C3 = CLBLL_L_X2Y107_SLICE_X1Y107_DQ;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C4 = CLBLM_R_X3Y106_SLICE_X3Y106_DO6;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C5 = CLBLL_L_X2Y108_SLICE_X1Y108_BO5;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_C6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D4 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D5 = 1'b1;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D6 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D2 = 1'b1;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D3 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C3 = CLBLM_R_X3Y109_SLICE_X3Y109_BQ;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D1 = CLBLL_L_X2Y106_SLICE_X0Y106_AQ;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D3 = CLBLL_L_X2Y107_SLICE_X1Y107_DQ;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D4 = LIOB33_X0Y103_IOB_X0Y103_I;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D5 = CLBLM_R_X3Y109_SLICE_X2Y109_B5Q;
  assign CLBLL_L_X2Y107_SLICE_X1Y107_D6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C4 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C5 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_C6 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D2 = 1'b1;
  assign CLBLM_R_X5Y105_SLICE_X7Y105_D3 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A2 = CLBLL_L_X4Y109_SLICE_X4Y109_BQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A3 = CLBLL_L_X4Y109_SLICE_X4Y109_AQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A4 = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A5 = CLBLL_L_X4Y109_SLICE_X4Y109_CO5;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_A6 = CLBLM_R_X3Y106_SLICE_X3Y106_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_AX = CLBLL_L_X4Y109_SLICE_X4Y109_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B2 = CLBLL_L_X4Y109_SLICE_X4Y109_BQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B3 = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B4 = CLBLM_R_X3Y109_SLICE_X3Y109_BQ;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A1 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A3 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_A6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C1 = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B5 = CLBLL_L_X4Y109_SLICE_X4Y109_A5Q;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_B6 = CLBLM_R_X3Y106_SLICE_X3Y106_CO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C4 = CLBLL_L_X4Y109_SLICE_X4Y109_A5Q;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_C6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B3 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_B6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C1 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C3 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_C6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D1 = CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D2 = LIOB33_X0Y109_IOB_X0Y110_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D3 = CLBLL_L_X2Y109_SLICE_X0Y109_AQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D4 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D5 = CLBLL_L_X2Y106_SLICE_X0Y106_CQ;
  assign CLBLL_L_X4Y109_SLICE_X4Y109_D6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D1 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D2 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D3 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D4 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X0Y108_D6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A1 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A2 = CLBLL_L_X4Y109_SLICE_X5Y109_BQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A3 = CLBLL_L_X2Y109_SLICE_X0Y109_BO5;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A4 = CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A5 = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_A6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_A6 = CLBLL_L_X4Y105_SLICE_X4Y105_DQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B2 = CLBLL_L_X4Y109_SLICE_X5Y109_BQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B3 = CLBLL_L_X2Y109_SLICE_X0Y109_BO5;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B4 = CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A1 = CLBLL_L_X2Y106_SLICE_X0Y106_DQ;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A4 = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A5 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_A6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B5 = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B1 = CLBLM_R_X3Y108_SLICE_X2Y108_BQ;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B2 = CLBLL_L_X2Y107_SLICE_X1Y107_BQ;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B3 = CLBLL_L_X2Y107_SLICE_X1Y107_AQ;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B5 = CLBLL_L_X2Y106_SLICE_X0Y106_CQ;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_B6 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C2 = CLBLM_R_X3Y110_SLICE_X2Y110_A5Q;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C3 = CLBLL_L_X4Y109_SLICE_X5Y109_BQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_C5 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C1 = CLBLL_L_X2Y107_SLICE_X1Y107_AQ;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C2 = CLBLM_R_X3Y108_SLICE_X2Y108_BQ;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C3 = CLBLL_L_X2Y106_SLICE_X0Y106_CQ;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C5 = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_C6 = CLBLL_L_X2Y107_SLICE_X1Y107_BQ;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D1 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D2 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D3 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D4 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D5 = 1'b1;
  assign CLBLL_L_X4Y109_SLICE_X5Y109_D6 = 1'b1;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D1 = CLBLL_L_X2Y107_SLICE_X1Y107_AQ;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D2 = CLBLM_R_X3Y108_SLICE_X2Y108_BQ;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D3 = CLBLL_L_X2Y106_SLICE_X0Y106_CQ;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D4 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D5 = LIOB33_X0Y101_IOB_X0Y101_I;
  assign CLBLL_L_X2Y108_SLICE_X1Y108_D6 = CLBLL_L_X2Y107_SLICE_X1Y107_BQ;
  assign LIOI3_X0Y105_ILOGIC_X0Y106_D = LIOB33_X0Y105_IOB_X0Y106_I;
  assign LIOI3_X0Y105_ILOGIC_X0Y105_D = LIOB33_X0Y105_IOB_X0Y105_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C2 = CLBLM_R_X5Y105_SLICE_X6Y105_AQ;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y114_D = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C3 = CLBLM_R_X3Y105_SLICE_X2Y105_DO6;
  assign LIOI3_TBYTETERM_X0Y113_ILOGIC_X0Y113_D = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C4 = CLBLM_R_X5Y105_SLICE_X6Y105_CQ;
  assign CLBLM_R_X5Y105_SLICE_X6Y105_C5 = CLBLM_R_X5Y105_SLICE_X6Y105_DO6;
  assign LIOI3_SING_X0Y100_ILOGIC_X0Y100_D = LIOB33_SING_X0Y100_IOB_X0Y100_I;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_D1 = CLBLL_L_X2Y107_SLICE_X1Y107_CQ;
  assign LIOI3_X0Y123_OLOGIC_X0Y124_T1 = 1'b1;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_D1 = CLBLL_L_X2Y107_SLICE_X1Y107_CQ;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A1 = CLBLL_L_X2Y109_SLICE_X0Y109_BO5;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A2 = CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A3 = CLBLL_L_X2Y109_SLICE_X0Y109_AQ;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A4 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_A6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign LIOI3_X0Y123_OLOGIC_X0Y123_T1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B1 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B2 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B3 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B4 = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B5 = CLBLL_L_X2Y106_SLICE_X0Y106_CQ;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_B6 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_C6 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D1 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D2 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D3 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D4 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D5 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X0Y109_D6 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A2 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A3 = CLBLL_L_X2Y109_SLICE_X1Y109_AQ;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A4 = CLBLM_R_X3Y107_SLICE_X2Y107_CO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A5 = CLBLL_L_X2Y109_SLICE_X0Y109_AQ;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_A6 = CLBLL_L_X2Y109_SLICE_X0Y109_BO5;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B1 = CLBLM_R_X3Y106_SLICE_X2Y106_CO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B2 = CLBLL_L_X2Y109_SLICE_X1Y109_BQ;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B3 = CLBLM_R_X3Y106_SLICE_X3Y106_BO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B4 = CLBLL_L_X2Y109_SLICE_X0Y109_BO5;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_B6 = CLBLL_L_X2Y110_SLICE_X0Y110_CQ;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C1 = CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C2 = CLBLL_L_X2Y109_SLICE_X1Y109_AQ;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C4 = CLBLM_R_X3Y110_SLICE_X2Y110_CQ;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C5 = CLBLL_L_X2Y106_SLICE_X0Y106_CQ;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_C6 = 1'b1;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D1 = CLBLL_L_X2Y108_SLICE_X1Y108_BO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D2 = CLBLL_L_X2Y109_SLICE_X1Y109_AQ;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D3 = LIOB33_X0Y111_IOB_X0Y111_I;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D4 = CLBLL_L_X4Y108_SLICE_X4Y108_AO6;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D5 = CLBLL_L_X2Y106_SLICE_X0Y106_CQ;
  assign CLBLL_L_X2Y109_SLICE_X1Y109_D6 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A1 = CLBLM_R_X3Y104_SLICE_X3Y104_DO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A3 = CLBLM_R_X3Y104_SLICE_X3Y104_AQ;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A4 = LIOB33_X0Y103_IOB_X0Y104_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_A6 = CLBLM_R_X3Y110_SLICE_X2Y110_CQ;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B2 = CLBLM_R_X3Y104_SLICE_X3Y104_BQ;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B3 = CLBLL_L_X4Y104_SLICE_X4Y104_AQ;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B5 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_B6 = CLBLM_R_X3Y104_SLICE_X3Y104_CO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C1 = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C2 = CLBLM_R_X3Y105_SLICE_X3Y105_AQ;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C3 = CLBLL_L_X2Y106_SLICE_X0Y106_DQ;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C4 = CLBLL_L_X4Y104_SLICE_X5Y104_BQ;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C5 = CLBLL_L_X4Y104_SLICE_X4Y104_AQ;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_C6 = CLBLL_L_X4Y104_SLICE_X5Y104_AQ;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D1 = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D2 = CLBLL_L_X4Y104_SLICE_X4Y104_BQ;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D3 = CLBLL_L_X2Y106_SLICE_X0Y106_DQ;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D4 = CLBLM_R_X3Y104_SLICE_X2Y104_CQ;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D5 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X3Y104_D6 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A1 = CLBLM_R_X3Y105_SLICE_X2Y105_CO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A2 = CLBLM_R_X3Y104_SLICE_X2Y104_BQ;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A3 = CLBLM_R_X3Y104_SLICE_X2Y104_AQ;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A5 = CLBLM_R_X3Y104_SLICE_X2Y104_CQ;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_A6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B1 = CLBLM_R_X3Y105_SLICE_X2Y105_CO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B2 = CLBLM_R_X3Y104_SLICE_X2Y104_BQ;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B3 = CLBLM_R_X3Y104_SLICE_X2Y104_AQ;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B4 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B5 = 1'b1;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_B6 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C1 = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C2 = CLBLM_R_X3Y104_SLICE_X2Y104_CQ;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C3 = CLBLM_R_X3Y104_SLICE_X2Y104_DQ;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C4 = CLBLL_L_X4Y104_SLICE_X4Y104_BQ;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_C6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D1 = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D2 = CLBLM_R_X3Y104_SLICE_X2Y104_CQ;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D3 = CLBLM_R_X3Y104_SLICE_X2Y104_DQ;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D4 = CLBLL_L_X4Y104_SLICE_X4Y104_BQ;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D5 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y104_SLICE_X2Y104_D6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D1 = CLBLM_R_X3Y110_SLICE_X2Y110_BQ;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y108_D = LIOB33_X0Y107_IOB_X0Y108_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D2 = CLBLM_R_X3Y108_SLICE_X3Y108_BO6;
  assign LIOI3_TBYTESRC_X0Y107_ILOGIC_X0Y107_D = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D3 = CLBLL_L_X4Y109_SLICE_X4Y109_DO6;
  assign CLBLL_L_X4Y108_SLICE_X4Y108_D5 = CLBLL_L_X2Y109_SLICE_X1Y109_CO6;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B5 = CLBLL_L_X2Y106_SLICE_X0Y106_BQ;
  assign CLBLL_L_X2Y106_SLICE_X0Y106_B6 = CLBLL_L_X2Y107_SLICE_X0Y107_AQ;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A1 = CLBLL_L_X2Y110_SLICE_X1Y110_AQ;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A3 = CLBLL_L_X2Y110_SLICE_X0Y110_AQ;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A4 = LIOB33_X0Y113_IOB_X0Y114_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A5 = CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_A6 = CLBLL_L_X2Y108_SLICE_X1Y108_AO5;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B2 = LIOB33_X0Y115_IOB_X0Y115_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B3 = CLBLL_L_X2Y110_SLICE_X0Y110_AQ;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B4 = CLBLL_L_X2Y108_SLICE_X1Y108_AO5;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B5 = CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_B6 = CLBLL_L_X2Y110_SLICE_X0Y110_BQ;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C1 = CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C2 = CLBLL_L_X2Y110_SLICE_X0Y110_CQ;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C3 = CLBLL_L_X2Y110_SLICE_X0Y110_BQ;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C5 = LIOB33_X0Y115_IOB_X0Y116_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_C6 = CLBLL_L_X2Y108_SLICE_X1Y108_AO5;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D3 = LIOB33_X0Y107_IOB_X0Y107_I;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D4 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X0Y110_D6 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A1 = CLBLL_L_X2Y110_SLICE_X1Y110_AQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A3 = LIOB33_X0Y113_IOB_X0Y113_I;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A4 = CLBLL_L_X2Y109_SLICE_X1Y109_AQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A5 = CLBLL_L_X2Y108_SLICE_X1Y108_AO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_A6 = CLBLL_L_X2Y108_SLICE_X1Y108_AO5;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B1 = CLBLM_R_X3Y109_SLICE_X3Y109_CQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B2 = CLBLL_L_X2Y109_SLICE_X0Y109_AQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B3 = CLBLL_L_X2Y110_SLICE_X1Y110_AQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B4 = CLBLL_L_X4Y109_SLICE_X5Y109_BQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B5 = CLBLL_L_X2Y110_SLICE_X0Y110_AQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_B6 = CLBLL_L_X2Y110_SLICE_X0Y110_CQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C1 = CLBLL_L_X2Y110_SLICE_X0Y110_AQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C2 = CLBLL_L_X2Y110_SLICE_X0Y110_BQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C3 = CLBLL_L_X4Y109_SLICE_X5Y109_AQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C4 = CLBLL_L_X2Y110_SLICE_X0Y110_CQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C5 = CLBLL_L_X2Y110_SLICE_X1Y110_AQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_C6 = CLBLL_L_X2Y109_SLICE_X1Y109_AQ;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D1 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D2 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D3 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D4 = CLBLL_L_X2Y110_SLICE_X1Y110_CO6;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D5 = 1'b1;
  assign CLBLL_L_X2Y110_SLICE_X1Y110_D6 = CLBLL_L_X2Y110_SLICE_X1Y110_BO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A1 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A2 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A3 = CLBLM_R_X3Y105_SLICE_X3Y105_AQ;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A4 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A5 = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_A6 = CLBLM_R_X3Y105_SLICE_X3Y105_A5Q;
  assign CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_CE = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_AX = CLBLM_R_X3Y105_SLICE_X3Y105_BO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B1 = CLBLM_R_X3Y105_SLICE_X3Y105_DO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B2 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B3 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B4 = CLBLM_R_X3Y104_SLICE_X3Y104_BQ;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B5 = CLBLM_R_X3Y105_SLICE_X3Y105_A5Q;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_B6 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C1 = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C2 = CLBLL_L_X2Y105_SLICE_X1Y105_AQ;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C3 = CLBLM_R_X3Y105_SLICE_X3Y105_A5Q;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C4 = CLBLM_R_X3Y104_SLICE_X2Y104_BQ;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C5 = CLBLM_R_X3Y105_SLICE_X3Y105_DO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_C6 = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D1 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D2 = CLBLL_L_X4Y104_SLICE_X5Y104_BQ;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D3 = CLBLL_L_X4Y104_SLICE_X4Y104_AQ;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D4 = CLBLL_L_X4Y105_SLICE_X5Y105_CO6;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D5 = CLBLL_L_X2Y106_SLICE_X0Y106_DQ;
  assign CLBLM_R_X3Y105_SLICE_X3Y105_D6 = CLBLM_R_X3Y104_SLICE_X3Y104_BQ;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A2 = CLBLM_R_X3Y105_SLICE_X2Y105_BQ;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A3 = CLBLM_R_X3Y105_SLICE_X2Y105_AQ;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A4 = CLBLM_R_X3Y105_SLICE_X2Y105_DO5;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A5 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_A6 = CLBLL_L_X2Y105_SLICE_X1Y105_AQ;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B1 = LIOB33_X0Y117_IOB_X0Y117_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B2 = CLBLM_R_X3Y105_SLICE_X2Y105_BQ;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B3 = CLBLM_R_X3Y105_SLICE_X2Y105_AQ;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C1 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B4 = CLBLM_R_X3Y105_SLICE_X2Y105_DO5;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B6 = LIOB33_X0Y105_IOB_X0Y106_I;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_B5 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C1 = CLBLM_R_X3Y104_SLICE_X2Y104_BQ;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C2 = CLBLM_R_X3Y105_SLICE_X3Y105_A5Q;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C3 = CLBLM_R_X3Y105_SLICE_X3Y105_DO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C4 = CLBLL_L_X4Y105_SLICE_X5Y105_BO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C5 = CLBLM_R_X3Y108_SLICE_X3Y108_DO6;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_C6 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_CLK = CLK_HROW_BOT_R_X139Y130_BUFHCE_X0Y32_O;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_C6 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D1 = CLBLM_R_X3Y105_SLICE_X2Y105_CO5;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D2 = CLBLM_R_X5Y105_SLICE_X6Y105_CQ;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D3 = CLBLL_L_X2Y106_SLICE_X0Y106_DQ;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D4 = 1'b1;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D5 = CLBLL_L_X2Y105_SLICE_X1Y105_AQ;
  assign CLBLM_R_X3Y105_SLICE_X2Y105_D6 = 1'b1;
  assign LIOI3_X0Y109_ILOGIC_X0Y110_D = LIOB33_X0Y109_IOB_X0Y110_I;
  assign LIOI3_X0Y109_ILOGIC_X0Y109_D = LIOB33_X0Y109_IOB_X0Y109_I;
  assign CLBLL_L_X4Y108_SLICE_X5Y108_D1 = 1'b1;
endmodule
